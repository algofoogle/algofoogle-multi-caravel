magic
tech gf180mcuD
magscale 1 5
timestamp 1702351428
<< obsm1 >>
rect 672 1538 65856 99206
<< metal2 >>
rect 2912 0 2968 400
rect 4256 0 4312 400
rect 5600 0 5656 400
rect 6944 0 7000 400
rect 8288 0 8344 400
rect 9632 0 9688 400
rect 10976 0 11032 400
rect 12320 0 12376 400
rect 13664 0 13720 400
rect 15008 0 15064 400
rect 16352 0 16408 400
rect 17696 0 17752 400
rect 19040 0 19096 400
rect 20384 0 20440 400
rect 21728 0 21784 400
rect 23072 0 23128 400
rect 24416 0 24472 400
rect 25760 0 25816 400
rect 27104 0 27160 400
rect 28448 0 28504 400
rect 29792 0 29848 400
rect 31136 0 31192 400
rect 32480 0 32536 400
rect 33824 0 33880 400
rect 35168 0 35224 400
rect 36512 0 36568 400
rect 37856 0 37912 400
rect 39200 0 39256 400
rect 40544 0 40600 400
rect 41888 0 41944 400
rect 43232 0 43288 400
rect 44576 0 44632 400
rect 45920 0 45976 400
rect 47264 0 47320 400
rect 48608 0 48664 400
rect 49952 0 50008 400
rect 51296 0 51352 400
rect 52640 0 52696 400
rect 53984 0 54040 400
rect 55328 0 55384 400
rect 56672 0 56728 400
rect 58016 0 58072 400
rect 59360 0 59416 400
rect 60704 0 60760 400
rect 62048 0 62104 400
rect 63392 0 63448 400
<< obsm2 >>
rect 518 430 65730 99195
rect 518 400 2882 430
rect 2998 400 4226 430
rect 4342 400 5570 430
rect 5686 400 6914 430
rect 7030 400 8258 430
rect 8374 400 9602 430
rect 9718 400 10946 430
rect 11062 400 12290 430
rect 12406 400 13634 430
rect 13750 400 14978 430
rect 15094 400 16322 430
rect 16438 400 17666 430
rect 17782 400 19010 430
rect 19126 400 20354 430
rect 20470 400 21698 430
rect 21814 400 23042 430
rect 23158 400 24386 430
rect 24502 400 25730 430
rect 25846 400 27074 430
rect 27190 400 28418 430
rect 28534 400 29762 430
rect 29878 400 31106 430
rect 31222 400 32450 430
rect 32566 400 33794 430
rect 33910 400 35138 430
rect 35254 400 36482 430
rect 36598 400 37826 430
rect 37942 400 39170 430
rect 39286 400 40514 430
rect 40630 400 41858 430
rect 41974 400 43202 430
rect 43318 400 44546 430
rect 44662 400 45890 430
rect 46006 400 47234 430
rect 47350 400 48578 430
rect 48694 400 49922 430
rect 50038 400 51266 430
rect 51382 400 52610 430
rect 52726 400 53954 430
rect 54070 400 55298 430
rect 55414 400 56642 430
rect 56758 400 57986 430
rect 58102 400 59330 430
rect 59446 400 60674 430
rect 60790 400 62018 430
rect 62134 400 63362 430
rect 63478 400 65730 430
<< obsm3 >>
rect 513 1246 65735 99190
<< metal4 >>
rect 2224 1538 2384 99206
rect 9904 1538 10064 99206
rect 17584 1538 17744 99206
rect 25264 1538 25424 99206
rect 32944 1538 33104 99206
rect 40624 1538 40784 99206
rect 48304 1538 48464 99206
rect 55984 1538 56144 99206
rect 63664 1538 63824 99206
<< obsm4 >>
rect 854 1801 2194 97879
rect 2414 1801 9874 97879
rect 10094 1801 17554 97879
rect 17774 1801 25234 97879
rect 25454 1801 32914 97879
rect 33134 1801 40594 97879
rect 40814 1801 48274 97879
rect 48494 1801 55954 97879
rect 56174 1801 63602 97879
<< labels >>
rlabel metal2 s 2912 0 2968 400 6 i_clk
port 1 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal2 s 47264 0 47320 400 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 49952 0 50008 400 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 20384 0 20440 400 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 19040 0 19096 400 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 17696 0 17752 400 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 16352 0 16408 400 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal2 s 15008 0 15064 400 6 i_gpout1_sel[0]
port 9 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 i_gpout1_sel[1]
port 10 nsew signal input
rlabel metal2 s 12320 0 12376 400 6 i_gpout1_sel[2]
port 11 nsew signal input
rlabel metal2 s 10976 0 11032 400 6 i_gpout1_sel[3]
port 12 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 i_gpout2_sel[0]
port 13 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 i_gpout2_sel[1]
port 14 nsew signal input
rlabel metal2 s 6944 0 7000 400 6 i_gpout2_sel[2]
port 15 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 i_gpout2_sel[3]
port 16 nsew signal input
rlabel metal2 s 44576 0 44632 400 6 i_mode[0]
port 17 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 i_mode[1]
port 18 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 i_mode[2]
port 19 nsew signal input
rlabel metal2 s 53984 0 54040 400 6 i_reg_csb
port 20 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 i_reg_mosi
port 21 nsew signal input
rlabel metal2 s 45920 0 45976 400 6 i_reg_outs_enb
port 22 nsew signal input
rlabel metal2 s 52640 0 52696 400 6 i_reg_sclk
port 23 nsew signal input
rlabel metal2 s 4256 0 4312 400 6 i_reset
port 24 nsew signal input
rlabel metal2 s 63392 0 63448 400 6 i_tex_in[0]
port 25 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 i_tex_in[1]
port 26 nsew signal input
rlabel metal2 s 60704 0 60760 400 6 i_tex_in[2]
port 27 nsew signal input
rlabel metal2 s 59360 0 59416 400 6 i_tex_in[3]
port 28 nsew signal input
rlabel metal2 s 58016 0 58072 400 6 i_vec_csb
port 29 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 i_vec_mosi
port 30 nsew signal input
rlabel metal2 s 56672 0 56728 400 6 i_vec_sclk
port 31 nsew signal input
rlabel metal2 s 24416 0 24472 400 6 o_gpout[0]
port 32 nsew signal output
rlabel metal2 s 23072 0 23128 400 6 o_gpout[1]
port 33 nsew signal output
rlabel metal2 s 21728 0 21784 400 6 o_gpout[2]
port 34 nsew signal output
rlabel metal2 s 40544 0 40600 400 6 o_hsync
port 35 nsew signal output
rlabel metal2 s 37856 0 37912 400 6 o_rgb[0]
port 36 nsew signal output
rlabel metal2 s 36512 0 36568 400 6 o_rgb[1]
port 37 nsew signal output
rlabel metal2 s 35168 0 35224 400 6 o_rgb[2]
port 38 nsew signal output
rlabel metal2 s 33824 0 33880 400 6 o_rgb[3]
port 39 nsew signal output
rlabel metal2 s 32480 0 32536 400 6 o_rgb[4]
port 40 nsew signal output
rlabel metal2 s 31136 0 31192 400 6 o_rgb[5]
port 41 nsew signal output
rlabel metal2 s 29792 0 29848 400 6 o_tex_csb
port 42 nsew signal output
rlabel metal2 s 25760 0 25816 400 6 o_tex_oeb0
port 43 nsew signal output
rlabel metal2 s 27104 0 27160 400 6 o_tex_out0
port 44 nsew signal output
rlabel metal2 s 28448 0 28504 400 6 o_tex_sclk
port 45 nsew signal output
rlabel metal2 s 39200 0 39256 400 6 o_vsync
port 46 nsew signal output
rlabel metal4 s 2224 1538 2384 99206 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 99206 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 99206 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 99206 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 99206 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 99206 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 99206 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 99206 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 99206 6 vss
port 48 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 66563 100965
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 25139744
string GDS_FILE /home/zerotoasic/anton/algofoogle-multi-caravel/openlane/top_raybox_zero_fsm/runs/23_12_12_13_43/results/signoff/top_raybox_zero_fsm.magic.gds
string GDS_START 599310
<< end >>

