magic
tech gf180mcuD
magscale 1 10
timestamp 1702302760
<< nwell >>
rect 1258 48985 48806 49824
rect 1258 48960 15677 48985
rect 1258 47417 48806 48256
rect 1258 47392 11197 47417
rect 1258 46663 14557 46688
rect 1258 45849 48806 46663
rect 1258 45824 9517 45849
rect 1258 45095 28221 45120
rect 1258 44281 48806 45095
rect 1258 44256 8733 44281
rect 1258 43527 5933 43552
rect 1258 42713 48806 43527
rect 1258 42688 16685 42713
rect 1258 41959 20605 41984
rect 1258 41145 48806 41959
rect 1258 41120 10749 41145
rect 1258 40391 3805 40416
rect 1258 39577 48806 40391
rect 1258 39552 18141 39577
rect 1258 38823 3021 38848
rect 1258 38009 48806 38823
rect 1258 37984 12181 38009
rect 1258 37255 3021 37280
rect 1258 36441 48806 37255
rect 1258 36416 16797 36441
rect 1258 35687 6829 35712
rect 1258 34873 48806 35687
rect 1258 34848 3021 34873
rect 1258 34119 15117 34144
rect 1258 33305 48806 34119
rect 1258 33280 7277 33305
rect 1258 32551 3021 32576
rect 1258 31737 48806 32551
rect 1258 31712 16461 31737
rect 1258 30983 7165 31008
rect 1258 30169 48806 30983
rect 1258 30144 3021 30169
rect 1258 29415 43229 29440
rect 1258 28601 48806 29415
rect 1258 28576 3133 28601
rect 1258 27847 7277 27872
rect 1258 27033 48806 27847
rect 1258 27008 5924 27033
rect 1258 26279 3021 26304
rect 1258 25465 48806 26279
rect 1258 25440 9063 25465
rect 1258 24711 3245 24736
rect 1258 23897 48806 24711
rect 1258 23872 11409 23897
rect 1258 23143 3021 23168
rect 1258 22329 48806 23143
rect 1258 22304 7949 22329
rect 1258 21575 3133 21600
rect 1258 20761 48806 21575
rect 1258 20736 13872 20761
rect 1258 20007 7277 20032
rect 1258 19193 48806 20007
rect 1258 19168 3021 19193
rect 1258 18439 18125 18464
rect 1258 17625 48806 18439
rect 1258 17600 29327 17625
rect 1258 16871 3021 16896
rect 1258 16057 48806 16871
rect 1258 16032 39165 16057
rect 1258 15303 12397 15328
rect 1258 14489 48806 15303
rect 1258 14464 3021 14489
rect 1258 13735 4813 13760
rect 1258 12921 48806 13735
rect 1258 12896 39880 12921
rect 1258 12167 3021 12192
rect 1258 11353 48806 12167
rect 1258 11328 9293 11353
rect 1258 10599 3021 10624
rect 1258 9785 48806 10599
rect 1258 9760 24941 9785
rect 1258 9031 20031 9056
rect 1258 8217 48806 9031
rect 1258 8192 3021 8217
rect 1258 7463 25303 7488
rect 1258 6649 48806 7463
rect 1258 6624 32669 6649
rect 1258 5895 3021 5920
rect 1258 5081 48806 5895
rect 1258 5056 9597 5081
rect 1258 4327 3133 4352
rect 1258 3488 48806 4327
<< pwell >>
rect 1258 49824 48806 50262
rect 1258 48256 48806 48960
rect 1258 46688 48806 47392
rect 1258 45120 48806 45824
rect 1258 43552 48806 44256
rect 1258 41984 48806 42688
rect 1258 40416 48806 41120
rect 1258 38848 48806 39552
rect 1258 37280 48806 37984
rect 1258 35712 48806 36416
rect 1258 34144 48806 34848
rect 1258 32576 48806 33280
rect 1258 31008 48806 31712
rect 1258 29440 48806 30144
rect 1258 27872 48806 28576
rect 1258 26304 48806 27008
rect 1258 24736 48806 25440
rect 1258 23168 48806 23872
rect 1258 21600 48806 22304
rect 1258 20032 48806 20736
rect 1258 18464 48806 19168
rect 1258 16896 48806 17600
rect 1258 15328 48806 16032
rect 1258 13760 48806 14464
rect 1258 12192 48806 12896
rect 1258 10624 48806 11328
rect 1258 9056 48806 9760
rect 1258 7488 48806 8192
rect 1258 5920 48806 6624
rect 1258 4352 48806 5056
rect 1258 3050 48806 3488
<< obsm1 >>
rect 1344 3076 48720 50370
<< metal2 >>
rect 2016 0 2128 800
rect 3136 0 3248 800
rect 4256 0 4368 800
rect 5376 0 5488 800
rect 6496 0 6608 800
rect 7616 0 7728 800
rect 8736 0 8848 800
rect 9856 0 9968 800
rect 10976 0 11088 800
rect 12096 0 12208 800
rect 13216 0 13328 800
rect 14336 0 14448 800
rect 15456 0 15568 800
rect 16576 0 16688 800
rect 17696 0 17808 800
rect 18816 0 18928 800
rect 19936 0 20048 800
rect 21056 0 21168 800
rect 22176 0 22288 800
rect 23296 0 23408 800
rect 24416 0 24528 800
rect 25536 0 25648 800
rect 26656 0 26768 800
rect 27776 0 27888 800
rect 28896 0 29008 800
rect 30016 0 30128 800
rect 31136 0 31248 800
rect 32256 0 32368 800
rect 33376 0 33488 800
rect 34496 0 34608 800
rect 35616 0 35728 800
rect 36736 0 36848 800
rect 37856 0 37968 800
rect 38976 0 39088 800
rect 40096 0 40208 800
rect 41216 0 41328 800
rect 42336 0 42448 800
rect 43456 0 43568 800
rect 44576 0 44688 800
rect 45696 0 45808 800
rect 46816 0 46928 800
rect 47936 0 48048 800
<< obsm2 >>
rect 1708 860 48468 50382
rect 1708 700 1956 860
rect 2188 700 3076 860
rect 3308 700 4196 860
rect 4428 700 5316 860
rect 5548 700 6436 860
rect 6668 700 7556 860
rect 7788 700 8676 860
rect 8908 700 9796 860
rect 10028 700 10916 860
rect 11148 700 12036 860
rect 12268 700 13156 860
rect 13388 700 14276 860
rect 14508 700 15396 860
rect 15628 700 16516 860
rect 16748 700 17636 860
rect 17868 700 18756 860
rect 18988 700 19876 860
rect 20108 700 20996 860
rect 21228 700 22116 860
rect 22348 700 23236 860
rect 23468 700 24356 860
rect 24588 700 25476 860
rect 25708 700 26596 860
rect 26828 700 27716 860
rect 27948 700 28836 860
rect 29068 700 29956 860
rect 30188 700 31076 860
rect 31308 700 32196 860
rect 32428 700 33316 860
rect 33548 700 34436 860
rect 34668 700 35556 860
rect 35788 700 36676 860
rect 36908 700 37796 860
rect 38028 700 38916 860
rect 39148 700 40036 860
rect 40268 700 41156 860
rect 41388 700 42276 860
rect 42508 700 43396 860
rect 43628 700 44516 860
rect 44748 700 45636 860
rect 45868 700 46756 860
rect 46988 700 47876 860
rect 48108 700 48468 860
<< obsm3 >>
rect 1698 2940 48478 50204
<< metal4 >>
rect 4448 3076 4768 50236
rect 19808 3076 20128 50236
rect 35168 3076 35488 50236
<< obsm4 >>
rect 9212 11890 19748 41310
rect 20188 11890 35108 41310
rect 35548 11890 37940 41310
<< labels >>
rlabel metal2 s 2016 0 2128 800 6 clk
port 1 nsew signal input
rlabel metal2 s 3136 0 3248 800 6 rst
port 2 nsew signal input
rlabel metal2 s 12096 0 12208 800 6 ui_in[0]
port 3 nsew signal input
rlabel metal2 s 10976 0 11088 800 6 ui_in[1]
port 4 nsew signal input
rlabel metal2 s 9856 0 9968 800 6 ui_in[2]
port 5 nsew signal input
rlabel metal2 s 8736 0 8848 800 6 ui_in[3]
port 6 nsew signal input
rlabel metal2 s 7616 0 7728 800 6 ui_in[4]
port 7 nsew signal input
rlabel metal2 s 6496 0 6608 800 6 ui_in[5]
port 8 nsew signal input
rlabel metal2 s 5376 0 5488 800 6 ui_in[6]
port 9 nsew signal input
rlabel metal2 s 4256 0 4368 800 6 ui_in[7]
port 10 nsew signal input
rlabel metal2 s 21056 0 21168 800 6 uio_in[0]
port 11 nsew signal input
rlabel metal2 s 19936 0 20048 800 6 uio_in[1]
port 12 nsew signal input
rlabel metal2 s 18816 0 18928 800 6 uio_in[2]
port 13 nsew signal input
rlabel metal2 s 17696 0 17808 800 6 uio_in[3]
port 14 nsew signal input
rlabel metal2 s 16576 0 16688 800 6 uio_in[4]
port 15 nsew signal input
rlabel metal2 s 15456 0 15568 800 6 uio_in[5]
port 16 nsew signal input
rlabel metal2 s 14336 0 14448 800 6 uio_in[6]
port 17 nsew signal input
rlabel metal2 s 13216 0 13328 800 6 uio_in[7]
port 18 nsew signal input
rlabel metal2 s 47936 0 48048 800 6 uio_oe[0]
port 19 nsew signal output
rlabel metal2 s 46816 0 46928 800 6 uio_oe[1]
port 20 nsew signal output
rlabel metal2 s 45696 0 45808 800 6 uio_oe[2]
port 21 nsew signal output
rlabel metal2 s 44576 0 44688 800 6 uio_oe[3]
port 22 nsew signal output
rlabel metal2 s 43456 0 43568 800 6 uio_oe[4]
port 23 nsew signal output
rlabel metal2 s 42336 0 42448 800 6 uio_oe[5]
port 24 nsew signal output
rlabel metal2 s 41216 0 41328 800 6 uio_oe[6]
port 25 nsew signal output
rlabel metal2 s 40096 0 40208 800 6 uio_oe[7]
port 26 nsew signal output
rlabel metal2 s 38976 0 39088 800 6 uio_out[0]
port 27 nsew signal output
rlabel metal2 s 37856 0 37968 800 6 uio_out[1]
port 28 nsew signal output
rlabel metal2 s 36736 0 36848 800 6 uio_out[2]
port 29 nsew signal output
rlabel metal2 s 35616 0 35728 800 6 uio_out[3]
port 30 nsew signal output
rlabel metal2 s 34496 0 34608 800 6 uio_out[4]
port 31 nsew signal output
rlabel metal2 s 33376 0 33488 800 6 uio_out[5]
port 32 nsew signal output
rlabel metal2 s 32256 0 32368 800 6 uio_out[6]
port 33 nsew signal output
rlabel metal2 s 31136 0 31248 800 6 uio_out[7]
port 34 nsew signal output
rlabel metal2 s 30016 0 30128 800 6 uo_out[0]
port 35 nsew signal output
rlabel metal2 s 28896 0 29008 800 6 uo_out[1]
port 36 nsew signal output
rlabel metal2 s 27776 0 27888 800 6 uo_out[2]
port 37 nsew signal output
rlabel metal2 s 26656 0 26768 800 6 uo_out[3]
port 38 nsew signal output
rlabel metal2 s 25536 0 25648 800 6 uo_out[4]
port 39 nsew signal output
rlabel metal2 s 24416 0 24528 800 6 uo_out[5]
port 40 nsew signal output
rlabel metal2 s 23296 0 23408 800 6 uo_out[6]
port 41 nsew signal output
rlabel metal2 s 22176 0 22288 800 6 uo_out[7]
port 42 nsew signal output
rlabel metal4 s 4448 3076 4768 50236 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 50236 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 50236 6 vss
port 44 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 50087 53671
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2226910
string GDS_FILE /home/zerotoasic/anton/algofoogle-multi-caravel/openlane/top_vga_spi_rom/runs/23_12_12_00_21/results/signoff/top_vga_spi_rom.magic.gds
string GDS_START 348292
<< end >>

