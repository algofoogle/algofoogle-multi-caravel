magic
tech gf180mcuD
magscale 1 10
timestamp 1702289012
<< nwell >>
rect 1258 41120 40070 41638
rect 1258 39577 40070 40416
rect 1258 39552 11880 39577
rect 1258 38009 40070 38848
rect 1258 37984 18464 38009
rect 1258 37255 27336 37280
rect 1258 36416 40070 37255
rect 1258 35687 6909 35712
rect 1258 34873 40070 35687
rect 1258 34848 6461 34873
rect 1258 34119 26061 34144
rect 1258 33305 40070 34119
rect 1258 33280 7870 33305
rect 1258 32551 22072 32576
rect 1258 31737 40070 32551
rect 1258 31712 8990 31737
rect 1258 30983 3661 31008
rect 1258 30169 40070 30983
rect 1258 30144 26686 30169
rect 1258 29415 2653 29440
rect 1258 28601 40070 29415
rect 1258 28576 11856 28601
rect 1258 27847 4669 27872
rect 1258 27033 40070 27847
rect 1258 27008 2541 27033
rect 1258 26279 20797 26304
rect 1258 25465 40070 26279
rect 1258 25440 15352 25465
rect 1258 24711 2998 24736
rect 1258 23897 40070 24711
rect 1258 23872 9149 23897
rect 1258 23143 14344 23168
rect 1258 22329 40070 23143
rect 1258 22304 7712 22329
rect 1258 21575 27853 21600
rect 1258 20761 40070 21575
rect 1258 20736 2541 20761
rect 1258 20007 23214 20032
rect 1258 19168 40070 20007
rect 1258 18439 33472 18464
rect 1258 17625 40070 18439
rect 1258 17600 2541 17625
rect 1258 16871 27517 16896
rect 1258 16057 40070 16871
rect 1258 16032 33496 16057
rect 1258 15303 14568 15328
rect 1258 14464 40070 15303
rect 1258 13735 2653 13760
rect 1258 12921 40070 13735
rect 1258 12896 26993 12921
rect 1258 12167 3101 12192
rect 1258 11353 40070 12167
rect 1258 11328 15576 11353
rect 1258 10599 21917 10624
rect 1258 9760 40070 10599
rect 1258 9031 2541 9056
rect 1258 8217 40070 9031
rect 1258 8192 18376 8217
rect 1258 7463 2765 7488
rect 1258 6649 40070 7463
rect 1258 6624 18669 6649
rect 1258 5081 40070 5920
rect 1258 5056 2653 5081
rect 1258 4327 21512 4352
rect 1258 3488 40070 4327
<< pwell >>
rect 1258 40416 40070 41120
rect 1258 38848 40070 39552
rect 1258 37280 40070 37984
rect 1258 35712 40070 36416
rect 1258 34144 40070 34848
rect 1258 32576 40070 33280
rect 1258 31008 40070 31712
rect 1258 29440 40070 30144
rect 1258 27872 40070 28576
rect 1258 26304 40070 27008
rect 1258 24736 40070 25440
rect 1258 23168 40070 23872
rect 1258 21600 40070 22304
rect 1258 20032 40070 20736
rect 1258 18464 40070 19168
rect 1258 16896 40070 17600
rect 1258 15328 40070 16032
rect 1258 13760 40070 14464
rect 1258 12192 40070 12896
rect 1258 10624 40070 11328
rect 1258 9056 40070 9760
rect 1258 7488 40070 8192
rect 1258 5920 40070 6624
rect 1258 4352 40070 5056
rect 1258 3050 40070 3488
<< obsm1 >>
rect 1344 3076 39984 41612
<< metal2 >>
rect 1792 0 1904 800
rect 3136 0 3248 800
rect 4480 0 4592 800
rect 5824 0 5936 800
rect 7168 0 7280 800
rect 8512 0 8624 800
rect 9856 0 9968 800
rect 11200 0 11312 800
rect 12544 0 12656 800
rect 13888 0 14000 800
rect 15232 0 15344 800
rect 16576 0 16688 800
rect 17920 0 18032 800
rect 19264 0 19376 800
rect 20608 0 20720 800
rect 21952 0 22064 800
rect 23296 0 23408 800
rect 24640 0 24752 800
rect 25984 0 26096 800
rect 27328 0 27440 800
rect 28672 0 28784 800
rect 30016 0 30128 800
rect 31360 0 31472 800
rect 32704 0 32816 800
rect 34048 0 34160 800
rect 35392 0 35504 800
rect 36736 0 36848 800
rect 38080 0 38192 800
rect 39424 0 39536 800
<< obsm2 >>
rect 1820 860 39732 41590
rect 1964 800 3076 860
rect 3308 800 4420 860
rect 4652 800 5764 860
rect 5996 800 7108 860
rect 7340 800 8452 860
rect 8684 800 9796 860
rect 10028 800 11140 860
rect 11372 800 12484 860
rect 12716 800 13828 860
rect 14060 800 15172 860
rect 15404 800 16516 860
rect 16748 800 17860 860
rect 18092 800 19204 860
rect 19436 800 20548 860
rect 20780 800 21892 860
rect 22124 800 23236 860
rect 23468 800 24580 860
rect 24812 800 25924 860
rect 26156 800 27268 860
rect 27500 800 28612 860
rect 28844 800 29956 860
rect 30188 800 31300 860
rect 31532 800 32644 860
rect 32876 800 33988 860
rect 34220 800 35332 860
rect 35564 800 36676 860
rect 36908 800 38020 860
rect 38252 800 39364 860
rect 39596 800 39732 860
<< obsm3 >>
rect 1810 3108 39742 41580
<< metal4 >>
rect 4448 3076 4768 41612
rect 19808 3076 20128 41612
rect 35168 3076 35488 41612
<< obsm4 >>
rect 8204 6290 19748 33246
rect 20188 6290 35108 33246
rect 35548 6290 37716 33246
<< labels >>
rlabel metal2 s 1792 0 1904 800 6 clk
port 1 nsew signal input
rlabel metal2 s 4480 0 4592 800 6 gpio_ready
port 2 nsew signal input
rlabel metal2 s 39424 0 39536 800 6 io_in[0]
port 3 nsew signal input
rlabel metal2 s 25984 0 26096 800 6 io_in[10]
port 4 nsew signal input
rlabel metal2 s 24640 0 24752 800 6 io_in[11]
port 5 nsew signal input
rlabel metal2 s 23296 0 23408 800 6 io_in[12]
port 6 nsew signal input
rlabel metal2 s 38080 0 38192 800 6 io_in[1]
port 7 nsew signal input
rlabel metal2 s 36736 0 36848 800 6 io_in[2]
port 8 nsew signal input
rlabel metal2 s 35392 0 35504 800 6 io_in[3]
port 9 nsew signal input
rlabel metal2 s 34048 0 34160 800 6 io_in[4]
port 10 nsew signal input
rlabel metal2 s 32704 0 32816 800 6 io_in[5]
port 11 nsew signal input
rlabel metal2 s 31360 0 31472 800 6 io_in[6]
port 12 nsew signal input
rlabel metal2 s 30016 0 30128 800 6 io_in[7]
port 13 nsew signal input
rlabel metal2 s 28672 0 28784 800 6 io_in[8]
port 14 nsew signal input
rlabel metal2 s 27328 0 27440 800 6 io_in[9]
port 15 nsew signal input
rlabel metal2 s 21952 0 22064 800 6 io_out[0]
port 16 nsew signal output
rlabel metal2 s 8512 0 8624 800 6 io_out[10]
port 17 nsew signal output
rlabel metal2 s 7168 0 7280 800 6 io_out[11]
port 18 nsew signal output
rlabel metal2 s 5824 0 5936 800 6 io_out[12]
port 19 nsew signal output
rlabel metal2 s 20608 0 20720 800 6 io_out[1]
port 20 nsew signal output
rlabel metal2 s 19264 0 19376 800 6 io_out[2]
port 21 nsew signal output
rlabel metal2 s 17920 0 18032 800 6 io_out[3]
port 22 nsew signal output
rlabel metal2 s 16576 0 16688 800 6 io_out[4]
port 23 nsew signal output
rlabel metal2 s 15232 0 15344 800 6 io_out[5]
port 24 nsew signal output
rlabel metal2 s 13888 0 14000 800 6 io_out[6]
port 25 nsew signal output
rlabel metal2 s 12544 0 12656 800 6 io_out[7]
port 26 nsew signal output
rlabel metal2 s 11200 0 11312 800 6 io_out[8]
port 27 nsew signal output
rlabel metal2 s 9856 0 9968 800 6 io_out[9]
port 28 nsew signal output
rlabel metal2 s 3136 0 3248 800 6 rst
port 29 nsew signal input
rlabel metal4 s 4448 3076 4768 41612 6 vdd
port 30 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 41612 6 vdd
port 30 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 41612 6 vss
port 31 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 41437 45021
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1326800
string GDS_FILE /home/zerotoasic/anton/algofoogle-multi-caravel/openlane/top_solo_squash/runs/23_12_11_20_32/results/signoff/top_solo_squash.magic.gds
string GDS_START 265422
<< end >>

