VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_design_mux
  CLASS BLOCK ;
  FOREIGN top_design_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 2400.000 BY 300.000 ;
  PIN diego_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1434.720 0.000 1435.280 4.000 ;
    END
  END diego_clk
  PIN diego_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1448.160 0.000 1448.720 4.000 ;
    END
  END diego_ena
  PIN diego_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1884.960 0.000 1885.520 4.000 ;
    END
  END diego_io_in[0]
  PIN diego_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1952.160 0.000 1952.720 4.000 ;
    END
  END diego_io_in[10]
  PIN diego_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1958.880 0.000 1959.440 4.000 ;
    END
  END diego_io_in[11]
  PIN diego_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1965.600 0.000 1966.160 4.000 ;
    END
  END diego_io_in[12]
  PIN diego_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1972.320 0.000 1972.880 4.000 ;
    END
  END diego_io_in[13]
  PIN diego_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1979.040 0.000 1979.600 4.000 ;
    END
  END diego_io_in[14]
  PIN diego_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1985.760 0.000 1986.320 4.000 ;
    END
  END diego_io_in[15]
  PIN diego_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1992.480 0.000 1993.040 4.000 ;
    END
  END diego_io_in[16]
  PIN diego_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1999.200 0.000 1999.760 4.000 ;
    END
  END diego_io_in[17]
  PIN diego_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2005.920 0.000 2006.480 4.000 ;
    END
  END diego_io_in[18]
  PIN diego_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2012.640 0.000 2013.200 4.000 ;
    END
  END diego_io_in[19]
  PIN diego_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1891.680 0.000 1892.240 4.000 ;
    END
  END diego_io_in[1]
  PIN diego_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2019.360 0.000 2019.920 4.000 ;
    END
  END diego_io_in[20]
  PIN diego_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2026.080 0.000 2026.640 4.000 ;
    END
  END diego_io_in[21]
  PIN diego_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2032.800 0.000 2033.360 4.000 ;
    END
  END diego_io_in[22]
  PIN diego_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2039.520 0.000 2040.080 4.000 ;
    END
  END diego_io_in[23]
  PIN diego_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2046.240 0.000 2046.800 4.000 ;
    END
  END diego_io_in[24]
  PIN diego_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2052.960 0.000 2053.520 4.000 ;
    END
  END diego_io_in[25]
  PIN diego_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2059.680 0.000 2060.240 4.000 ;
    END
  END diego_io_in[26]
  PIN diego_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2066.400 0.000 2066.960 4.000 ;
    END
  END diego_io_in[27]
  PIN diego_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2073.120 0.000 2073.680 4.000 ;
    END
  END diego_io_in[28]
  PIN diego_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2079.840 0.000 2080.400 4.000 ;
    END
  END diego_io_in[29]
  PIN diego_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1898.400 0.000 1898.960 4.000 ;
    END
  END diego_io_in[2]
  PIN diego_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2086.560 0.000 2087.120 4.000 ;
    END
  END diego_io_in[30]
  PIN diego_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2093.280 0.000 2093.840 4.000 ;
    END
  END diego_io_in[31]
  PIN diego_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2100.000 0.000 2100.560 4.000 ;
    END
  END diego_io_in[32]
  PIN diego_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2106.720 0.000 2107.280 4.000 ;
    END
  END diego_io_in[33]
  PIN diego_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2113.440 0.000 2114.000 4.000 ;
    END
  END diego_io_in[34]
  PIN diego_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2120.160 0.000 2120.720 4.000 ;
    END
  END diego_io_in[35]
  PIN diego_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2126.880 0.000 2127.440 4.000 ;
    END
  END diego_io_in[36]
  PIN diego_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2133.600 0.000 2134.160 4.000 ;
    END
  END diego_io_in[37]
  PIN diego_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1905.120 0.000 1905.680 4.000 ;
    END
  END diego_io_in[3]
  PIN diego_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1911.840 0.000 1912.400 4.000 ;
    END
  END diego_io_in[4]
  PIN diego_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1918.560 0.000 1919.120 4.000 ;
    END
  END diego_io_in[5]
  PIN diego_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1925.280 0.000 1925.840 4.000 ;
    END
  END diego_io_in[6]
  PIN diego_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1932.000 0.000 1932.560 4.000 ;
    END
  END diego_io_in[7]
  PIN diego_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1938.720 0.000 1939.280 4.000 ;
    END
  END diego_io_in[8]
  PIN diego_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1945.440 0.000 1946.000 4.000 ;
    END
  END diego_io_in[9]
  PIN diego_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1669.920 0.000 1670.480 4.000 ;
    END
  END diego_io_oeb[0]
  PIN diego_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1737.120 0.000 1737.680 4.000 ;
    END
  END diego_io_oeb[10]
  PIN diego_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1743.840 0.000 1744.400 4.000 ;
    END
  END diego_io_oeb[11]
  PIN diego_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1750.560 0.000 1751.120 4.000 ;
    END
  END diego_io_oeb[12]
  PIN diego_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1757.280 0.000 1757.840 4.000 ;
    END
  END diego_io_oeb[13]
  PIN diego_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1764.000 0.000 1764.560 4.000 ;
    END
  END diego_io_oeb[14]
  PIN diego_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1770.720 0.000 1771.280 4.000 ;
    END
  END diego_io_oeb[15]
  PIN diego_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1777.440 0.000 1778.000 4.000 ;
    END
  END diego_io_oeb[16]
  PIN diego_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1784.160 0.000 1784.720 4.000 ;
    END
  END diego_io_oeb[17]
  PIN diego_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1790.880 0.000 1791.440 4.000 ;
    END
  END diego_io_oeb[18]
  PIN diego_io_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1797.600 0.000 1798.160 4.000 ;
    END
  END diego_io_oeb[19]
  PIN diego_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1676.640 0.000 1677.200 4.000 ;
    END
  END diego_io_oeb[1]
  PIN diego_io_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1804.320 0.000 1804.880 4.000 ;
    END
  END diego_io_oeb[20]
  PIN diego_io_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1811.040 0.000 1811.600 4.000 ;
    END
  END diego_io_oeb[21]
  PIN diego_io_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1817.760 0.000 1818.320 4.000 ;
    END
  END diego_io_oeb[22]
  PIN diego_io_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1824.480 0.000 1825.040 4.000 ;
    END
  END diego_io_oeb[23]
  PIN diego_io_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1831.200 0.000 1831.760 4.000 ;
    END
  END diego_io_oeb[24]
  PIN diego_io_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1837.920 0.000 1838.480 4.000 ;
    END
  END diego_io_oeb[25]
  PIN diego_io_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1844.640 0.000 1845.200 4.000 ;
    END
  END diego_io_oeb[26]
  PIN diego_io_oeb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1851.360 0.000 1851.920 4.000 ;
    END
  END diego_io_oeb[27]
  PIN diego_io_oeb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1858.080 0.000 1858.640 4.000 ;
    END
  END diego_io_oeb[28]
  PIN diego_io_oeb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1864.800 0.000 1865.360 4.000 ;
    END
  END diego_io_oeb[29]
  PIN diego_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1683.360 0.000 1683.920 4.000 ;
    END
  END diego_io_oeb[2]
  PIN diego_io_oeb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1871.520 0.000 1872.080 4.000 ;
    END
  END diego_io_oeb[30]
  PIN diego_io_oeb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1878.240 0.000 1878.800 4.000 ;
    END
  END diego_io_oeb[31]
  PIN diego_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1690.080 0.000 1690.640 4.000 ;
    END
  END diego_io_oeb[3]
  PIN diego_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1696.800 0.000 1697.360 4.000 ;
    END
  END diego_io_oeb[4]
  PIN diego_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1703.520 0.000 1704.080 4.000 ;
    END
  END diego_io_oeb[5]
  PIN diego_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1710.240 0.000 1710.800 4.000 ;
    END
  END diego_io_oeb[6]
  PIN diego_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1716.960 0.000 1717.520 4.000 ;
    END
  END diego_io_oeb[7]
  PIN diego_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1723.680 0.000 1724.240 4.000 ;
    END
  END diego_io_oeb[8]
  PIN diego_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1730.400 0.000 1730.960 4.000 ;
    END
  END diego_io_oeb[9]
  PIN diego_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1454.880 0.000 1455.440 4.000 ;
    END
  END diego_io_out[0]
  PIN diego_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1522.080 0.000 1522.640 4.000 ;
    END
  END diego_io_out[10]
  PIN diego_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1528.800 0.000 1529.360 4.000 ;
    END
  END diego_io_out[11]
  PIN diego_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1535.520 0.000 1536.080 4.000 ;
    END
  END diego_io_out[12]
  PIN diego_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1542.240 0.000 1542.800 4.000 ;
    END
  END diego_io_out[13]
  PIN diego_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1548.960 0.000 1549.520 4.000 ;
    END
  END diego_io_out[14]
  PIN diego_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1555.680 0.000 1556.240 4.000 ;
    END
  END diego_io_out[15]
  PIN diego_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1562.400 0.000 1562.960 4.000 ;
    END
  END diego_io_out[16]
  PIN diego_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1569.120 0.000 1569.680 4.000 ;
    END
  END diego_io_out[17]
  PIN diego_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1575.840 0.000 1576.400 4.000 ;
    END
  END diego_io_out[18]
  PIN diego_io_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1582.560 0.000 1583.120 4.000 ;
    END
  END diego_io_out[19]
  PIN diego_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1461.600 0.000 1462.160 4.000 ;
    END
  END diego_io_out[1]
  PIN diego_io_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1589.280 0.000 1589.840 4.000 ;
    END
  END diego_io_out[20]
  PIN diego_io_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1596.000 0.000 1596.560 4.000 ;
    END
  END diego_io_out[21]
  PIN diego_io_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1602.720 0.000 1603.280 4.000 ;
    END
  END diego_io_out[22]
  PIN diego_io_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1609.440 0.000 1610.000 4.000 ;
    END
  END diego_io_out[23]
  PIN diego_io_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1616.160 0.000 1616.720 4.000 ;
    END
  END diego_io_out[24]
  PIN diego_io_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1622.880 0.000 1623.440 4.000 ;
    END
  END diego_io_out[25]
  PIN diego_io_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1629.600 0.000 1630.160 4.000 ;
    END
  END diego_io_out[26]
  PIN diego_io_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1636.320 0.000 1636.880 4.000 ;
    END
  END diego_io_out[27]
  PIN diego_io_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1643.040 0.000 1643.600 4.000 ;
    END
  END diego_io_out[28]
  PIN diego_io_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1649.760 0.000 1650.320 4.000 ;
    END
  END diego_io_out[29]
  PIN diego_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1468.320 0.000 1468.880 4.000 ;
    END
  END diego_io_out[2]
  PIN diego_io_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1656.480 0.000 1657.040 4.000 ;
    END
  END diego_io_out[30]
  PIN diego_io_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1663.200 0.000 1663.760 4.000 ;
    END
  END diego_io_out[31]
  PIN diego_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1475.040 0.000 1475.600 4.000 ;
    END
  END diego_io_out[3]
  PIN diego_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1481.760 0.000 1482.320 4.000 ;
    END
  END diego_io_out[4]
  PIN diego_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1488.480 0.000 1489.040 4.000 ;
    END
  END diego_io_out[5]
  PIN diego_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1495.200 0.000 1495.760 4.000 ;
    END
  END diego_io_out[6]
  PIN diego_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1501.920 0.000 1502.480 4.000 ;
    END
  END diego_io_out[7]
  PIN diego_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1508.640 0.000 1509.200 4.000 ;
    END
  END diego_io_out[8]
  PIN diego_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1515.360 0.000 1515.920 4.000 ;
    END
  END diego_io_out[9]
  PIN diego_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1441.440 0.000 1442.000 4.000 ;
    END
  END diego_rst
  PIN i_design_reset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 39.200 2400.000 39.760 ;
    END
  END i_design_reset[0]
  PIN i_design_reset[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 43.680 2400.000 44.240 ;
    END
  END i_design_reset[1]
  PIN i_design_reset[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 48.160 2400.000 48.720 ;
    END
  END i_design_reset[2]
  PIN i_design_reset[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 52.640 2400.000 53.200 ;
    END
  END i_design_reset[3]
  PIN i_design_reset[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 57.120 2400.000 57.680 ;
    END
  END i_design_reset[4]
  PIN i_design_reset[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 61.600 2400.000 62.160 ;
    END
  END i_design_reset[5]
  PIN i_design_reset[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 66.080 2400.000 66.640 ;
    END
  END i_design_reset[6]
  PIN i_design_reset[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 70.560 2400.000 71.120 ;
    END
  END i_design_reset[7]
  PIN i_mux_auto_reset_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 34.720 2400.000 35.280 ;
    END
  END i_mux_auto_reset_enb
  PIN i_mux_io5_reset_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 7.840 2400.000 8.400 ;
    END
  END i_mux_io5_reset_enb
  PIN i_mux_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 12.320 2400.000 12.880 ;
    END
  END i_mux_sel[0]
  PIN i_mux_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 16.800 2400.000 17.360 ;
    END
  END i_mux_sel[1]
  PIN i_mux_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 21.280 2400.000 21.840 ;
    END
  END i_mux_sel[2]
  PIN i_mux_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 25.760 2400.000 26.320 ;
    END
  END i_mux_sel[3]
  PIN i_mux_sys_reset_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 30.240 2400.000 30.800 ;
    END
  END i_mux_sys_reset_enb
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 79.520 2400.000 80.080 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 213.920 2400.000 214.480 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 227.360 2400.000 227.920 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 240.800 2400.000 241.360 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 254.240 2400.000 254.800 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 267.680 2400.000 268.240 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 281.120 2400.000 281.680 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1962.240 296.000 1962.800 300.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1942.080 296.000 1942.640 300.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1921.920 296.000 1922.480 300.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 296.000 638.960 300.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 92.960 2400.000 93.520 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 296.000 618.800 300.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 296.000 598.640 300.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 296.000 578.480 300.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 277.760 4.000 278.320 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 4.000 261.520 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.160 4.000 244.720 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 227.360 4.000 227.920 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 210.560 4.000 211.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 193.760 4.000 194.320 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.960 4.000 177.520 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 106.400 2400.000 106.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.160 4.000 160.720 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 143.360 4.000 143.920 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.560 4.000 127.120 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.760 4.000 110.320 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.960 4.000 93.520 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 76.160 4.000 76.720 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 4.000 59.920 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 4.000 43.120 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 119.840 2400.000 120.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 133.280 2400.000 133.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 146.720 2400.000 147.280 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 160.160 2400.000 160.720 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 173.600 2400.000 174.160 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 187.040 2400.000 187.600 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 200.480 2400.000 201.040 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 88.480 2400.000 89.040 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 222.880 2400.000 223.440 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 236.320 2400.000 236.880 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 249.760 2400.000 250.320 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 263.200 2400.000 263.760 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 276.640 2400.000 277.200 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 290.080 2400.000 290.640 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1948.800 296.000 1949.360 300.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1928.640 296.000 1929.200 300.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1908.480 296.000 1909.040 300.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 296.000 625.520 300.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 101.920 2400.000 102.480 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 296.000 605.360 300.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 296.000 585.200 300.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 296.000 565.040 300.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 266.560 4.000 267.120 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 249.760 4.000 250.320 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.960 4.000 233.520 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.160 4.000 216.720 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.360 4.000 199.920 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.560 4.000 183.120 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 165.760 4.000 166.320 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 115.360 2400.000 115.920 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.960 4.000 149.520 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.160 4.000 132.720 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 98.560 4.000 99.120 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.760 4.000 82.320 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.960 4.000 65.520 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 4.000 48.720 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.360 4.000 31.920 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 128.800 2400.000 129.360 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 142.240 2400.000 142.800 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 155.680 2400.000 156.240 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 169.120 2400.000 169.680 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 182.560 2400.000 183.120 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 196.000 2400.000 196.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 209.440 2400.000 210.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 84.000 2400.000 84.560 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 218.400 2400.000 218.960 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 231.840 2400.000 232.400 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 245.280 2400.000 245.840 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 258.720 2400.000 259.280 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 272.160 2400.000 272.720 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 285.600 2400.000 286.160 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1955.520 296.000 1956.080 300.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1935.360 296.000 1935.920 300.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1915.200 296.000 1915.760 300.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 296.000 632.240 300.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 97.440 2400.000 98.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 296.000 612.080 300.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 296.000 591.920 300.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 296.000 571.760 300.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 4.000 272.720 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.360 4.000 255.920 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 4.000 171.920 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 110.880 2400.000 111.440 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 4.000 71.120 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.960 4.000 37.520 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 124.320 2400.000 124.880 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 137.760 2400.000 138.320 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 151.200 2400.000 151.760 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 164.640 2400.000 165.200 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 178.080 2400.000 178.640 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 191.520 2400.000 192.080 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 204.960 2400.000 205.520 ;
    END
  END io_out[9]
  PIN la_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1125.600 0.000 1126.160 4.000 ;
    END
  END la_in[0]
  PIN la_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1192.800 0.000 1193.360 4.000 ;
    END
  END la_in[10]
  PIN la_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1199.520 0.000 1200.080 4.000 ;
    END
  END la_in[11]
  PIN la_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1206.240 0.000 1206.800 4.000 ;
    END
  END la_in[12]
  PIN la_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1212.960 0.000 1213.520 4.000 ;
    END
  END la_in[13]
  PIN la_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1219.680 0.000 1220.240 4.000 ;
    END
  END la_in[14]
  PIN la_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1226.400 0.000 1226.960 4.000 ;
    END
  END la_in[15]
  PIN la_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1132.320 0.000 1132.880 4.000 ;
    END
  END la_in[1]
  PIN la_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1139.040 0.000 1139.600 4.000 ;
    END
  END la_in[2]
  PIN la_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1145.760 0.000 1146.320 4.000 ;
    END
  END la_in[3]
  PIN la_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1152.480 0.000 1153.040 4.000 ;
    END
  END la_in[4]
  PIN la_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1159.200 0.000 1159.760 4.000 ;
    END
  END la_in[5]
  PIN la_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 0.000 1166.480 4.000 ;
    END
  END la_in[6]
  PIN la_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1172.640 0.000 1173.200 4.000 ;
    END
  END la_in[7]
  PIN la_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1179.360 0.000 1179.920 4.000 ;
    END
  END la_in[8]
  PIN la_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1186.080 0.000 1186.640 4.000 ;
    END
  END la_in[9]
  PIN mux_conf_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2396.000 75.040 2400.000 75.600 ;
    END
  END mux_conf_clk
  PIN pawel_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END pawel_clk
  PIN pawel_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END pawel_ena
  PIN pawel_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END pawel_io_in[0]
  PIN pawel_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 4.000 ;
    END
  END pawel_io_in[10]
  PIN pawel_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END pawel_io_in[11]
  PIN pawel_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 0.000 306.320 4.000 ;
    END
  END pawel_io_in[12]
  PIN pawel_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 0.000 326.480 4.000 ;
    END
  END pawel_io_in[13]
  PIN pawel_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 0.000 333.200 4.000 ;
    END
  END pawel_io_in[14]
  PIN pawel_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 0.000 339.920 4.000 ;
    END
  END pawel_io_in[15]
  PIN pawel_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 0.000 346.640 4.000 ;
    END
  END pawel_io_in[16]
  PIN pawel_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END pawel_io_in[17]
  PIN pawel_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 0.000 360.080 4.000 ;
    END
  END pawel_io_in[18]
  PIN pawel_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END pawel_io_in[19]
  PIN pawel_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END pawel_io_in[1]
  PIN pawel_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 0.000 373.520 4.000 ;
    END
  END pawel_io_in[20]
  PIN pawel_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 0.000 380.240 4.000 ;
    END
  END pawel_io_in[21]
  PIN pawel_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END pawel_io_in[22]
  PIN pawel_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 0.000 393.680 4.000 ;
    END
  END pawel_io_in[23]
  PIN pawel_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 0.000 400.400 4.000 ;
    END
  END pawel_io_in[24]
  PIN pawel_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 0.000 407.120 4.000 ;
    END
  END pawel_io_in[25]
  PIN pawel_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 0.000 413.840 4.000 ;
    END
  END pawel_io_in[26]
  PIN pawel_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 0.000 420.560 4.000 ;
    END
  END pawel_io_in[27]
  PIN pawel_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 0.000 427.280 4.000 ;
    END
  END pawel_io_in[28]
  PIN pawel_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 0.000 434.000 4.000 ;
    END
  END pawel_io_in[29]
  PIN pawel_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END pawel_io_in[2]
  PIN pawel_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 0.000 440.720 4.000 ;
    END
  END pawel_io_in[30]
  PIN pawel_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 0.000 447.440 4.000 ;
    END
  END pawel_io_in[31]
  PIN pawel_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 0.000 454.160 4.000 ;
    END
  END pawel_io_in[32]
  PIN pawel_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 0.000 460.880 4.000 ;
    END
  END pawel_io_in[33]
  PIN pawel_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 0.000 467.600 4.000 ;
    END
  END pawel_io_in[34]
  PIN pawel_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 0.000 474.320 4.000 ;
    END
  END pawel_io_in[35]
  PIN pawel_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 0.000 481.040 4.000 ;
    END
  END pawel_io_in[36]
  PIN pawel_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 0.000 487.760 4.000 ;
    END
  END pawel_io_in[37]
  PIN pawel_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END pawel_io_in[3]
  PIN pawel_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END pawel_io_in[4]
  PIN pawel_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END pawel_io_in[5]
  PIN pawel_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END pawel_io_in[6]
  PIN pawel_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END pawel_io_in[7]
  PIN pawel_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END pawel_io_in[8]
  PIN pawel_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 4.000 ;
    END
  END pawel_io_in[9]
  PIN pawel_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END pawel_io_oeb[0]
  PIN pawel_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 0.000 272.720 4.000 ;
    END
  END pawel_io_oeb[10]
  PIN pawel_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 0.000 292.880 4.000 ;
    END
  END pawel_io_oeb[11]
  PIN pawel_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END pawel_io_oeb[12]
  PIN pawel_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END pawel_io_oeb[1]
  PIN pawel_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END pawel_io_oeb[2]
  PIN pawel_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END pawel_io_oeb[3]
  PIN pawel_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END pawel_io_oeb[4]
  PIN pawel_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END pawel_io_oeb[5]
  PIN pawel_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END pawel_io_oeb[6]
  PIN pawel_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END pawel_io_oeb[7]
  PIN pawel_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 0.000 232.400 4.000 ;
    END
  END pawel_io_oeb[8]
  PIN pawel_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 4.000 ;
    END
  END pawel_io_oeb[9]
  PIN pawel_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END pawel_io_out[0]
  PIN pawel_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 4.000 ;
    END
  END pawel_io_out[10]
  PIN pawel_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 0.000 299.600 4.000 ;
    END
  END pawel_io_out[11]
  PIN pawel_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 0.000 319.760 4.000 ;
    END
  END pawel_io_out[12]
  PIN pawel_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END pawel_io_out[1]
  PIN pawel_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END pawel_io_out[2]
  PIN pawel_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END pawel_io_out[3]
  PIN pawel_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END pawel_io_out[4]
  PIN pawel_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END pawel_io_out[5]
  PIN pawel_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 4.000 ;
    END
  END pawel_io_out[6]
  PIN pawel_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END pawel_io_out[7]
  PIN pawel_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END pawel_io_out[8]
  PIN pawel_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 0.000 259.280 4.000 ;
    END
  END pawel_io_out[9]
  PIN pawel_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END pawel_rst
  PIN solos_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2002.560 296.000 2003.120 300.000 ;
    END
  END solos_clk
  PIN solos_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2016.000 296.000 2016.560 300.000 ;
    END
  END solos_ena
  PIN solos_gpio_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2022.720 296.000 2023.280 300.000 ;
    END
  END solos_gpio_ready
  PIN solos_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2365.440 296.000 2366.000 300.000 ;
    END
  END solos_io_in[0]
  PIN solos_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2298.240 296.000 2298.800 300.000 ;
    END
  END solos_io_in[10]
  PIN solos_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2291.520 296.000 2292.080 300.000 ;
    END
  END solos_io_in[11]
  PIN solos_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2284.800 296.000 2285.360 300.000 ;
    END
  END solos_io_in[12]
  PIN solos_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2278.080 296.000 2278.640 300.000 ;
    END
  END solos_io_in[13]
  PIN solos_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2271.360 296.000 2271.920 300.000 ;
    END
  END solos_io_in[14]
  PIN solos_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2264.640 296.000 2265.200 300.000 ;
    END
  END solos_io_in[15]
  PIN solos_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2257.920 296.000 2258.480 300.000 ;
    END
  END solos_io_in[16]
  PIN solos_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2251.200 296.000 2251.760 300.000 ;
    END
  END solos_io_in[17]
  PIN solos_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2244.480 296.000 2245.040 300.000 ;
    END
  END solos_io_in[18]
  PIN solos_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2237.760 296.000 2238.320 300.000 ;
    END
  END solos_io_in[19]
  PIN solos_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2358.720 296.000 2359.280 300.000 ;
    END
  END solos_io_in[1]
  PIN solos_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2231.040 296.000 2231.600 300.000 ;
    END
  END solos_io_in[20]
  PIN solos_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2224.320 296.000 2224.880 300.000 ;
    END
  END solos_io_in[21]
  PIN solos_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2217.600 296.000 2218.160 300.000 ;
    END
  END solos_io_in[22]
  PIN solos_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2210.880 296.000 2211.440 300.000 ;
    END
  END solos_io_in[23]
  PIN solos_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2204.160 296.000 2204.720 300.000 ;
    END
  END solos_io_in[24]
  PIN solos_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2197.440 296.000 2198.000 300.000 ;
    END
  END solos_io_in[25]
  PIN solos_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2190.720 296.000 2191.280 300.000 ;
    END
  END solos_io_in[26]
  PIN solos_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2184.000 296.000 2184.560 300.000 ;
    END
  END solos_io_in[27]
  PIN solos_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2177.280 296.000 2177.840 300.000 ;
    END
  END solos_io_in[28]
  PIN solos_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2170.560 296.000 2171.120 300.000 ;
    END
  END solos_io_in[29]
  PIN solos_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2352.000 296.000 2352.560 300.000 ;
    END
  END solos_io_in[2]
  PIN solos_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2163.840 296.000 2164.400 300.000 ;
    END
  END solos_io_in[30]
  PIN solos_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2157.120 296.000 2157.680 300.000 ;
    END
  END solos_io_in[31]
  PIN solos_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2150.400 296.000 2150.960 300.000 ;
    END
  END solos_io_in[32]
  PIN solos_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2143.680 296.000 2144.240 300.000 ;
    END
  END solos_io_in[33]
  PIN solos_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2136.960 296.000 2137.520 300.000 ;
    END
  END solos_io_in[34]
  PIN solos_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2130.240 296.000 2130.800 300.000 ;
    END
  END solos_io_in[35]
  PIN solos_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2123.520 296.000 2124.080 300.000 ;
    END
  END solos_io_in[36]
  PIN solos_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2116.800 296.000 2117.360 300.000 ;
    END
  END solos_io_in[37]
  PIN solos_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2345.280 296.000 2345.840 300.000 ;
    END
  END solos_io_in[3]
  PIN solos_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2338.560 296.000 2339.120 300.000 ;
    END
  END solos_io_in[4]
  PIN solos_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2331.840 296.000 2332.400 300.000 ;
    END
  END solos_io_in[5]
  PIN solos_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2325.120 296.000 2325.680 300.000 ;
    END
  END solos_io_in[6]
  PIN solos_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2318.400 296.000 2318.960 300.000 ;
    END
  END solos_io_in[7]
  PIN solos_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2311.680 296.000 2312.240 300.000 ;
    END
  END solos_io_in[8]
  PIN solos_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2304.960 296.000 2305.520 300.000 ;
    END
  END solos_io_in[9]
  PIN solos_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2110.080 296.000 2110.640 300.000 ;
    END
  END solos_io_out[0]
  PIN solos_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2042.880 296.000 2043.440 300.000 ;
    END
  END solos_io_out[10]
  PIN solos_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2036.160 296.000 2036.720 300.000 ;
    END
  END solos_io_out[11]
  PIN solos_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2029.440 296.000 2030.000 300.000 ;
    END
  END solos_io_out[12]
  PIN solos_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2103.360 296.000 2103.920 300.000 ;
    END
  END solos_io_out[1]
  PIN solos_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2096.640 296.000 2097.200 300.000 ;
    END
  END solos_io_out[2]
  PIN solos_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2089.920 296.000 2090.480 300.000 ;
    END
  END solos_io_out[3]
  PIN solos_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2083.200 296.000 2083.760 300.000 ;
    END
  END solos_io_out[4]
  PIN solos_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2076.480 296.000 2077.040 300.000 ;
    END
  END solos_io_out[5]
  PIN solos_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2069.760 296.000 2070.320 300.000 ;
    END
  END solos_io_out[6]
  PIN solos_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2063.040 296.000 2063.600 300.000 ;
    END
  END solos_io_out[7]
  PIN solos_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2056.320 296.000 2056.880 300.000 ;
    END
  END solos_io_out[8]
  PIN solos_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2049.600 296.000 2050.160 300.000 ;
    END
  END solos_io_out[9]
  PIN solos_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2009.280 296.000 2009.840 300.000 ;
    END
  END solos_rst
  PIN trzf2_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 296.000 719.600 300.000 ;
    END
  END trzf2_clk
  PIN trzf2_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 296.000 712.880 300.000 ;
    END
  END trzf2_ena
  PIN trzf2_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1169.280 296.000 1169.840 300.000 ;
    END
  END trzf2_io_in[0]
  PIN trzf2_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1102.080 296.000 1102.640 300.000 ;
    END
  END trzf2_io_in[10]
  PIN trzf2_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1095.360 296.000 1095.920 300.000 ;
    END
  END trzf2_io_in[11]
  PIN trzf2_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1088.640 296.000 1089.200 300.000 ;
    END
  END trzf2_io_in[12]
  PIN trzf2_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1081.920 296.000 1082.480 300.000 ;
    END
  END trzf2_io_in[13]
  PIN trzf2_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1075.200 296.000 1075.760 300.000 ;
    END
  END trzf2_io_in[14]
  PIN trzf2_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1068.480 296.000 1069.040 300.000 ;
    END
  END trzf2_io_in[15]
  PIN trzf2_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1061.760 296.000 1062.320 300.000 ;
    END
  END trzf2_io_in[16]
  PIN trzf2_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 296.000 1055.600 300.000 ;
    END
  END trzf2_io_in[17]
  PIN trzf2_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1048.320 296.000 1048.880 300.000 ;
    END
  END trzf2_io_in[18]
  PIN trzf2_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1041.600 296.000 1042.160 300.000 ;
    END
  END trzf2_io_in[19]
  PIN trzf2_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1162.560 296.000 1163.120 300.000 ;
    END
  END trzf2_io_in[1]
  PIN trzf2_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1034.880 296.000 1035.440 300.000 ;
    END
  END trzf2_io_in[20]
  PIN trzf2_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1028.160 296.000 1028.720 300.000 ;
    END
  END trzf2_io_in[21]
  PIN trzf2_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1021.440 296.000 1022.000 300.000 ;
    END
  END trzf2_io_in[22]
  PIN trzf2_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1014.720 296.000 1015.280 300.000 ;
    END
  END trzf2_io_in[23]
  PIN trzf2_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1008.000 296.000 1008.560 300.000 ;
    END
  END trzf2_io_in[24]
  PIN trzf2_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1001.280 296.000 1001.840 300.000 ;
    END
  END trzf2_io_in[25]
  PIN trzf2_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 296.000 995.120 300.000 ;
    END
  END trzf2_io_in[26]
  PIN trzf2_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 987.840 296.000 988.400 300.000 ;
    END
  END trzf2_io_in[27]
  PIN trzf2_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 296.000 981.680 300.000 ;
    END
  END trzf2_io_in[28]
  PIN trzf2_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 296.000 974.960 300.000 ;
    END
  END trzf2_io_in[29]
  PIN trzf2_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1155.840 296.000 1156.400 300.000 ;
    END
  END trzf2_io_in[2]
  PIN trzf2_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 967.680 296.000 968.240 300.000 ;
    END
  END trzf2_io_in[30]
  PIN trzf2_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 296.000 961.520 300.000 ;
    END
  END trzf2_io_in[31]
  PIN trzf2_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 296.000 954.800 300.000 ;
    END
  END trzf2_io_in[32]
  PIN trzf2_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 296.000 948.080 300.000 ;
    END
  END trzf2_io_in[33]
  PIN trzf2_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 940.800 296.000 941.360 300.000 ;
    END
  END trzf2_io_in[34]
  PIN trzf2_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 296.000 934.640 300.000 ;
    END
  END trzf2_io_in[35]
  PIN trzf2_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 296.000 927.920 300.000 ;
    END
  END trzf2_io_in[36]
  PIN trzf2_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 920.640 296.000 921.200 300.000 ;
    END
  END trzf2_io_in[37]
  PIN trzf2_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1149.120 296.000 1149.680 300.000 ;
    END
  END trzf2_io_in[3]
  PIN trzf2_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1142.400 296.000 1142.960 300.000 ;
    END
  END trzf2_io_in[4]
  PIN trzf2_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1135.680 296.000 1136.240 300.000 ;
    END
  END trzf2_io_in[5]
  PIN trzf2_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1128.960 296.000 1129.520 300.000 ;
    END
  END trzf2_io_in[6]
  PIN trzf2_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1122.240 296.000 1122.800 300.000 ;
    END
  END trzf2_io_in[7]
  PIN trzf2_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1115.520 296.000 1116.080 300.000 ;
    END
  END trzf2_io_in[8]
  PIN trzf2_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1108.800 296.000 1109.360 300.000 ;
    END
  END trzf2_io_in[9]
  PIN trzf2_la_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 296.000 813.680 300.000 ;
    END
  END trzf2_la_in[0]
  PIN trzf2_la_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 296.000 746.480 300.000 ;
    END
  END trzf2_la_in[10]
  PIN trzf2_la_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 296.000 739.760 300.000 ;
    END
  END trzf2_la_in[11]
  PIN trzf2_la_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 296.000 733.040 300.000 ;
    END
  END trzf2_la_in[12]
  PIN trzf2_la_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 806.400 296.000 806.960 300.000 ;
    END
  END trzf2_la_in[1]
  PIN trzf2_la_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 296.000 800.240 300.000 ;
    END
  END trzf2_la_in[2]
  PIN trzf2_la_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 792.960 296.000 793.520 300.000 ;
    END
  END trzf2_la_in[3]
  PIN trzf2_la_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 786.240 296.000 786.800 300.000 ;
    END
  END trzf2_la_in[4]
  PIN trzf2_la_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 296.000 780.080 300.000 ;
    END
  END trzf2_la_in[5]
  PIN trzf2_la_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 296.000 773.360 300.000 ;
    END
  END trzf2_la_in[6]
  PIN trzf2_la_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 766.080 296.000 766.640 300.000 ;
    END
  END trzf2_la_in[7]
  PIN trzf2_la_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 296.000 759.920 300.000 ;
    END
  END trzf2_la_in[8]
  PIN trzf2_la_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 296.000 753.200 300.000 ;
    END
  END trzf2_la_in[9]
  PIN trzf2_o_gpout[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 833.280 296.000 833.840 300.000 ;
    END
  END trzf2_o_gpout[0]
  PIN trzf2_o_gpout[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 826.560 296.000 827.120 300.000 ;
    END
  END trzf2_o_gpout[1]
  PIN trzf2_o_gpout[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 819.840 296.000 820.400 300.000 ;
    END
  END trzf2_o_gpout[2]
  PIN trzf2_o_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 913.920 296.000 914.480 300.000 ;
    END
  END trzf2_o_hsync
  PIN trzf2_o_rgb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 900.480 296.000 901.040 300.000 ;
    END
  END trzf2_o_rgb[0]
  PIN trzf2_o_rgb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 893.760 296.000 894.320 300.000 ;
    END
  END trzf2_o_rgb[1]
  PIN trzf2_o_rgb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 887.040 296.000 887.600 300.000 ;
    END
  END trzf2_o_rgb[2]
  PIN trzf2_o_rgb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 880.320 296.000 880.880 300.000 ;
    END
  END trzf2_o_rgb[3]
  PIN trzf2_o_rgb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 873.600 296.000 874.160 300.000 ;
    END
  END trzf2_o_rgb[4]
  PIN trzf2_o_rgb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 866.880 296.000 867.440 300.000 ;
    END
  END trzf2_o_rgb[5]
  PIN trzf2_o_tex_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 860.160 296.000 860.720 300.000 ;
    END
  END trzf2_o_tex_csb
  PIN trzf2_o_tex_oeb0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 296.000 840.560 300.000 ;
    END
  END trzf2_o_tex_oeb0
  PIN trzf2_o_tex_out0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 846.720 296.000 847.280 300.000 ;
    END
  END trzf2_o_tex_out0
  PIN trzf2_o_tex_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 296.000 854.000 300.000 ;
    END
  END trzf2_o_tex_sclk
  PIN trzf2_o_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 296.000 907.760 300.000 ;
    END
  END trzf2_o_vsync
  PIN trzf2_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 296.000 726.320 300.000 ;
    END
  END trzf2_rst
  PIN trzf_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 296.000 40.880 300.000 ;
    END
  END trzf_clk
  PIN trzf_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 296.000 34.160 300.000 ;
    END
  END trzf_ena
  PIN trzf_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 296.000 491.120 300.000 ;
    END
  END trzf_io_in[0]
  PIN trzf_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 296.000 423.920 300.000 ;
    END
  END trzf_io_in[10]
  PIN trzf_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 296.000 417.200 300.000 ;
    END
  END trzf_io_in[11]
  PIN trzf_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 296.000 410.480 300.000 ;
    END
  END trzf_io_in[12]
  PIN trzf_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 296.000 403.760 300.000 ;
    END
  END trzf_io_in[13]
  PIN trzf_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 296.000 397.040 300.000 ;
    END
  END trzf_io_in[14]
  PIN trzf_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 296.000 390.320 300.000 ;
    END
  END trzf_io_in[15]
  PIN trzf_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 296.000 383.600 300.000 ;
    END
  END trzf_io_in[16]
  PIN trzf_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 296.000 376.880 300.000 ;
    END
  END trzf_io_in[17]
  PIN trzf_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 296.000 370.160 300.000 ;
    END
  END trzf_io_in[18]
  PIN trzf_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 296.000 363.440 300.000 ;
    END
  END trzf_io_in[19]
  PIN trzf_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 296.000 484.400 300.000 ;
    END
  END trzf_io_in[1]
  PIN trzf_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 296.000 356.720 300.000 ;
    END
  END trzf_io_in[20]
  PIN trzf_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 296.000 350.000 300.000 ;
    END
  END trzf_io_in[21]
  PIN trzf_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 296.000 343.280 300.000 ;
    END
  END trzf_io_in[22]
  PIN trzf_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 296.000 336.560 300.000 ;
    END
  END trzf_io_in[23]
  PIN trzf_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 296.000 329.840 300.000 ;
    END
  END trzf_io_in[24]
  PIN trzf_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 296.000 323.120 300.000 ;
    END
  END trzf_io_in[25]
  PIN trzf_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 296.000 316.400 300.000 ;
    END
  END trzf_io_in[26]
  PIN trzf_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 296.000 309.680 300.000 ;
    END
  END trzf_io_in[27]
  PIN trzf_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 296.000 302.960 300.000 ;
    END
  END trzf_io_in[28]
  PIN trzf_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 296.000 296.240 300.000 ;
    END
  END trzf_io_in[29]
  PIN trzf_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 296.000 477.680 300.000 ;
    END
  END trzf_io_in[2]
  PIN trzf_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 296.000 289.520 300.000 ;
    END
  END trzf_io_in[30]
  PIN trzf_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 296.000 282.800 300.000 ;
    END
  END trzf_io_in[31]
  PIN trzf_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 296.000 276.080 300.000 ;
    END
  END trzf_io_in[32]
  PIN trzf_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 296.000 269.360 300.000 ;
    END
  END trzf_io_in[33]
  PIN trzf_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 296.000 262.640 300.000 ;
    END
  END trzf_io_in[34]
  PIN trzf_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 296.000 255.920 300.000 ;
    END
  END trzf_io_in[35]
  PIN trzf_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 296.000 249.200 300.000 ;
    END
  END trzf_io_in[36]
  PIN trzf_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 296.000 242.480 300.000 ;
    END
  END trzf_io_in[37]
  PIN trzf_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 296.000 470.960 300.000 ;
    END
  END trzf_io_in[3]
  PIN trzf_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 296.000 464.240 300.000 ;
    END
  END trzf_io_in[4]
  PIN trzf_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 296.000 457.520 300.000 ;
    END
  END trzf_io_in[5]
  PIN trzf_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 296.000 450.800 300.000 ;
    END
  END trzf_io_in[6]
  PIN trzf_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 296.000 444.080 300.000 ;
    END
  END trzf_io_in[7]
  PIN trzf_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 296.000 437.360 300.000 ;
    END
  END trzf_io_in[8]
  PIN trzf_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 296.000 430.640 300.000 ;
    END
  END trzf_io_in[9]
  PIN trzf_la_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 296.000 134.960 300.000 ;
    END
  END trzf_la_in[0]
  PIN trzf_la_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 296.000 67.760 300.000 ;
    END
  END trzf_la_in[10]
  PIN trzf_la_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 296.000 61.040 300.000 ;
    END
  END trzf_la_in[11]
  PIN trzf_la_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 296.000 54.320 300.000 ;
    END
  END trzf_la_in[12]
  PIN trzf_la_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 296.000 128.240 300.000 ;
    END
  END trzf_la_in[1]
  PIN trzf_la_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 296.000 121.520 300.000 ;
    END
  END trzf_la_in[2]
  PIN trzf_la_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 296.000 114.800 300.000 ;
    END
  END trzf_la_in[3]
  PIN trzf_la_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 296.000 108.080 300.000 ;
    END
  END trzf_la_in[4]
  PIN trzf_la_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 296.000 101.360 300.000 ;
    END
  END trzf_la_in[5]
  PIN trzf_la_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 296.000 94.640 300.000 ;
    END
  END trzf_la_in[6]
  PIN trzf_la_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 296.000 87.920 300.000 ;
    END
  END trzf_la_in[7]
  PIN trzf_la_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 296.000 81.200 300.000 ;
    END
  END trzf_la_in[8]
  PIN trzf_la_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 296.000 74.480 300.000 ;
    END
  END trzf_la_in[9]
  PIN trzf_o_gpout[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 296.000 155.120 300.000 ;
    END
  END trzf_o_gpout[0]
  PIN trzf_o_gpout[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 296.000 148.400 300.000 ;
    END
  END trzf_o_gpout[1]
  PIN trzf_o_gpout[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 296.000 141.680 300.000 ;
    END
  END trzf_o_gpout[2]
  PIN trzf_o_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 296.000 235.760 300.000 ;
    END
  END trzf_o_hsync
  PIN trzf_o_rgb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 296.000 222.320 300.000 ;
    END
  END trzf_o_rgb[0]
  PIN trzf_o_rgb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 296.000 215.600 300.000 ;
    END
  END trzf_o_rgb[1]
  PIN trzf_o_rgb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 296.000 208.880 300.000 ;
    END
  END trzf_o_rgb[2]
  PIN trzf_o_rgb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 296.000 202.160 300.000 ;
    END
  END trzf_o_rgb[3]
  PIN trzf_o_rgb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 296.000 195.440 300.000 ;
    END
  END trzf_o_rgb[4]
  PIN trzf_o_rgb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 296.000 188.720 300.000 ;
    END
  END trzf_o_rgb[5]
  PIN trzf_o_tex_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 296.000 182.000 300.000 ;
    END
  END trzf_o_tex_csb
  PIN trzf_o_tex_oeb0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 296.000 161.840 300.000 ;
    END
  END trzf_o_tex_oeb0
  PIN trzf_o_tex_out0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 296.000 168.560 300.000 ;
    END
  END trzf_o_tex_out0
  PIN trzf_o_tex_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 296.000 175.280 300.000 ;
    END
  END trzf_o_tex_sclk
  PIN trzf_o_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 296.000 229.040 300.000 ;
    END
  END trzf_o_vsync
  PIN trzf_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 296.000 47.600 300.000 ;
    END
  END trzf_rst
  PIN uri_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 0.000 528.080 4.000 ;
    END
  END uri_clk
  PIN uri_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 0.000 541.520 4.000 ;
    END
  END uri_ena
  PIN uri_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 0.000 548.240 4.000 ;
    END
  END uri_io_in[0]
  PIN uri_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 0.000 749.840 4.000 ;
    END
  END uri_io_in[10]
  PIN uri_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 0.000 770.000 4.000 ;
    END
  END uri_io_in[11]
  PIN uri_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 0.000 790.160 4.000 ;
    END
  END uri_io_in[12]
  PIN uri_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 0.000 810.320 4.000 ;
    END
  END uri_io_in[13]
  PIN uri_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 0.000 830.480 4.000 ;
    END
  END uri_io_in[14]
  PIN uri_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 0.000 850.640 4.000 ;
    END
  END uri_io_in[15]
  PIN uri_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 0.000 870.800 4.000 ;
    END
  END uri_io_in[16]
  PIN uri_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 0.000 890.960 4.000 ;
    END
  END uri_io_in[17]
  PIN uri_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 910.560 0.000 911.120 4.000 ;
    END
  END uri_io_in[18]
  PIN uri_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 930.720 0.000 931.280 4.000 ;
    END
  END uri_io_in[19]
  PIN uri_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 0.000 568.400 4.000 ;
    END
  END uri_io_in[1]
  PIN uri_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 0.000 938.000 4.000 ;
    END
  END uri_io_in[20]
  PIN uri_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 0.000 944.720 4.000 ;
    END
  END uri_io_in[21]
  PIN uri_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 950.880 0.000 951.440 4.000 ;
    END
  END uri_io_in[22]
  PIN uri_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 0.000 958.160 4.000 ;
    END
  END uri_io_in[23]
  PIN uri_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 964.320 0.000 964.880 4.000 ;
    END
  END uri_io_in[24]
  PIN uri_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 0.000 971.600 4.000 ;
    END
  END uri_io_in[25]
  PIN uri_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 977.760 0.000 978.320 4.000 ;
    END
  END uri_io_in[26]
  PIN uri_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 0.000 985.040 4.000 ;
    END
  END uri_io_in[27]
  PIN uri_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 0.000 991.760 4.000 ;
    END
  END uri_io_in[28]
  PIN uri_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 997.920 0.000 998.480 4.000 ;
    END
  END uri_io_in[29]
  PIN uri_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 0.000 588.560 4.000 ;
    END
  END uri_io_in[2]
  PIN uri_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1004.640 0.000 1005.200 4.000 ;
    END
  END uri_io_in[30]
  PIN uri_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1011.360 0.000 1011.920 4.000 ;
    END
  END uri_io_in[31]
  PIN uri_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 0.000 1018.640 4.000 ;
    END
  END uri_io_in[32]
  PIN uri_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1024.800 0.000 1025.360 4.000 ;
    END
  END uri_io_in[33]
  PIN uri_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1031.520 0.000 1032.080 4.000 ;
    END
  END uri_io_in[34]
  PIN uri_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1038.240 0.000 1038.800 4.000 ;
    END
  END uri_io_in[35]
  PIN uri_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1044.960 0.000 1045.520 4.000 ;
    END
  END uri_io_in[36]
  PIN uri_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1051.680 0.000 1052.240 4.000 ;
    END
  END uri_io_in[37]
  PIN uri_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 0.000 608.720 4.000 ;
    END
  END uri_io_in[3]
  PIN uri_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 0.000 628.880 4.000 ;
    END
  END uri_io_in[4]
  PIN uri_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 0.000 649.040 4.000 ;
    END
  END uri_io_in[5]
  PIN uri_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 0.000 669.200 4.000 ;
    END
  END uri_io_in[6]
  PIN uri_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 0.000 689.360 4.000 ;
    END
  END uri_io_in[7]
  PIN uri_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 0.000 709.520 4.000 ;
    END
  END uri_io_in[8]
  PIN uri_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 0.000 729.680 4.000 ;
    END
  END uri_io_in[9]
  PIN uri_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 0.000 554.960 4.000 ;
    END
  END uri_io_oeb[0]
  PIN uri_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 0.000 756.560 4.000 ;
    END
  END uri_io_oeb[10]
  PIN uri_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 0.000 776.720 4.000 ;
    END
  END uri_io_oeb[11]
  PIN uri_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 0.000 796.880 4.000 ;
    END
  END uri_io_oeb[12]
  PIN uri_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 0.000 817.040 4.000 ;
    END
  END uri_io_oeb[13]
  PIN uri_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 0.000 837.200 4.000 ;
    END
  END uri_io_oeb[14]
  PIN uri_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 0.000 857.360 4.000 ;
    END
  END uri_io_oeb[15]
  PIN uri_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 0.000 877.520 4.000 ;
    END
  END uri_io_oeb[16]
  PIN uri_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 0.000 897.680 4.000 ;
    END
  END uri_io_oeb[17]
  PIN uri_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 0.000 917.840 4.000 ;
    END
  END uri_io_oeb[18]
  PIN uri_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 0.000 575.120 4.000 ;
    END
  END uri_io_oeb[1]
  PIN uri_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 0.000 595.280 4.000 ;
    END
  END uri_io_oeb[2]
  PIN uri_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 0.000 615.440 4.000 ;
    END
  END uri_io_oeb[3]
  PIN uri_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 0.000 635.600 4.000 ;
    END
  END uri_io_oeb[4]
  PIN uri_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 0.000 655.760 4.000 ;
    END
  END uri_io_oeb[5]
  PIN uri_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 0.000 675.920 4.000 ;
    END
  END uri_io_oeb[6]
  PIN uri_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 695.520 0.000 696.080 4.000 ;
    END
  END uri_io_oeb[7]
  PIN uri_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 0.000 716.240 4.000 ;
    END
  END uri_io_oeb[8]
  PIN uri_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 0.000 736.400 4.000 ;
    END
  END uri_io_oeb[9]
  PIN uri_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 0.000 561.680 4.000 ;
    END
  END uri_io_out[0]
  PIN uri_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 0.000 763.280 4.000 ;
    END
  END uri_io_out[10]
  PIN uri_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 0.000 783.440 4.000 ;
    END
  END uri_io_out[11]
  PIN uri_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 0.000 803.600 4.000 ;
    END
  END uri_io_out[12]
  PIN uri_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 0.000 823.760 4.000 ;
    END
  END uri_io_out[13]
  PIN uri_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 0.000 843.920 4.000 ;
    END
  END uri_io_out[14]
  PIN uri_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 0.000 864.080 4.000 ;
    END
  END uri_io_out[15]
  PIN uri_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 0.000 884.240 4.000 ;
    END
  END uri_io_out[16]
  PIN uri_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 0.000 904.400 4.000 ;
    END
  END uri_io_out[17]
  PIN uri_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 0.000 924.560 4.000 ;
    END
  END uri_io_out[18]
  PIN uri_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 0.000 581.840 4.000 ;
    END
  END uri_io_out[1]
  PIN uri_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 0.000 602.000 4.000 ;
    END
  END uri_io_out[2]
  PIN uri_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 0.000 622.160 4.000 ;
    END
  END uri_io_out[3]
  PIN uri_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 0.000 642.320 4.000 ;
    END
  END uri_io_out[4]
  PIN uri_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 0.000 662.480 4.000 ;
    END
  END uri_io_out[5]
  PIN uri_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 0.000 682.640 4.000 ;
    END
  END uri_io_out[6]
  PIN uri_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 0.000 702.800 4.000 ;
    END
  END uri_io_out[7]
  PIN uri_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 0.000 722.960 4.000 ;
    END
  END uri_io_out[8]
  PIN uri_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 0.000 743.120 4.000 ;
    END
  END uri_io_out[9]
  PIN uri_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 0.000 534.800 4.000 ;
    END
  END uri_rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 282.540 ;
    END
  END vdd
  PIN vgasp_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1444.800 296.000 1445.360 300.000 ;
    END
  END vgasp_clk
  PIN vgasp_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1706.880 296.000 1707.440 300.000 ;
    END
  END vgasp_io_in[0]
  PIN vgasp_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1639.680 296.000 1640.240 300.000 ;
    END
  END vgasp_io_in[10]
  PIN vgasp_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1632.960 296.000 1633.520 300.000 ;
    END
  END vgasp_io_in[11]
  PIN vgasp_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1626.240 296.000 1626.800 300.000 ;
    END
  END vgasp_io_in[12]
  PIN vgasp_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1619.520 296.000 1620.080 300.000 ;
    END
  END vgasp_io_in[13]
  PIN vgasp_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1612.800 296.000 1613.360 300.000 ;
    END
  END vgasp_io_in[14]
  PIN vgasp_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1606.080 296.000 1606.640 300.000 ;
    END
  END vgasp_io_in[15]
  PIN vgasp_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1599.360 296.000 1599.920 300.000 ;
    END
  END vgasp_io_in[16]
  PIN vgasp_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1592.640 296.000 1593.200 300.000 ;
    END
  END vgasp_io_in[17]
  PIN vgasp_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1585.920 296.000 1586.480 300.000 ;
    END
  END vgasp_io_in[18]
  PIN vgasp_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1579.200 296.000 1579.760 300.000 ;
    END
  END vgasp_io_in[19]
  PIN vgasp_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1700.160 296.000 1700.720 300.000 ;
    END
  END vgasp_io_in[1]
  PIN vgasp_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1572.480 296.000 1573.040 300.000 ;
    END
  END vgasp_io_in[20]
  PIN vgasp_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1565.760 296.000 1566.320 300.000 ;
    END
  END vgasp_io_in[21]
  PIN vgasp_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1559.040 296.000 1559.600 300.000 ;
    END
  END vgasp_io_in[22]
  PIN vgasp_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1552.320 296.000 1552.880 300.000 ;
    END
  END vgasp_io_in[23]
  PIN vgasp_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1545.600 296.000 1546.160 300.000 ;
    END
  END vgasp_io_in[24]
  PIN vgasp_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1538.880 296.000 1539.440 300.000 ;
    END
  END vgasp_io_in[25]
  PIN vgasp_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1532.160 296.000 1532.720 300.000 ;
    END
  END vgasp_io_in[26]
  PIN vgasp_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1525.440 296.000 1526.000 300.000 ;
    END
  END vgasp_io_in[27]
  PIN vgasp_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1518.720 296.000 1519.280 300.000 ;
    END
  END vgasp_io_in[28]
  PIN vgasp_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1512.000 296.000 1512.560 300.000 ;
    END
  END vgasp_io_in[29]
  PIN vgasp_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1693.440 296.000 1694.000 300.000 ;
    END
  END vgasp_io_in[2]
  PIN vgasp_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1505.280 296.000 1505.840 300.000 ;
    END
  END vgasp_io_in[30]
  PIN vgasp_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1498.560 296.000 1499.120 300.000 ;
    END
  END vgasp_io_in[31]
  PIN vgasp_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1491.840 296.000 1492.400 300.000 ;
    END
  END vgasp_io_in[32]
  PIN vgasp_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1485.120 296.000 1485.680 300.000 ;
    END
  END vgasp_io_in[33]
  PIN vgasp_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1478.400 296.000 1478.960 300.000 ;
    END
  END vgasp_io_in[34]
  PIN vgasp_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1471.680 296.000 1472.240 300.000 ;
    END
  END vgasp_io_in[35]
  PIN vgasp_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1464.960 296.000 1465.520 300.000 ;
    END
  END vgasp_io_in[36]
  PIN vgasp_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1458.240 296.000 1458.800 300.000 ;
    END
  END vgasp_io_in[37]
  PIN vgasp_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1686.720 296.000 1687.280 300.000 ;
    END
  END vgasp_io_in[3]
  PIN vgasp_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1680.000 296.000 1680.560 300.000 ;
    END
  END vgasp_io_in[4]
  PIN vgasp_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1673.280 296.000 1673.840 300.000 ;
    END
  END vgasp_io_in[5]
  PIN vgasp_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1666.560 296.000 1667.120 300.000 ;
    END
  END vgasp_io_in[6]
  PIN vgasp_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1659.840 296.000 1660.400 300.000 ;
    END
  END vgasp_io_in[7]
  PIN vgasp_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1653.120 296.000 1653.680 300.000 ;
    END
  END vgasp_io_in[8]
  PIN vgasp_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1646.400 296.000 1646.960 300.000 ;
    END
  END vgasp_io_in[9]
  PIN vgasp_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1451.520 296.000 1452.080 300.000 ;
    END
  END vgasp_rst
  PIN vgasp_uio_oe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1868.160 296.000 1868.720 300.000 ;
    END
  END vgasp_uio_oe[0]
  PIN vgasp_uio_oe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1861.440 296.000 1862.000 300.000 ;
    END
  END vgasp_uio_oe[1]
  PIN vgasp_uio_oe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1854.720 296.000 1855.280 300.000 ;
    END
  END vgasp_uio_oe[2]
  PIN vgasp_uio_oe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1848.000 296.000 1848.560 300.000 ;
    END
  END vgasp_uio_oe[3]
  PIN vgasp_uio_oe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1841.280 296.000 1841.840 300.000 ;
    END
  END vgasp_uio_oe[4]
  PIN vgasp_uio_oe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1834.560 296.000 1835.120 300.000 ;
    END
  END vgasp_uio_oe[5]
  PIN vgasp_uio_oe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1827.840 296.000 1828.400 300.000 ;
    END
  END vgasp_uio_oe[6]
  PIN vgasp_uio_oe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1821.120 296.000 1821.680 300.000 ;
    END
  END vgasp_uio_oe[7]
  PIN vgasp_uio_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1814.400 296.000 1814.960 300.000 ;
    END
  END vgasp_uio_out[0]
  PIN vgasp_uio_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1807.680 296.000 1808.240 300.000 ;
    END
  END vgasp_uio_out[1]
  PIN vgasp_uio_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1800.960 296.000 1801.520 300.000 ;
    END
  END vgasp_uio_out[2]
  PIN vgasp_uio_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1794.240 296.000 1794.800 300.000 ;
    END
  END vgasp_uio_out[3]
  PIN vgasp_uio_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1787.520 296.000 1788.080 300.000 ;
    END
  END vgasp_uio_out[4]
  PIN vgasp_uio_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1780.800 296.000 1781.360 300.000 ;
    END
  END vgasp_uio_out[5]
  PIN vgasp_uio_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1774.080 296.000 1774.640 300.000 ;
    END
  END vgasp_uio_out[6]
  PIN vgasp_uio_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1767.360 296.000 1767.920 300.000 ;
    END
  END vgasp_uio_out[7]
  PIN vgasp_uo_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1760.640 296.000 1761.200 300.000 ;
    END
  END vgasp_uo_out[0]
  PIN vgasp_uo_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1753.920 296.000 1754.480 300.000 ;
    END
  END vgasp_uo_out[1]
  PIN vgasp_uo_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1747.200 296.000 1747.760 300.000 ;
    END
  END vgasp_uo_out[2]
  PIN vgasp_uo_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1740.480 296.000 1741.040 300.000 ;
    END
  END vgasp_uo_out[3]
  PIN vgasp_uo_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1733.760 296.000 1734.320 300.000 ;
    END
  END vgasp_uo_out[4]
  PIN vgasp_uo_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1727.040 296.000 1727.600 300.000 ;
    END
  END vgasp_uo_out[5]
  PIN vgasp_uo_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1720.320 296.000 1720.880 300.000 ;
    END
  END vgasp_uo_out[6]
  PIN vgasp_uo_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1713.600 296.000 1714.160 300.000 ;
    END
  END vgasp_uo_out[7]
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 282.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.760 4.000 26.320 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END wb_rst_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 4.630 2392.880 285.450 ;
      LAYER Metal2 ;
        RECT 8.540 295.700 33.300 296.660 ;
        RECT 34.460 295.700 40.020 296.660 ;
        RECT 41.180 295.700 46.740 296.660 ;
        RECT 47.900 295.700 53.460 296.660 ;
        RECT 54.620 295.700 60.180 296.660 ;
        RECT 61.340 295.700 66.900 296.660 ;
        RECT 68.060 295.700 73.620 296.660 ;
        RECT 74.780 295.700 80.340 296.660 ;
        RECT 81.500 295.700 87.060 296.660 ;
        RECT 88.220 295.700 93.780 296.660 ;
        RECT 94.940 295.700 100.500 296.660 ;
        RECT 101.660 295.700 107.220 296.660 ;
        RECT 108.380 295.700 113.940 296.660 ;
        RECT 115.100 295.700 120.660 296.660 ;
        RECT 121.820 295.700 127.380 296.660 ;
        RECT 128.540 295.700 134.100 296.660 ;
        RECT 135.260 295.700 140.820 296.660 ;
        RECT 141.980 295.700 147.540 296.660 ;
        RECT 148.700 295.700 154.260 296.660 ;
        RECT 155.420 295.700 160.980 296.660 ;
        RECT 162.140 295.700 167.700 296.660 ;
        RECT 168.860 295.700 174.420 296.660 ;
        RECT 175.580 295.700 181.140 296.660 ;
        RECT 182.300 295.700 187.860 296.660 ;
        RECT 189.020 295.700 194.580 296.660 ;
        RECT 195.740 295.700 201.300 296.660 ;
        RECT 202.460 295.700 208.020 296.660 ;
        RECT 209.180 295.700 214.740 296.660 ;
        RECT 215.900 295.700 221.460 296.660 ;
        RECT 222.620 295.700 228.180 296.660 ;
        RECT 229.340 295.700 234.900 296.660 ;
        RECT 236.060 295.700 241.620 296.660 ;
        RECT 242.780 295.700 248.340 296.660 ;
        RECT 249.500 295.700 255.060 296.660 ;
        RECT 256.220 295.700 261.780 296.660 ;
        RECT 262.940 295.700 268.500 296.660 ;
        RECT 269.660 295.700 275.220 296.660 ;
        RECT 276.380 295.700 281.940 296.660 ;
        RECT 283.100 295.700 288.660 296.660 ;
        RECT 289.820 295.700 295.380 296.660 ;
        RECT 296.540 295.700 302.100 296.660 ;
        RECT 303.260 295.700 308.820 296.660 ;
        RECT 309.980 295.700 315.540 296.660 ;
        RECT 316.700 295.700 322.260 296.660 ;
        RECT 323.420 295.700 328.980 296.660 ;
        RECT 330.140 295.700 335.700 296.660 ;
        RECT 336.860 295.700 342.420 296.660 ;
        RECT 343.580 295.700 349.140 296.660 ;
        RECT 350.300 295.700 355.860 296.660 ;
        RECT 357.020 295.700 362.580 296.660 ;
        RECT 363.740 295.700 369.300 296.660 ;
        RECT 370.460 295.700 376.020 296.660 ;
        RECT 377.180 295.700 382.740 296.660 ;
        RECT 383.900 295.700 389.460 296.660 ;
        RECT 390.620 295.700 396.180 296.660 ;
        RECT 397.340 295.700 402.900 296.660 ;
        RECT 404.060 295.700 409.620 296.660 ;
        RECT 410.780 295.700 416.340 296.660 ;
        RECT 417.500 295.700 423.060 296.660 ;
        RECT 424.220 295.700 429.780 296.660 ;
        RECT 430.940 295.700 436.500 296.660 ;
        RECT 437.660 295.700 443.220 296.660 ;
        RECT 444.380 295.700 449.940 296.660 ;
        RECT 451.100 295.700 456.660 296.660 ;
        RECT 457.820 295.700 463.380 296.660 ;
        RECT 464.540 295.700 470.100 296.660 ;
        RECT 471.260 295.700 476.820 296.660 ;
        RECT 477.980 295.700 483.540 296.660 ;
        RECT 484.700 295.700 490.260 296.660 ;
        RECT 491.420 295.700 564.180 296.660 ;
        RECT 565.340 295.700 570.900 296.660 ;
        RECT 572.060 295.700 577.620 296.660 ;
        RECT 578.780 295.700 584.340 296.660 ;
        RECT 585.500 295.700 591.060 296.660 ;
        RECT 592.220 295.700 597.780 296.660 ;
        RECT 598.940 295.700 604.500 296.660 ;
        RECT 605.660 295.700 611.220 296.660 ;
        RECT 612.380 295.700 617.940 296.660 ;
        RECT 619.100 295.700 624.660 296.660 ;
        RECT 625.820 295.700 631.380 296.660 ;
        RECT 632.540 295.700 638.100 296.660 ;
        RECT 639.260 295.700 712.020 296.660 ;
        RECT 713.180 295.700 718.740 296.660 ;
        RECT 719.900 295.700 725.460 296.660 ;
        RECT 726.620 295.700 732.180 296.660 ;
        RECT 733.340 295.700 738.900 296.660 ;
        RECT 740.060 295.700 745.620 296.660 ;
        RECT 746.780 295.700 752.340 296.660 ;
        RECT 753.500 295.700 759.060 296.660 ;
        RECT 760.220 295.700 765.780 296.660 ;
        RECT 766.940 295.700 772.500 296.660 ;
        RECT 773.660 295.700 779.220 296.660 ;
        RECT 780.380 295.700 785.940 296.660 ;
        RECT 787.100 295.700 792.660 296.660 ;
        RECT 793.820 295.700 799.380 296.660 ;
        RECT 800.540 295.700 806.100 296.660 ;
        RECT 807.260 295.700 812.820 296.660 ;
        RECT 813.980 295.700 819.540 296.660 ;
        RECT 820.700 295.700 826.260 296.660 ;
        RECT 827.420 295.700 832.980 296.660 ;
        RECT 834.140 295.700 839.700 296.660 ;
        RECT 840.860 295.700 846.420 296.660 ;
        RECT 847.580 295.700 853.140 296.660 ;
        RECT 854.300 295.700 859.860 296.660 ;
        RECT 861.020 295.700 866.580 296.660 ;
        RECT 867.740 295.700 873.300 296.660 ;
        RECT 874.460 295.700 880.020 296.660 ;
        RECT 881.180 295.700 886.740 296.660 ;
        RECT 887.900 295.700 893.460 296.660 ;
        RECT 894.620 295.700 900.180 296.660 ;
        RECT 901.340 295.700 906.900 296.660 ;
        RECT 908.060 295.700 913.620 296.660 ;
        RECT 914.780 295.700 920.340 296.660 ;
        RECT 921.500 295.700 927.060 296.660 ;
        RECT 928.220 295.700 933.780 296.660 ;
        RECT 934.940 295.700 940.500 296.660 ;
        RECT 941.660 295.700 947.220 296.660 ;
        RECT 948.380 295.700 953.940 296.660 ;
        RECT 955.100 295.700 960.660 296.660 ;
        RECT 961.820 295.700 967.380 296.660 ;
        RECT 968.540 295.700 974.100 296.660 ;
        RECT 975.260 295.700 980.820 296.660 ;
        RECT 981.980 295.700 987.540 296.660 ;
        RECT 988.700 295.700 994.260 296.660 ;
        RECT 995.420 295.700 1000.980 296.660 ;
        RECT 1002.140 295.700 1007.700 296.660 ;
        RECT 1008.860 295.700 1014.420 296.660 ;
        RECT 1015.580 295.700 1021.140 296.660 ;
        RECT 1022.300 295.700 1027.860 296.660 ;
        RECT 1029.020 295.700 1034.580 296.660 ;
        RECT 1035.740 295.700 1041.300 296.660 ;
        RECT 1042.460 295.700 1048.020 296.660 ;
        RECT 1049.180 295.700 1054.740 296.660 ;
        RECT 1055.900 295.700 1061.460 296.660 ;
        RECT 1062.620 295.700 1068.180 296.660 ;
        RECT 1069.340 295.700 1074.900 296.660 ;
        RECT 1076.060 295.700 1081.620 296.660 ;
        RECT 1082.780 295.700 1088.340 296.660 ;
        RECT 1089.500 295.700 1095.060 296.660 ;
        RECT 1096.220 295.700 1101.780 296.660 ;
        RECT 1102.940 295.700 1108.500 296.660 ;
        RECT 1109.660 295.700 1115.220 296.660 ;
        RECT 1116.380 295.700 1121.940 296.660 ;
        RECT 1123.100 295.700 1128.660 296.660 ;
        RECT 1129.820 295.700 1135.380 296.660 ;
        RECT 1136.540 295.700 1142.100 296.660 ;
        RECT 1143.260 295.700 1148.820 296.660 ;
        RECT 1149.980 295.700 1155.540 296.660 ;
        RECT 1156.700 295.700 1162.260 296.660 ;
        RECT 1163.420 295.700 1168.980 296.660 ;
        RECT 1170.140 295.700 1444.500 296.660 ;
        RECT 1445.660 295.700 1451.220 296.660 ;
        RECT 1452.380 295.700 1457.940 296.660 ;
        RECT 1459.100 295.700 1464.660 296.660 ;
        RECT 1465.820 295.700 1471.380 296.660 ;
        RECT 1472.540 295.700 1478.100 296.660 ;
        RECT 1479.260 295.700 1484.820 296.660 ;
        RECT 1485.980 295.700 1491.540 296.660 ;
        RECT 1492.700 295.700 1498.260 296.660 ;
        RECT 1499.420 295.700 1504.980 296.660 ;
        RECT 1506.140 295.700 1511.700 296.660 ;
        RECT 1512.860 295.700 1518.420 296.660 ;
        RECT 1519.580 295.700 1525.140 296.660 ;
        RECT 1526.300 295.700 1531.860 296.660 ;
        RECT 1533.020 295.700 1538.580 296.660 ;
        RECT 1539.740 295.700 1545.300 296.660 ;
        RECT 1546.460 295.700 1552.020 296.660 ;
        RECT 1553.180 295.700 1558.740 296.660 ;
        RECT 1559.900 295.700 1565.460 296.660 ;
        RECT 1566.620 295.700 1572.180 296.660 ;
        RECT 1573.340 295.700 1578.900 296.660 ;
        RECT 1580.060 295.700 1585.620 296.660 ;
        RECT 1586.780 295.700 1592.340 296.660 ;
        RECT 1593.500 295.700 1599.060 296.660 ;
        RECT 1600.220 295.700 1605.780 296.660 ;
        RECT 1606.940 295.700 1612.500 296.660 ;
        RECT 1613.660 295.700 1619.220 296.660 ;
        RECT 1620.380 295.700 1625.940 296.660 ;
        RECT 1627.100 295.700 1632.660 296.660 ;
        RECT 1633.820 295.700 1639.380 296.660 ;
        RECT 1640.540 295.700 1646.100 296.660 ;
        RECT 1647.260 295.700 1652.820 296.660 ;
        RECT 1653.980 295.700 1659.540 296.660 ;
        RECT 1660.700 295.700 1666.260 296.660 ;
        RECT 1667.420 295.700 1672.980 296.660 ;
        RECT 1674.140 295.700 1679.700 296.660 ;
        RECT 1680.860 295.700 1686.420 296.660 ;
        RECT 1687.580 295.700 1693.140 296.660 ;
        RECT 1694.300 295.700 1699.860 296.660 ;
        RECT 1701.020 295.700 1706.580 296.660 ;
        RECT 1707.740 295.700 1713.300 296.660 ;
        RECT 1714.460 295.700 1720.020 296.660 ;
        RECT 1721.180 295.700 1726.740 296.660 ;
        RECT 1727.900 295.700 1733.460 296.660 ;
        RECT 1734.620 295.700 1740.180 296.660 ;
        RECT 1741.340 295.700 1746.900 296.660 ;
        RECT 1748.060 295.700 1753.620 296.660 ;
        RECT 1754.780 295.700 1760.340 296.660 ;
        RECT 1761.500 295.700 1767.060 296.660 ;
        RECT 1768.220 295.700 1773.780 296.660 ;
        RECT 1774.940 295.700 1780.500 296.660 ;
        RECT 1781.660 295.700 1787.220 296.660 ;
        RECT 1788.380 295.700 1793.940 296.660 ;
        RECT 1795.100 295.700 1800.660 296.660 ;
        RECT 1801.820 295.700 1807.380 296.660 ;
        RECT 1808.540 295.700 1814.100 296.660 ;
        RECT 1815.260 295.700 1820.820 296.660 ;
        RECT 1821.980 295.700 1827.540 296.660 ;
        RECT 1828.700 295.700 1834.260 296.660 ;
        RECT 1835.420 295.700 1840.980 296.660 ;
        RECT 1842.140 295.700 1847.700 296.660 ;
        RECT 1848.860 295.700 1854.420 296.660 ;
        RECT 1855.580 295.700 1861.140 296.660 ;
        RECT 1862.300 295.700 1867.860 296.660 ;
        RECT 1869.020 295.700 1908.180 296.660 ;
        RECT 1909.340 295.700 1914.900 296.660 ;
        RECT 1916.060 295.700 1921.620 296.660 ;
        RECT 1922.780 295.700 1928.340 296.660 ;
        RECT 1929.500 295.700 1935.060 296.660 ;
        RECT 1936.220 295.700 1941.780 296.660 ;
        RECT 1942.940 295.700 1948.500 296.660 ;
        RECT 1949.660 295.700 1955.220 296.660 ;
        RECT 1956.380 295.700 1961.940 296.660 ;
        RECT 1963.100 295.700 2002.260 296.660 ;
        RECT 2003.420 295.700 2008.980 296.660 ;
        RECT 2010.140 295.700 2015.700 296.660 ;
        RECT 2016.860 295.700 2022.420 296.660 ;
        RECT 2023.580 295.700 2029.140 296.660 ;
        RECT 2030.300 295.700 2035.860 296.660 ;
        RECT 2037.020 295.700 2042.580 296.660 ;
        RECT 2043.740 295.700 2049.300 296.660 ;
        RECT 2050.460 295.700 2056.020 296.660 ;
        RECT 2057.180 295.700 2062.740 296.660 ;
        RECT 2063.900 295.700 2069.460 296.660 ;
        RECT 2070.620 295.700 2076.180 296.660 ;
        RECT 2077.340 295.700 2082.900 296.660 ;
        RECT 2084.060 295.700 2089.620 296.660 ;
        RECT 2090.780 295.700 2096.340 296.660 ;
        RECT 2097.500 295.700 2103.060 296.660 ;
        RECT 2104.220 295.700 2109.780 296.660 ;
        RECT 2110.940 295.700 2116.500 296.660 ;
        RECT 2117.660 295.700 2123.220 296.660 ;
        RECT 2124.380 295.700 2129.940 296.660 ;
        RECT 2131.100 295.700 2136.660 296.660 ;
        RECT 2137.820 295.700 2143.380 296.660 ;
        RECT 2144.540 295.700 2150.100 296.660 ;
        RECT 2151.260 295.700 2156.820 296.660 ;
        RECT 2157.980 295.700 2163.540 296.660 ;
        RECT 2164.700 295.700 2170.260 296.660 ;
        RECT 2171.420 295.700 2176.980 296.660 ;
        RECT 2178.140 295.700 2183.700 296.660 ;
        RECT 2184.860 295.700 2190.420 296.660 ;
        RECT 2191.580 295.700 2197.140 296.660 ;
        RECT 2198.300 295.700 2203.860 296.660 ;
        RECT 2205.020 295.700 2210.580 296.660 ;
        RECT 2211.740 295.700 2217.300 296.660 ;
        RECT 2218.460 295.700 2224.020 296.660 ;
        RECT 2225.180 295.700 2230.740 296.660 ;
        RECT 2231.900 295.700 2237.460 296.660 ;
        RECT 2238.620 295.700 2244.180 296.660 ;
        RECT 2245.340 295.700 2250.900 296.660 ;
        RECT 2252.060 295.700 2257.620 296.660 ;
        RECT 2258.780 295.700 2264.340 296.660 ;
        RECT 2265.500 295.700 2271.060 296.660 ;
        RECT 2272.220 295.700 2277.780 296.660 ;
        RECT 2278.940 295.700 2284.500 296.660 ;
        RECT 2285.660 295.700 2291.220 296.660 ;
        RECT 2292.380 295.700 2297.940 296.660 ;
        RECT 2299.100 295.700 2304.660 296.660 ;
        RECT 2305.820 295.700 2311.380 296.660 ;
        RECT 2312.540 295.700 2318.100 296.660 ;
        RECT 2319.260 295.700 2324.820 296.660 ;
        RECT 2325.980 295.700 2331.540 296.660 ;
        RECT 2332.700 295.700 2338.260 296.660 ;
        RECT 2339.420 295.700 2344.980 296.660 ;
        RECT 2346.140 295.700 2351.700 296.660 ;
        RECT 2352.860 295.700 2358.420 296.660 ;
        RECT 2359.580 295.700 2365.140 296.660 ;
        RECT 2366.300 295.700 2391.620 296.660 ;
        RECT 8.540 4.300 2391.620 295.700 ;
        RECT 8.540 2.330 43.380 4.300 ;
        RECT 44.540 2.330 50.100 4.300 ;
        RECT 51.260 2.330 56.820 4.300 ;
        RECT 57.980 2.330 63.540 4.300 ;
        RECT 64.700 2.330 70.260 4.300 ;
        RECT 71.420 2.330 76.980 4.300 ;
        RECT 78.140 2.330 83.700 4.300 ;
        RECT 84.860 2.330 90.420 4.300 ;
        RECT 91.580 2.330 97.140 4.300 ;
        RECT 98.300 2.330 103.860 4.300 ;
        RECT 105.020 2.330 110.580 4.300 ;
        RECT 111.740 2.330 117.300 4.300 ;
        RECT 118.460 2.330 124.020 4.300 ;
        RECT 125.180 2.330 130.740 4.300 ;
        RECT 131.900 2.330 137.460 4.300 ;
        RECT 138.620 2.330 144.180 4.300 ;
        RECT 145.340 2.330 150.900 4.300 ;
        RECT 152.060 2.330 157.620 4.300 ;
        RECT 158.780 2.330 164.340 4.300 ;
        RECT 165.500 2.330 171.060 4.300 ;
        RECT 172.220 2.330 177.780 4.300 ;
        RECT 178.940 2.330 184.500 4.300 ;
        RECT 185.660 2.330 191.220 4.300 ;
        RECT 192.380 2.330 197.940 4.300 ;
        RECT 199.100 2.330 204.660 4.300 ;
        RECT 205.820 2.330 211.380 4.300 ;
        RECT 212.540 2.330 218.100 4.300 ;
        RECT 219.260 2.330 224.820 4.300 ;
        RECT 225.980 2.330 231.540 4.300 ;
        RECT 232.700 2.330 238.260 4.300 ;
        RECT 239.420 2.330 244.980 4.300 ;
        RECT 246.140 2.330 251.700 4.300 ;
        RECT 252.860 2.330 258.420 4.300 ;
        RECT 259.580 2.330 265.140 4.300 ;
        RECT 266.300 2.330 271.860 4.300 ;
        RECT 273.020 2.330 278.580 4.300 ;
        RECT 279.740 2.330 285.300 4.300 ;
        RECT 286.460 2.330 292.020 4.300 ;
        RECT 293.180 2.330 298.740 4.300 ;
        RECT 299.900 2.330 305.460 4.300 ;
        RECT 306.620 2.330 312.180 4.300 ;
        RECT 313.340 2.330 318.900 4.300 ;
        RECT 320.060 2.330 325.620 4.300 ;
        RECT 326.780 2.330 332.340 4.300 ;
        RECT 333.500 2.330 339.060 4.300 ;
        RECT 340.220 2.330 345.780 4.300 ;
        RECT 346.940 2.330 352.500 4.300 ;
        RECT 353.660 2.330 359.220 4.300 ;
        RECT 360.380 2.330 365.940 4.300 ;
        RECT 367.100 2.330 372.660 4.300 ;
        RECT 373.820 2.330 379.380 4.300 ;
        RECT 380.540 2.330 386.100 4.300 ;
        RECT 387.260 2.330 392.820 4.300 ;
        RECT 393.980 2.330 399.540 4.300 ;
        RECT 400.700 2.330 406.260 4.300 ;
        RECT 407.420 2.330 412.980 4.300 ;
        RECT 414.140 2.330 419.700 4.300 ;
        RECT 420.860 2.330 426.420 4.300 ;
        RECT 427.580 2.330 433.140 4.300 ;
        RECT 434.300 2.330 439.860 4.300 ;
        RECT 441.020 2.330 446.580 4.300 ;
        RECT 447.740 2.330 453.300 4.300 ;
        RECT 454.460 2.330 460.020 4.300 ;
        RECT 461.180 2.330 466.740 4.300 ;
        RECT 467.900 2.330 473.460 4.300 ;
        RECT 474.620 2.330 480.180 4.300 ;
        RECT 481.340 2.330 486.900 4.300 ;
        RECT 488.060 2.330 527.220 4.300 ;
        RECT 528.380 2.330 533.940 4.300 ;
        RECT 535.100 2.330 540.660 4.300 ;
        RECT 541.820 2.330 547.380 4.300 ;
        RECT 548.540 2.330 554.100 4.300 ;
        RECT 555.260 2.330 560.820 4.300 ;
        RECT 561.980 2.330 567.540 4.300 ;
        RECT 568.700 2.330 574.260 4.300 ;
        RECT 575.420 2.330 580.980 4.300 ;
        RECT 582.140 2.330 587.700 4.300 ;
        RECT 588.860 2.330 594.420 4.300 ;
        RECT 595.580 2.330 601.140 4.300 ;
        RECT 602.300 2.330 607.860 4.300 ;
        RECT 609.020 2.330 614.580 4.300 ;
        RECT 615.740 2.330 621.300 4.300 ;
        RECT 622.460 2.330 628.020 4.300 ;
        RECT 629.180 2.330 634.740 4.300 ;
        RECT 635.900 2.330 641.460 4.300 ;
        RECT 642.620 2.330 648.180 4.300 ;
        RECT 649.340 2.330 654.900 4.300 ;
        RECT 656.060 2.330 661.620 4.300 ;
        RECT 662.780 2.330 668.340 4.300 ;
        RECT 669.500 2.330 675.060 4.300 ;
        RECT 676.220 2.330 681.780 4.300 ;
        RECT 682.940 2.330 688.500 4.300 ;
        RECT 689.660 2.330 695.220 4.300 ;
        RECT 696.380 2.330 701.940 4.300 ;
        RECT 703.100 2.330 708.660 4.300 ;
        RECT 709.820 2.330 715.380 4.300 ;
        RECT 716.540 2.330 722.100 4.300 ;
        RECT 723.260 2.330 728.820 4.300 ;
        RECT 729.980 2.330 735.540 4.300 ;
        RECT 736.700 2.330 742.260 4.300 ;
        RECT 743.420 2.330 748.980 4.300 ;
        RECT 750.140 2.330 755.700 4.300 ;
        RECT 756.860 2.330 762.420 4.300 ;
        RECT 763.580 2.330 769.140 4.300 ;
        RECT 770.300 2.330 775.860 4.300 ;
        RECT 777.020 2.330 782.580 4.300 ;
        RECT 783.740 2.330 789.300 4.300 ;
        RECT 790.460 2.330 796.020 4.300 ;
        RECT 797.180 2.330 802.740 4.300 ;
        RECT 803.900 2.330 809.460 4.300 ;
        RECT 810.620 2.330 816.180 4.300 ;
        RECT 817.340 2.330 822.900 4.300 ;
        RECT 824.060 2.330 829.620 4.300 ;
        RECT 830.780 2.330 836.340 4.300 ;
        RECT 837.500 2.330 843.060 4.300 ;
        RECT 844.220 2.330 849.780 4.300 ;
        RECT 850.940 2.330 856.500 4.300 ;
        RECT 857.660 2.330 863.220 4.300 ;
        RECT 864.380 2.330 869.940 4.300 ;
        RECT 871.100 2.330 876.660 4.300 ;
        RECT 877.820 2.330 883.380 4.300 ;
        RECT 884.540 2.330 890.100 4.300 ;
        RECT 891.260 2.330 896.820 4.300 ;
        RECT 897.980 2.330 903.540 4.300 ;
        RECT 904.700 2.330 910.260 4.300 ;
        RECT 911.420 2.330 916.980 4.300 ;
        RECT 918.140 2.330 923.700 4.300 ;
        RECT 924.860 2.330 930.420 4.300 ;
        RECT 931.580 2.330 937.140 4.300 ;
        RECT 938.300 2.330 943.860 4.300 ;
        RECT 945.020 2.330 950.580 4.300 ;
        RECT 951.740 2.330 957.300 4.300 ;
        RECT 958.460 2.330 964.020 4.300 ;
        RECT 965.180 2.330 970.740 4.300 ;
        RECT 971.900 2.330 977.460 4.300 ;
        RECT 978.620 2.330 984.180 4.300 ;
        RECT 985.340 2.330 990.900 4.300 ;
        RECT 992.060 2.330 997.620 4.300 ;
        RECT 998.780 2.330 1004.340 4.300 ;
        RECT 1005.500 2.330 1011.060 4.300 ;
        RECT 1012.220 2.330 1017.780 4.300 ;
        RECT 1018.940 2.330 1024.500 4.300 ;
        RECT 1025.660 2.330 1031.220 4.300 ;
        RECT 1032.380 2.330 1037.940 4.300 ;
        RECT 1039.100 2.330 1044.660 4.300 ;
        RECT 1045.820 2.330 1051.380 4.300 ;
        RECT 1052.540 2.330 1125.300 4.300 ;
        RECT 1126.460 2.330 1132.020 4.300 ;
        RECT 1133.180 2.330 1138.740 4.300 ;
        RECT 1139.900 2.330 1145.460 4.300 ;
        RECT 1146.620 2.330 1152.180 4.300 ;
        RECT 1153.340 2.330 1158.900 4.300 ;
        RECT 1160.060 2.330 1165.620 4.300 ;
        RECT 1166.780 2.330 1172.340 4.300 ;
        RECT 1173.500 2.330 1179.060 4.300 ;
        RECT 1180.220 2.330 1185.780 4.300 ;
        RECT 1186.940 2.330 1192.500 4.300 ;
        RECT 1193.660 2.330 1199.220 4.300 ;
        RECT 1200.380 2.330 1205.940 4.300 ;
        RECT 1207.100 2.330 1212.660 4.300 ;
        RECT 1213.820 2.330 1219.380 4.300 ;
        RECT 1220.540 2.330 1226.100 4.300 ;
        RECT 1227.260 2.330 1434.420 4.300 ;
        RECT 1435.580 2.330 1441.140 4.300 ;
        RECT 1442.300 2.330 1447.860 4.300 ;
        RECT 1449.020 2.330 1454.580 4.300 ;
        RECT 1455.740 2.330 1461.300 4.300 ;
        RECT 1462.460 2.330 1468.020 4.300 ;
        RECT 1469.180 2.330 1474.740 4.300 ;
        RECT 1475.900 2.330 1481.460 4.300 ;
        RECT 1482.620 2.330 1488.180 4.300 ;
        RECT 1489.340 2.330 1494.900 4.300 ;
        RECT 1496.060 2.330 1501.620 4.300 ;
        RECT 1502.780 2.330 1508.340 4.300 ;
        RECT 1509.500 2.330 1515.060 4.300 ;
        RECT 1516.220 2.330 1521.780 4.300 ;
        RECT 1522.940 2.330 1528.500 4.300 ;
        RECT 1529.660 2.330 1535.220 4.300 ;
        RECT 1536.380 2.330 1541.940 4.300 ;
        RECT 1543.100 2.330 1548.660 4.300 ;
        RECT 1549.820 2.330 1555.380 4.300 ;
        RECT 1556.540 2.330 1562.100 4.300 ;
        RECT 1563.260 2.330 1568.820 4.300 ;
        RECT 1569.980 2.330 1575.540 4.300 ;
        RECT 1576.700 2.330 1582.260 4.300 ;
        RECT 1583.420 2.330 1588.980 4.300 ;
        RECT 1590.140 2.330 1595.700 4.300 ;
        RECT 1596.860 2.330 1602.420 4.300 ;
        RECT 1603.580 2.330 1609.140 4.300 ;
        RECT 1610.300 2.330 1615.860 4.300 ;
        RECT 1617.020 2.330 1622.580 4.300 ;
        RECT 1623.740 2.330 1629.300 4.300 ;
        RECT 1630.460 2.330 1636.020 4.300 ;
        RECT 1637.180 2.330 1642.740 4.300 ;
        RECT 1643.900 2.330 1649.460 4.300 ;
        RECT 1650.620 2.330 1656.180 4.300 ;
        RECT 1657.340 2.330 1662.900 4.300 ;
        RECT 1664.060 2.330 1669.620 4.300 ;
        RECT 1670.780 2.330 1676.340 4.300 ;
        RECT 1677.500 2.330 1683.060 4.300 ;
        RECT 1684.220 2.330 1689.780 4.300 ;
        RECT 1690.940 2.330 1696.500 4.300 ;
        RECT 1697.660 2.330 1703.220 4.300 ;
        RECT 1704.380 2.330 1709.940 4.300 ;
        RECT 1711.100 2.330 1716.660 4.300 ;
        RECT 1717.820 2.330 1723.380 4.300 ;
        RECT 1724.540 2.330 1730.100 4.300 ;
        RECT 1731.260 2.330 1736.820 4.300 ;
        RECT 1737.980 2.330 1743.540 4.300 ;
        RECT 1744.700 2.330 1750.260 4.300 ;
        RECT 1751.420 2.330 1756.980 4.300 ;
        RECT 1758.140 2.330 1763.700 4.300 ;
        RECT 1764.860 2.330 1770.420 4.300 ;
        RECT 1771.580 2.330 1777.140 4.300 ;
        RECT 1778.300 2.330 1783.860 4.300 ;
        RECT 1785.020 2.330 1790.580 4.300 ;
        RECT 1791.740 2.330 1797.300 4.300 ;
        RECT 1798.460 2.330 1804.020 4.300 ;
        RECT 1805.180 2.330 1810.740 4.300 ;
        RECT 1811.900 2.330 1817.460 4.300 ;
        RECT 1818.620 2.330 1824.180 4.300 ;
        RECT 1825.340 2.330 1830.900 4.300 ;
        RECT 1832.060 2.330 1837.620 4.300 ;
        RECT 1838.780 2.330 1844.340 4.300 ;
        RECT 1845.500 2.330 1851.060 4.300 ;
        RECT 1852.220 2.330 1857.780 4.300 ;
        RECT 1858.940 2.330 1864.500 4.300 ;
        RECT 1865.660 2.330 1871.220 4.300 ;
        RECT 1872.380 2.330 1877.940 4.300 ;
        RECT 1879.100 2.330 1884.660 4.300 ;
        RECT 1885.820 2.330 1891.380 4.300 ;
        RECT 1892.540 2.330 1898.100 4.300 ;
        RECT 1899.260 2.330 1904.820 4.300 ;
        RECT 1905.980 2.330 1911.540 4.300 ;
        RECT 1912.700 2.330 1918.260 4.300 ;
        RECT 1919.420 2.330 1924.980 4.300 ;
        RECT 1926.140 2.330 1931.700 4.300 ;
        RECT 1932.860 2.330 1938.420 4.300 ;
        RECT 1939.580 2.330 1945.140 4.300 ;
        RECT 1946.300 2.330 1951.860 4.300 ;
        RECT 1953.020 2.330 1958.580 4.300 ;
        RECT 1959.740 2.330 1965.300 4.300 ;
        RECT 1966.460 2.330 1972.020 4.300 ;
        RECT 1973.180 2.330 1978.740 4.300 ;
        RECT 1979.900 2.330 1985.460 4.300 ;
        RECT 1986.620 2.330 1992.180 4.300 ;
        RECT 1993.340 2.330 1998.900 4.300 ;
        RECT 2000.060 2.330 2005.620 4.300 ;
        RECT 2006.780 2.330 2012.340 4.300 ;
        RECT 2013.500 2.330 2019.060 4.300 ;
        RECT 2020.220 2.330 2025.780 4.300 ;
        RECT 2026.940 2.330 2032.500 4.300 ;
        RECT 2033.660 2.330 2039.220 4.300 ;
        RECT 2040.380 2.330 2045.940 4.300 ;
        RECT 2047.100 2.330 2052.660 4.300 ;
        RECT 2053.820 2.330 2059.380 4.300 ;
        RECT 2060.540 2.330 2066.100 4.300 ;
        RECT 2067.260 2.330 2072.820 4.300 ;
        RECT 2073.980 2.330 2079.540 4.300 ;
        RECT 2080.700 2.330 2086.260 4.300 ;
        RECT 2087.420 2.330 2092.980 4.300 ;
        RECT 2094.140 2.330 2099.700 4.300 ;
        RECT 2100.860 2.330 2106.420 4.300 ;
        RECT 2107.580 2.330 2113.140 4.300 ;
        RECT 2114.300 2.330 2119.860 4.300 ;
        RECT 2121.020 2.330 2126.580 4.300 ;
        RECT 2127.740 2.330 2133.300 4.300 ;
        RECT 2134.460 2.330 2391.620 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 289.780 2395.700 290.500 ;
        RECT 4.000 286.460 2396.660 289.780 ;
        RECT 4.000 285.300 2395.700 286.460 ;
        RECT 4.000 281.980 2396.660 285.300 ;
        RECT 4.000 280.820 2395.700 281.980 ;
        RECT 4.000 278.620 2396.660 280.820 ;
        RECT 4.300 277.500 2396.660 278.620 ;
        RECT 4.300 277.460 2395.700 277.500 ;
        RECT 4.000 276.340 2395.700 277.460 ;
        RECT 4.000 273.020 2396.660 276.340 ;
        RECT 4.300 271.860 2395.700 273.020 ;
        RECT 4.000 268.540 2396.660 271.860 ;
        RECT 4.000 267.420 2395.700 268.540 ;
        RECT 4.300 267.380 2395.700 267.420 ;
        RECT 4.300 266.260 2396.660 267.380 ;
        RECT 4.000 264.060 2396.660 266.260 ;
        RECT 4.000 262.900 2395.700 264.060 ;
        RECT 4.000 261.820 2396.660 262.900 ;
        RECT 4.300 260.660 2396.660 261.820 ;
        RECT 4.000 259.580 2396.660 260.660 ;
        RECT 4.000 258.420 2395.700 259.580 ;
        RECT 4.000 256.220 2396.660 258.420 ;
        RECT 4.300 255.100 2396.660 256.220 ;
        RECT 4.300 255.060 2395.700 255.100 ;
        RECT 4.000 253.940 2395.700 255.060 ;
        RECT 4.000 250.620 2396.660 253.940 ;
        RECT 4.300 249.460 2395.700 250.620 ;
        RECT 4.000 246.140 2396.660 249.460 ;
        RECT 4.000 245.020 2395.700 246.140 ;
        RECT 4.300 244.980 2395.700 245.020 ;
        RECT 4.300 243.860 2396.660 244.980 ;
        RECT 4.000 241.660 2396.660 243.860 ;
        RECT 4.000 240.500 2395.700 241.660 ;
        RECT 4.000 239.420 2396.660 240.500 ;
        RECT 4.300 238.260 2396.660 239.420 ;
        RECT 4.000 237.180 2396.660 238.260 ;
        RECT 4.000 236.020 2395.700 237.180 ;
        RECT 4.000 233.820 2396.660 236.020 ;
        RECT 4.300 232.700 2396.660 233.820 ;
        RECT 4.300 232.660 2395.700 232.700 ;
        RECT 4.000 231.540 2395.700 232.660 ;
        RECT 4.000 228.220 2396.660 231.540 ;
        RECT 4.300 227.060 2395.700 228.220 ;
        RECT 4.000 223.740 2396.660 227.060 ;
        RECT 4.000 222.620 2395.700 223.740 ;
        RECT 4.300 222.580 2395.700 222.620 ;
        RECT 4.300 221.460 2396.660 222.580 ;
        RECT 4.000 219.260 2396.660 221.460 ;
        RECT 4.000 218.100 2395.700 219.260 ;
        RECT 4.000 217.020 2396.660 218.100 ;
        RECT 4.300 215.860 2396.660 217.020 ;
        RECT 4.000 214.780 2396.660 215.860 ;
        RECT 4.000 213.620 2395.700 214.780 ;
        RECT 4.000 211.420 2396.660 213.620 ;
        RECT 4.300 210.300 2396.660 211.420 ;
        RECT 4.300 210.260 2395.700 210.300 ;
        RECT 4.000 209.140 2395.700 210.260 ;
        RECT 4.000 205.820 2396.660 209.140 ;
        RECT 4.300 204.660 2395.700 205.820 ;
        RECT 4.000 201.340 2396.660 204.660 ;
        RECT 4.000 200.220 2395.700 201.340 ;
        RECT 4.300 200.180 2395.700 200.220 ;
        RECT 4.300 199.060 2396.660 200.180 ;
        RECT 4.000 196.860 2396.660 199.060 ;
        RECT 4.000 195.700 2395.700 196.860 ;
        RECT 4.000 194.620 2396.660 195.700 ;
        RECT 4.300 193.460 2396.660 194.620 ;
        RECT 4.000 192.380 2396.660 193.460 ;
        RECT 4.000 191.220 2395.700 192.380 ;
        RECT 4.000 189.020 2396.660 191.220 ;
        RECT 4.300 187.900 2396.660 189.020 ;
        RECT 4.300 187.860 2395.700 187.900 ;
        RECT 4.000 186.740 2395.700 187.860 ;
        RECT 4.000 183.420 2396.660 186.740 ;
        RECT 4.300 182.260 2395.700 183.420 ;
        RECT 4.000 178.940 2396.660 182.260 ;
        RECT 4.000 177.820 2395.700 178.940 ;
        RECT 4.300 177.780 2395.700 177.820 ;
        RECT 4.300 176.660 2396.660 177.780 ;
        RECT 4.000 174.460 2396.660 176.660 ;
        RECT 4.000 173.300 2395.700 174.460 ;
        RECT 4.000 172.220 2396.660 173.300 ;
        RECT 4.300 171.060 2396.660 172.220 ;
        RECT 4.000 169.980 2396.660 171.060 ;
        RECT 4.000 168.820 2395.700 169.980 ;
        RECT 4.000 166.620 2396.660 168.820 ;
        RECT 4.300 165.500 2396.660 166.620 ;
        RECT 4.300 165.460 2395.700 165.500 ;
        RECT 4.000 164.340 2395.700 165.460 ;
        RECT 4.000 161.020 2396.660 164.340 ;
        RECT 4.300 159.860 2395.700 161.020 ;
        RECT 4.000 156.540 2396.660 159.860 ;
        RECT 4.000 155.420 2395.700 156.540 ;
        RECT 4.300 155.380 2395.700 155.420 ;
        RECT 4.300 154.260 2396.660 155.380 ;
        RECT 4.000 152.060 2396.660 154.260 ;
        RECT 4.000 150.900 2395.700 152.060 ;
        RECT 4.000 149.820 2396.660 150.900 ;
        RECT 4.300 148.660 2396.660 149.820 ;
        RECT 4.000 147.580 2396.660 148.660 ;
        RECT 4.000 146.420 2395.700 147.580 ;
        RECT 4.000 144.220 2396.660 146.420 ;
        RECT 4.300 143.100 2396.660 144.220 ;
        RECT 4.300 143.060 2395.700 143.100 ;
        RECT 4.000 141.940 2395.700 143.060 ;
        RECT 4.000 138.620 2396.660 141.940 ;
        RECT 4.300 137.460 2395.700 138.620 ;
        RECT 4.000 134.140 2396.660 137.460 ;
        RECT 4.000 133.020 2395.700 134.140 ;
        RECT 4.300 132.980 2395.700 133.020 ;
        RECT 4.300 131.860 2396.660 132.980 ;
        RECT 4.000 129.660 2396.660 131.860 ;
        RECT 4.000 128.500 2395.700 129.660 ;
        RECT 4.000 127.420 2396.660 128.500 ;
        RECT 4.300 126.260 2396.660 127.420 ;
        RECT 4.000 125.180 2396.660 126.260 ;
        RECT 4.000 124.020 2395.700 125.180 ;
        RECT 4.000 121.820 2396.660 124.020 ;
        RECT 4.300 120.700 2396.660 121.820 ;
        RECT 4.300 120.660 2395.700 120.700 ;
        RECT 4.000 119.540 2395.700 120.660 ;
        RECT 4.000 116.220 2396.660 119.540 ;
        RECT 4.300 115.060 2395.700 116.220 ;
        RECT 4.000 111.740 2396.660 115.060 ;
        RECT 4.000 110.620 2395.700 111.740 ;
        RECT 4.300 110.580 2395.700 110.620 ;
        RECT 4.300 109.460 2396.660 110.580 ;
        RECT 4.000 107.260 2396.660 109.460 ;
        RECT 4.000 106.100 2395.700 107.260 ;
        RECT 4.000 105.020 2396.660 106.100 ;
        RECT 4.300 103.860 2396.660 105.020 ;
        RECT 4.000 102.780 2396.660 103.860 ;
        RECT 4.000 101.620 2395.700 102.780 ;
        RECT 4.000 99.420 2396.660 101.620 ;
        RECT 4.300 98.300 2396.660 99.420 ;
        RECT 4.300 98.260 2395.700 98.300 ;
        RECT 4.000 97.140 2395.700 98.260 ;
        RECT 4.000 93.820 2396.660 97.140 ;
        RECT 4.300 92.660 2395.700 93.820 ;
        RECT 4.000 89.340 2396.660 92.660 ;
        RECT 4.000 88.220 2395.700 89.340 ;
        RECT 4.300 88.180 2395.700 88.220 ;
        RECT 4.300 87.060 2396.660 88.180 ;
        RECT 4.000 84.860 2396.660 87.060 ;
        RECT 4.000 83.700 2395.700 84.860 ;
        RECT 4.000 82.620 2396.660 83.700 ;
        RECT 4.300 81.460 2396.660 82.620 ;
        RECT 4.000 80.380 2396.660 81.460 ;
        RECT 4.000 79.220 2395.700 80.380 ;
        RECT 4.000 77.020 2396.660 79.220 ;
        RECT 4.300 75.900 2396.660 77.020 ;
        RECT 4.300 75.860 2395.700 75.900 ;
        RECT 4.000 74.740 2395.700 75.860 ;
        RECT 4.000 71.420 2396.660 74.740 ;
        RECT 4.300 70.260 2395.700 71.420 ;
        RECT 4.000 66.940 2396.660 70.260 ;
        RECT 4.000 65.820 2395.700 66.940 ;
        RECT 4.300 65.780 2395.700 65.820 ;
        RECT 4.300 64.660 2396.660 65.780 ;
        RECT 4.000 62.460 2396.660 64.660 ;
        RECT 4.000 61.300 2395.700 62.460 ;
        RECT 4.000 60.220 2396.660 61.300 ;
        RECT 4.300 59.060 2396.660 60.220 ;
        RECT 4.000 57.980 2396.660 59.060 ;
        RECT 4.000 56.820 2395.700 57.980 ;
        RECT 4.000 54.620 2396.660 56.820 ;
        RECT 4.300 53.500 2396.660 54.620 ;
        RECT 4.300 53.460 2395.700 53.500 ;
        RECT 4.000 52.340 2395.700 53.460 ;
        RECT 4.000 49.020 2396.660 52.340 ;
        RECT 4.300 47.860 2395.700 49.020 ;
        RECT 4.000 44.540 2396.660 47.860 ;
        RECT 4.000 43.420 2395.700 44.540 ;
        RECT 4.300 43.380 2395.700 43.420 ;
        RECT 4.300 42.260 2396.660 43.380 ;
        RECT 4.000 40.060 2396.660 42.260 ;
        RECT 4.000 38.900 2395.700 40.060 ;
        RECT 4.000 37.820 2396.660 38.900 ;
        RECT 4.300 36.660 2396.660 37.820 ;
        RECT 4.000 35.580 2396.660 36.660 ;
        RECT 4.000 34.420 2395.700 35.580 ;
        RECT 4.000 32.220 2396.660 34.420 ;
        RECT 4.300 31.100 2396.660 32.220 ;
        RECT 4.300 31.060 2395.700 31.100 ;
        RECT 4.000 29.940 2395.700 31.060 ;
        RECT 4.000 26.620 2396.660 29.940 ;
        RECT 4.300 25.460 2395.700 26.620 ;
        RECT 4.000 22.140 2396.660 25.460 ;
        RECT 4.000 21.020 2395.700 22.140 ;
        RECT 4.300 20.980 2395.700 21.020 ;
        RECT 4.300 19.860 2396.660 20.980 ;
        RECT 4.000 17.660 2396.660 19.860 ;
        RECT 4.000 16.500 2395.700 17.660 ;
        RECT 4.000 13.180 2396.660 16.500 ;
        RECT 4.000 12.020 2395.700 13.180 ;
        RECT 4.000 8.700 2396.660 12.020 ;
        RECT 4.000 7.540 2395.700 8.700 ;
        RECT 4.000 2.380 2396.660 7.540 ;
      LAYER Metal4 ;
        RECT 693.980 20.810 713.140 277.110 ;
        RECT 715.340 20.810 789.940 277.110 ;
        RECT 792.140 20.810 866.740 277.110 ;
        RECT 868.940 20.810 943.540 277.110 ;
        RECT 945.740 20.810 1020.340 277.110 ;
        RECT 1022.540 20.810 1097.140 277.110 ;
        RECT 1099.340 20.810 1173.940 277.110 ;
        RECT 1176.140 20.810 1250.740 277.110 ;
        RECT 1252.940 20.810 1327.540 277.110 ;
        RECT 1329.740 20.810 1404.340 277.110 ;
        RECT 1406.540 20.810 1481.140 277.110 ;
        RECT 1483.340 20.810 1557.940 277.110 ;
        RECT 1560.140 20.810 1634.740 277.110 ;
        RECT 1636.940 20.810 1711.540 277.110 ;
        RECT 1713.740 20.810 1720.180 277.110 ;
  END
END top_design_mux
END LIBRARY

