magic
tech gf180mcuD
magscale 1 10
timestamp 1702319510
<< metal1 >>
rect 1344 41578 39984 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 39984 41578
rect 1344 41492 39984 41526
rect 1344 40794 39984 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 39984 40794
rect 1344 40708 39984 40742
rect 1344 40010 39984 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 39984 40010
rect 1344 39924 39984 39958
rect 9986 39678 9998 39730
rect 10050 39678 10062 39730
rect 18610 39678 18622 39730
rect 18674 39678 18686 39730
rect 21298 39678 21310 39730
rect 21362 39678 21374 39730
rect 24670 39618 24722 39630
rect 12898 39566 12910 39618
rect 12962 39566 12974 39618
rect 15698 39566 15710 39618
rect 15762 39566 15774 39618
rect 24210 39566 24222 39618
rect 24274 39566 24286 39618
rect 24670 39554 24722 39566
rect 12114 39454 12126 39506
rect 12178 39454 12190 39506
rect 16482 39454 16494 39506
rect 16546 39454 16558 39506
rect 23426 39454 23438 39506
rect 23490 39454 23502 39506
rect 13582 39394 13634 39406
rect 13582 39330 13634 39342
rect 15374 39394 15426 39406
rect 15374 39330 15426 39342
rect 1344 39226 39984 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 39984 39226
rect 1344 39140 39984 39174
rect 12126 39058 12178 39070
rect 16482 39006 16494 39058
rect 16546 39006 16558 39058
rect 12126 38994 12178 39006
rect 12014 38946 12066 38958
rect 17726 38946 17778 38958
rect 15026 38894 15038 38946
rect 15090 38894 15102 38946
rect 16594 38894 16606 38946
rect 16658 38894 16670 38946
rect 12014 38882 12066 38894
rect 17726 38882 17778 38894
rect 18286 38946 18338 38958
rect 18286 38882 18338 38894
rect 22878 38946 22930 38958
rect 22878 38882 22930 38894
rect 12686 38834 12738 38846
rect 18062 38834 18114 38846
rect 13122 38782 13134 38834
rect 13186 38782 13198 38834
rect 17378 38782 17390 38834
rect 17442 38782 17454 38834
rect 12686 38770 12738 38782
rect 18062 38770 18114 38782
rect 18174 38834 18226 38846
rect 18174 38770 18226 38782
rect 18734 38834 18786 38846
rect 20974 38834 21026 38846
rect 20178 38782 20190 38834
rect 20242 38782 20254 38834
rect 20402 38782 20414 38834
rect 20466 38782 20478 38834
rect 21634 38782 21646 38834
rect 21698 38782 21710 38834
rect 18734 38770 18786 38782
rect 20974 38770 21026 38782
rect 11678 38722 11730 38734
rect 11678 38658 11730 38670
rect 13582 38722 13634 38734
rect 17614 38722 17666 38734
rect 14690 38670 14702 38722
rect 14754 38670 14766 38722
rect 13582 38658 13634 38670
rect 17614 38658 17666 38670
rect 20638 38722 20690 38734
rect 21298 38670 21310 38722
rect 21362 38670 21374 38722
rect 22418 38670 22430 38722
rect 22482 38670 22494 38722
rect 20638 38658 20690 38670
rect 12238 38610 12290 38622
rect 12238 38546 12290 38558
rect 1344 38442 39984 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 39984 38442
rect 1344 38356 39984 38390
rect 18174 38274 18226 38286
rect 18174 38210 18226 38222
rect 22654 38274 22706 38286
rect 22654 38210 22706 38222
rect 10558 38162 10610 38174
rect 9986 38110 9998 38162
rect 10050 38110 10062 38162
rect 10558 38098 10610 38110
rect 13806 38162 13858 38174
rect 13806 38098 13858 38110
rect 17166 38162 17218 38174
rect 17166 38098 17218 38110
rect 20638 38162 20690 38174
rect 22318 38162 22370 38174
rect 21858 38110 21870 38162
rect 21922 38110 21934 38162
rect 20638 38098 20690 38110
rect 22318 38098 22370 38110
rect 13918 38050 13970 38062
rect 16158 38050 16210 38062
rect 9650 37998 9662 38050
rect 9714 37998 9726 38050
rect 11330 37998 11342 38050
rect 11394 37998 11406 38050
rect 14130 37998 14142 38050
rect 14194 37998 14206 38050
rect 15922 37998 15934 38050
rect 15986 37998 15998 38050
rect 13918 37986 13970 37998
rect 16158 37986 16210 37998
rect 16382 38050 16434 38062
rect 18398 38050 18450 38062
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 16382 37986 16434 37998
rect 18398 37986 18450 37998
rect 18734 38050 18786 38062
rect 18734 37986 18786 37998
rect 19854 38050 19906 38062
rect 19854 37986 19906 37998
rect 21534 38050 21586 38062
rect 22642 37998 22654 38050
rect 22706 37998 22718 38050
rect 21534 37986 21586 37998
rect 12238 37938 12290 37950
rect 11554 37886 11566 37938
rect 11618 37886 11630 37938
rect 12238 37874 12290 37886
rect 12350 37938 12402 37950
rect 12350 37874 12402 37886
rect 12686 37938 12738 37950
rect 12686 37874 12738 37886
rect 13470 37938 13522 37950
rect 13470 37874 13522 37886
rect 16606 37938 16658 37950
rect 16606 37874 16658 37886
rect 18622 37938 18674 37950
rect 18622 37874 18674 37886
rect 18958 37938 19010 37950
rect 20078 37938 20130 37950
rect 19282 37886 19294 37938
rect 19346 37886 19358 37938
rect 18958 37874 19010 37886
rect 20078 37874 20130 37886
rect 20190 37938 20242 37950
rect 20190 37874 20242 37886
rect 21310 37938 21362 37950
rect 21310 37874 21362 37886
rect 21870 37938 21922 37950
rect 21870 37874 21922 37886
rect 12798 37826 12850 37838
rect 12798 37762 12850 37774
rect 13022 37826 13074 37838
rect 13022 37762 13074 37774
rect 13694 37826 13746 37838
rect 13694 37762 13746 37774
rect 16270 37826 16322 37838
rect 16270 37762 16322 37774
rect 19630 37826 19682 37838
rect 19630 37762 19682 37774
rect 20526 37826 20578 37838
rect 20526 37762 20578 37774
rect 21758 37826 21810 37838
rect 21758 37762 21810 37774
rect 23102 37826 23154 37838
rect 23102 37762 23154 37774
rect 1344 37658 39984 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 39984 37658
rect 1344 37572 39984 37606
rect 13470 37490 13522 37502
rect 13470 37426 13522 37438
rect 13582 37490 13634 37502
rect 17502 37490 17554 37502
rect 16818 37438 16830 37490
rect 16882 37438 16894 37490
rect 13582 37426 13634 37438
rect 17502 37426 17554 37438
rect 18062 37490 18114 37502
rect 18062 37426 18114 37438
rect 18174 37490 18226 37502
rect 18174 37426 18226 37438
rect 17390 37378 17442 37390
rect 17390 37314 17442 37326
rect 17614 37378 17666 37390
rect 17614 37314 17666 37326
rect 24446 37378 24498 37390
rect 24446 37314 24498 37326
rect 28814 37378 28866 37390
rect 28814 37314 28866 37326
rect 13358 37266 13410 37278
rect 14366 37266 14418 37278
rect 13906 37214 13918 37266
rect 13970 37214 13982 37266
rect 13358 37202 13410 37214
rect 14366 37202 14418 37214
rect 16494 37266 16546 37278
rect 16494 37202 16546 37214
rect 18286 37266 18338 37278
rect 18286 37202 18338 37214
rect 18734 37266 18786 37278
rect 28242 37214 28254 37266
rect 28306 37214 28318 37266
rect 18734 37202 18786 37214
rect 19070 37154 19122 37166
rect 19070 37090 19122 37102
rect 20414 37154 20466 37166
rect 20414 37090 20466 37102
rect 22206 37154 22258 37166
rect 22206 37090 22258 37102
rect 23550 37154 23602 37166
rect 23550 37090 23602 37102
rect 24558 37154 24610 37166
rect 25330 37102 25342 37154
rect 25394 37102 25406 37154
rect 27570 37102 27582 37154
rect 27634 37102 27646 37154
rect 24558 37090 24610 37102
rect 24670 37042 24722 37054
rect 24670 36978 24722 36990
rect 1344 36874 39984 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 39984 36874
rect 1344 36788 39984 36822
rect 17726 36594 17778 36606
rect 17726 36530 17778 36542
rect 21422 36594 21474 36606
rect 26238 36594 26290 36606
rect 25218 36542 25230 36594
rect 25282 36542 25294 36594
rect 21422 36530 21474 36542
rect 26238 36530 26290 36542
rect 13694 36482 13746 36494
rect 13694 36418 13746 36430
rect 21646 36482 21698 36494
rect 23886 36482 23938 36494
rect 25342 36482 25394 36494
rect 21970 36430 21982 36482
rect 22034 36430 22046 36482
rect 22306 36430 22318 36482
rect 22370 36430 22382 36482
rect 23426 36430 23438 36482
rect 23490 36430 23502 36482
rect 24098 36430 24110 36482
rect 24162 36430 24174 36482
rect 21646 36418 21698 36430
rect 23886 36418 23938 36430
rect 25342 36418 25394 36430
rect 13470 36370 13522 36382
rect 13470 36306 13522 36318
rect 14030 36370 14082 36382
rect 24782 36370 24834 36382
rect 23314 36318 23326 36370
rect 23378 36318 23390 36370
rect 14030 36306 14082 36318
rect 24782 36306 24834 36318
rect 25566 36370 25618 36382
rect 25566 36306 25618 36318
rect 25790 36370 25842 36382
rect 25790 36306 25842 36318
rect 12574 36258 12626 36270
rect 12574 36194 12626 36206
rect 13806 36258 13858 36270
rect 25230 36258 25282 36270
rect 22418 36206 22430 36258
rect 22482 36206 22494 36258
rect 13806 36194 13858 36206
rect 25230 36194 25282 36206
rect 33070 36258 33122 36270
rect 33742 36258 33794 36270
rect 33394 36206 33406 36258
rect 33458 36206 33470 36258
rect 33070 36194 33122 36206
rect 33742 36194 33794 36206
rect 1344 36090 39984 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 39984 36090
rect 1344 36004 39984 36038
rect 24098 35870 24110 35922
rect 24162 35870 24174 35922
rect 12126 35810 12178 35822
rect 12126 35746 12178 35758
rect 14478 35810 14530 35822
rect 14478 35746 14530 35758
rect 14702 35810 14754 35822
rect 22766 35810 22818 35822
rect 19842 35758 19854 35810
rect 19906 35758 19918 35810
rect 14702 35746 14754 35758
rect 22766 35746 22818 35758
rect 13694 35698 13746 35710
rect 6178 35646 6190 35698
rect 6242 35646 6254 35698
rect 13234 35646 13246 35698
rect 13298 35646 13310 35698
rect 13694 35634 13746 35646
rect 14142 35698 14194 35710
rect 14142 35634 14194 35646
rect 14254 35698 14306 35710
rect 14254 35634 14306 35646
rect 19518 35698 19570 35710
rect 22194 35646 22206 35698
rect 22258 35646 22270 35698
rect 24322 35646 24334 35698
rect 24386 35646 24398 35698
rect 28242 35646 28254 35698
rect 28306 35646 28318 35698
rect 19518 35634 19570 35646
rect 9662 35586 9714 35598
rect 6850 35534 6862 35586
rect 6914 35534 6926 35586
rect 8978 35534 8990 35586
rect 9042 35534 9054 35586
rect 9662 35522 9714 35534
rect 12350 35586 12402 35598
rect 14366 35586 14418 35598
rect 23214 35586 23266 35598
rect 31502 35586 31554 35598
rect 13346 35534 13358 35586
rect 13410 35534 13422 35586
rect 21858 35534 21870 35586
rect 21922 35534 21934 35586
rect 28914 35534 28926 35586
rect 28978 35534 28990 35586
rect 31042 35534 31054 35586
rect 31106 35534 31118 35586
rect 12350 35522 12402 35534
rect 14366 35522 14418 35534
rect 23214 35522 23266 35534
rect 31502 35522 31554 35534
rect 12014 35474 12066 35486
rect 12014 35410 12066 35422
rect 1344 35306 39984 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 39984 35306
rect 1344 35220 39984 35254
rect 11566 35138 11618 35150
rect 11566 35074 11618 35086
rect 9662 35026 9714 35038
rect 17502 35026 17554 35038
rect 28366 35026 28418 35038
rect 6402 34974 6414 35026
rect 6466 34974 6478 35026
rect 8530 34974 8542 35026
rect 8594 34974 8606 35026
rect 12114 34974 12126 35026
rect 12178 34974 12190 35026
rect 14242 34974 14254 35026
rect 14306 34974 14318 35026
rect 22866 34974 22878 35026
rect 22930 34974 22942 35026
rect 34402 34974 34414 35026
rect 34466 34974 34478 35026
rect 35746 34974 35758 35026
rect 35810 34974 35822 35026
rect 9662 34962 9714 34974
rect 17502 34962 17554 34974
rect 28366 34962 28418 34974
rect 8878 34914 8930 34926
rect 14926 34914 14978 34926
rect 5618 34862 5630 34914
rect 5682 34862 5694 34914
rect 11554 34862 11566 34914
rect 11618 34862 11630 34914
rect 12450 34862 12462 34914
rect 12514 34862 12526 34914
rect 14130 34862 14142 34914
rect 14194 34862 14206 34914
rect 8878 34850 8930 34862
rect 14926 34850 14978 34862
rect 17278 34914 17330 34926
rect 17938 34862 17950 34914
rect 18002 34862 18014 34914
rect 34738 34862 34750 34914
rect 34802 34862 34814 34914
rect 17278 34850 17330 34862
rect 11230 34802 11282 34814
rect 11230 34738 11282 34750
rect 12910 34802 12962 34814
rect 12910 34738 12962 34750
rect 13470 34802 13522 34814
rect 13470 34738 13522 34750
rect 14814 34802 14866 34814
rect 34078 34802 34130 34814
rect 17826 34750 17838 34802
rect 17890 34750 17902 34802
rect 18386 34750 18398 34802
rect 18450 34750 18462 34802
rect 14814 34738 14866 34750
rect 34078 34738 34130 34750
rect 35422 34802 35474 34814
rect 35422 34738 35474 34750
rect 23326 34690 23378 34702
rect 9202 34638 9214 34690
rect 9266 34638 9278 34690
rect 16930 34638 16942 34690
rect 16994 34638 17006 34690
rect 23326 34626 23378 34638
rect 29374 34690 29426 34702
rect 29374 34626 29426 34638
rect 35646 34690 35698 34702
rect 35646 34626 35698 34638
rect 1344 34522 39984 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 39984 34522
rect 1344 34436 39984 34470
rect 12462 34354 12514 34366
rect 17614 34354 17666 34366
rect 12786 34302 12798 34354
rect 12850 34302 12862 34354
rect 12462 34290 12514 34302
rect 17614 34290 17666 34302
rect 18286 34354 18338 34366
rect 19742 34354 19794 34366
rect 18610 34302 18622 34354
rect 18674 34302 18686 34354
rect 18286 34290 18338 34302
rect 19742 34290 19794 34302
rect 28926 34354 28978 34366
rect 28926 34290 28978 34302
rect 29150 34354 29202 34366
rect 29150 34290 29202 34302
rect 17838 34242 17890 34254
rect 30830 34242 30882 34254
rect 14690 34190 14702 34242
rect 14754 34190 14766 34242
rect 16146 34190 16158 34242
rect 16210 34190 16222 34242
rect 29586 34190 29598 34242
rect 29650 34190 29662 34242
rect 17838 34178 17890 34190
rect 30830 34178 30882 34190
rect 32174 34242 32226 34254
rect 36530 34190 36542 34242
rect 36594 34190 36606 34242
rect 32174 34178 32226 34190
rect 14142 34130 14194 34142
rect 17278 34130 17330 34142
rect 19182 34130 19234 34142
rect 13458 34078 13470 34130
rect 13522 34078 13534 34130
rect 13906 34078 13918 34130
rect 13970 34078 13982 34130
rect 14578 34078 14590 34130
rect 14642 34078 14654 34130
rect 15586 34078 15598 34130
rect 15650 34078 15662 34130
rect 18834 34078 18846 34130
rect 18898 34078 18910 34130
rect 14142 34066 14194 34078
rect 17278 34066 17330 34078
rect 19182 34066 19234 34078
rect 19630 34130 19682 34142
rect 19630 34066 19682 34078
rect 19854 34130 19906 34142
rect 29262 34130 29314 34142
rect 25330 34078 25342 34130
rect 25394 34078 25406 34130
rect 19854 34066 19906 34078
rect 29262 34066 29314 34078
rect 29934 34130 29986 34142
rect 29934 34066 29986 34078
rect 30270 34130 30322 34142
rect 30270 34066 30322 34078
rect 30606 34130 30658 34142
rect 34078 34130 34130 34142
rect 31714 34078 31726 34130
rect 31778 34078 31790 34130
rect 37202 34078 37214 34130
rect 37266 34078 37278 34130
rect 30606 34066 30658 34078
rect 34078 34066 34130 34078
rect 10446 34018 10498 34030
rect 20974 34018 21026 34030
rect 28814 34018 28866 34030
rect 15922 33966 15934 34018
rect 15986 33966 15998 34018
rect 26002 33966 26014 34018
rect 26066 33966 26078 34018
rect 28130 33966 28142 34018
rect 28194 33966 28206 34018
rect 10446 33954 10498 33966
rect 20974 33954 21026 33966
rect 28814 33954 28866 33966
rect 30382 34018 30434 34030
rect 31266 33966 31278 34018
rect 31330 33966 31342 34018
rect 34402 33966 34414 34018
rect 34466 33966 34478 34018
rect 30382 33954 30434 33966
rect 10558 33906 10610 33918
rect 10558 33842 10610 33854
rect 17502 33906 17554 33918
rect 17502 33842 17554 33854
rect 1344 33738 39984 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 39984 33738
rect 1344 33652 39984 33686
rect 14030 33570 14082 33582
rect 14030 33506 14082 33518
rect 9214 33458 9266 33470
rect 7970 33406 7982 33458
rect 8034 33406 8046 33458
rect 9214 33394 9266 33406
rect 15038 33458 15090 33470
rect 15038 33394 15090 33406
rect 17390 33458 17442 33470
rect 25566 33458 25618 33470
rect 19618 33406 19630 33458
rect 19682 33406 19694 33458
rect 17390 33394 17442 33406
rect 25566 33394 25618 33406
rect 25678 33458 25730 33470
rect 26114 33406 26126 33458
rect 26178 33406 26190 33458
rect 31154 33406 31166 33458
rect 31218 33406 31230 33458
rect 25678 33394 25730 33406
rect 9998 33346 10050 33358
rect 10894 33346 10946 33358
rect 15710 33346 15762 33358
rect 7298 33294 7310 33346
rect 7362 33294 7374 33346
rect 9314 33294 9326 33346
rect 9378 33294 9390 33346
rect 10434 33294 10446 33346
rect 10498 33294 10510 33346
rect 14242 33294 14254 33346
rect 14306 33294 14318 33346
rect 14914 33294 14926 33346
rect 14978 33294 14990 33346
rect 9998 33282 10050 33294
rect 10894 33282 10946 33294
rect 15710 33282 15762 33294
rect 16270 33346 16322 33358
rect 16270 33282 16322 33294
rect 16942 33346 16994 33358
rect 16942 33282 16994 33294
rect 17278 33346 17330 33358
rect 17278 33282 17330 33294
rect 17502 33346 17554 33358
rect 20078 33346 20130 33358
rect 18610 33294 18622 33346
rect 18674 33294 18686 33346
rect 19058 33294 19070 33346
rect 19122 33294 19134 33346
rect 17502 33282 17554 33294
rect 20078 33282 20130 33294
rect 20302 33346 20354 33358
rect 20302 33282 20354 33294
rect 20526 33346 20578 33358
rect 20526 33282 20578 33294
rect 21534 33346 21586 33358
rect 34862 33346 34914 33358
rect 26674 33294 26686 33346
rect 26738 33294 26750 33346
rect 29138 33294 29150 33346
rect 29202 33294 29214 33346
rect 35298 33294 35310 33346
rect 35362 33294 35374 33346
rect 21534 33282 21586 33294
rect 34862 33282 34914 33294
rect 8206 33234 8258 33246
rect 8206 33170 8258 33182
rect 9102 33234 9154 33246
rect 9102 33170 9154 33182
rect 9550 33234 9602 33246
rect 9550 33170 9602 33182
rect 11342 33234 11394 33246
rect 11342 33170 11394 33182
rect 11454 33234 11506 33246
rect 11454 33170 11506 33182
rect 12574 33234 12626 33246
rect 12574 33170 12626 33182
rect 12798 33234 12850 33246
rect 12798 33170 12850 33182
rect 20638 33234 20690 33246
rect 20638 33170 20690 33182
rect 28590 33234 28642 33246
rect 28590 33170 28642 33182
rect 35758 33234 35810 33246
rect 35758 33170 35810 33182
rect 11118 33122 11170 33134
rect 11118 33058 11170 33070
rect 12686 33122 12738 33134
rect 12686 33058 12738 33070
rect 15598 33122 15650 33134
rect 15598 33058 15650 33070
rect 15822 33122 15874 33134
rect 15822 33058 15874 33070
rect 16718 33122 16770 33134
rect 16718 33058 16770 33070
rect 21310 33122 21362 33134
rect 21310 33058 21362 33070
rect 21422 33122 21474 33134
rect 21422 33058 21474 33070
rect 21758 33122 21810 33134
rect 21758 33058 21810 33070
rect 25454 33122 25506 33134
rect 25454 33058 25506 33070
rect 26126 33122 26178 33134
rect 26126 33058 26178 33070
rect 26238 33122 26290 33134
rect 26238 33058 26290 33070
rect 26462 33122 26514 33134
rect 26462 33058 26514 33070
rect 28142 33122 28194 33134
rect 28142 33058 28194 33070
rect 28254 33122 28306 33134
rect 28254 33058 28306 33070
rect 28478 33122 28530 33134
rect 28478 33058 28530 33070
rect 1344 32954 39984 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 39984 32954
rect 1344 32868 39984 32902
rect 17502 32786 17554 32798
rect 17502 32722 17554 32734
rect 17726 32786 17778 32798
rect 17726 32722 17778 32734
rect 18062 32786 18114 32798
rect 18062 32722 18114 32734
rect 18286 32786 18338 32798
rect 18286 32722 18338 32734
rect 19630 32786 19682 32798
rect 19630 32722 19682 32734
rect 23550 32786 23602 32798
rect 23550 32722 23602 32734
rect 25230 32786 25282 32798
rect 25230 32722 25282 32734
rect 30382 32786 30434 32798
rect 30382 32722 30434 32734
rect 32958 32786 33010 32798
rect 32958 32722 33010 32734
rect 33182 32786 33234 32798
rect 33182 32722 33234 32734
rect 35310 32786 35362 32798
rect 35310 32722 35362 32734
rect 36318 32786 36370 32798
rect 36318 32722 36370 32734
rect 26798 32674 26850 32686
rect 35086 32674 35138 32686
rect 11778 32622 11790 32674
rect 11842 32622 11854 32674
rect 22306 32622 22318 32674
rect 22370 32622 22382 32674
rect 25554 32622 25566 32674
rect 25618 32622 25630 32674
rect 26114 32622 26126 32674
rect 26178 32622 26190 32674
rect 28690 32622 28702 32674
rect 28754 32622 28766 32674
rect 26798 32610 26850 32622
rect 35086 32610 35138 32622
rect 17390 32562 17442 32574
rect 15474 32510 15486 32562
rect 15538 32510 15550 32562
rect 17390 32498 17442 32510
rect 17950 32562 18002 32574
rect 26462 32562 26514 32574
rect 29486 32562 29538 32574
rect 19842 32510 19854 32562
rect 19906 32510 19918 32562
rect 23090 32510 23102 32562
rect 23154 32510 23166 32562
rect 27458 32510 27470 32562
rect 27522 32510 27534 32562
rect 28130 32510 28142 32562
rect 28194 32510 28206 32562
rect 17950 32498 18002 32510
rect 26462 32498 26514 32510
rect 29486 32498 29538 32510
rect 29822 32562 29874 32574
rect 30270 32562 30322 32574
rect 30146 32510 30158 32562
rect 30210 32510 30222 32562
rect 29822 32498 29874 32510
rect 30270 32498 30322 32510
rect 30494 32562 30546 32574
rect 30494 32498 30546 32510
rect 31278 32562 31330 32574
rect 31278 32498 31330 32510
rect 31838 32562 31890 32574
rect 31838 32498 31890 32510
rect 32062 32562 32114 32574
rect 32062 32498 32114 32510
rect 33294 32562 33346 32574
rect 33294 32498 33346 32510
rect 34526 32562 34578 32574
rect 34526 32498 34578 32510
rect 35422 32562 35474 32574
rect 35422 32498 35474 32510
rect 35534 32562 35586 32574
rect 35746 32510 35758 32562
rect 35810 32510 35822 32562
rect 36642 32510 36654 32562
rect 36706 32510 36718 32562
rect 35534 32498 35586 32510
rect 15934 32450 15986 32462
rect 15934 32386 15986 32398
rect 19294 32450 19346 32462
rect 31502 32450 31554 32462
rect 20178 32398 20190 32450
rect 20242 32398 20254 32450
rect 19294 32386 19346 32398
rect 31502 32386 31554 32398
rect 34750 32450 34802 32462
rect 37426 32398 37438 32450
rect 37490 32398 37502 32450
rect 39554 32398 39566 32450
rect 39618 32398 39630 32450
rect 34750 32386 34802 32398
rect 19518 32338 19570 32350
rect 19518 32274 19570 32286
rect 30942 32338 30994 32350
rect 32386 32286 32398 32338
rect 32450 32286 32462 32338
rect 34178 32286 34190 32338
rect 34242 32286 34254 32338
rect 30942 32274 30994 32286
rect 1344 32170 39984 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 39984 32170
rect 1344 32084 39984 32118
rect 30830 32002 30882 32014
rect 30830 31938 30882 31950
rect 37326 32002 37378 32014
rect 37326 31938 37378 31950
rect 12574 31890 12626 31902
rect 8418 31838 8430 31890
rect 8482 31838 8494 31890
rect 10434 31838 10446 31890
rect 10498 31838 10510 31890
rect 12574 31826 12626 31838
rect 17166 31890 17218 31902
rect 36990 31890 37042 31902
rect 35522 31838 35534 31890
rect 35586 31838 35598 31890
rect 17166 31826 17218 31838
rect 36990 31826 37042 31838
rect 11566 31778 11618 31790
rect 8866 31726 8878 31778
rect 8930 31726 8942 31778
rect 10098 31726 10110 31778
rect 10162 31726 10174 31778
rect 11566 31714 11618 31726
rect 12126 31778 12178 31790
rect 12126 31714 12178 31726
rect 14254 31778 14306 31790
rect 14254 31714 14306 31726
rect 14926 31778 14978 31790
rect 14926 31714 14978 31726
rect 16382 31778 16434 31790
rect 16382 31714 16434 31726
rect 16942 31778 16994 31790
rect 16942 31714 16994 31726
rect 17726 31778 17778 31790
rect 31502 31778 31554 31790
rect 20514 31726 20526 31778
rect 20578 31726 20590 31778
rect 31154 31726 31166 31778
rect 31218 31726 31230 31778
rect 17726 31714 17778 31726
rect 31502 31714 31554 31726
rect 31950 31778 32002 31790
rect 31950 31714 32002 31726
rect 34414 31778 34466 31790
rect 35074 31726 35086 31778
rect 35138 31726 35150 31778
rect 34414 31714 34466 31726
rect 9326 31666 9378 31678
rect 9326 31602 9378 31614
rect 9662 31666 9714 31678
rect 9662 31602 9714 31614
rect 12014 31666 12066 31678
rect 12014 31602 12066 31614
rect 14814 31666 14866 31678
rect 14814 31602 14866 31614
rect 16158 31666 16210 31678
rect 16158 31602 16210 31614
rect 17950 31666 18002 31678
rect 17950 31602 18002 31614
rect 18062 31666 18114 31678
rect 35534 31666 35586 31678
rect 20290 31614 20302 31666
rect 20354 31614 20366 31666
rect 21746 31614 21758 31666
rect 21810 31614 21822 31666
rect 34738 31614 34750 31666
rect 34802 31614 34814 31666
rect 18062 31602 18114 31614
rect 35534 31602 35586 31614
rect 11790 31554 11842 31566
rect 11218 31502 11230 31554
rect 11282 31502 11294 31554
rect 11790 31490 11842 31502
rect 14702 31554 14754 31566
rect 14702 31490 14754 31502
rect 16270 31554 16322 31566
rect 16270 31490 16322 31502
rect 16606 31554 16658 31566
rect 16606 31490 16658 31502
rect 17278 31554 17330 31566
rect 17278 31490 17330 31502
rect 17502 31554 17554 31566
rect 17502 31490 17554 31502
rect 18622 31554 18674 31566
rect 18622 31490 18674 31502
rect 18958 31554 19010 31566
rect 18958 31490 19010 31502
rect 22094 31554 22146 31566
rect 22094 31490 22146 31502
rect 30942 31554 30994 31566
rect 30942 31490 30994 31502
rect 31614 31554 31666 31566
rect 31614 31490 31666 31502
rect 31838 31554 31890 31566
rect 31838 31490 31890 31502
rect 35310 31554 35362 31566
rect 35310 31490 35362 31502
rect 35646 31554 35698 31566
rect 35646 31490 35698 31502
rect 37214 31554 37266 31566
rect 37214 31490 37266 31502
rect 1344 31386 39984 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 39984 31386
rect 1344 31300 39984 31334
rect 16942 31218 16994 31230
rect 14018 31166 14030 31218
rect 14082 31166 14094 31218
rect 16942 31154 16994 31166
rect 29710 31218 29762 31230
rect 29710 31154 29762 31166
rect 32286 31218 32338 31230
rect 33170 31166 33182 31218
rect 33234 31166 33246 31218
rect 35858 31166 35870 31218
rect 35922 31166 35934 31218
rect 32286 31154 32338 31166
rect 7198 31106 7250 31118
rect 17390 31106 17442 31118
rect 9650 31054 9662 31106
rect 9714 31054 9726 31106
rect 7198 31042 7250 31054
rect 17390 31042 17442 31054
rect 18846 31106 18898 31118
rect 18846 31042 18898 31054
rect 23214 31106 23266 31118
rect 23214 31042 23266 31054
rect 29934 31106 29986 31118
rect 29934 31042 29986 31054
rect 30270 31106 30322 31118
rect 34290 31054 34302 31106
rect 34354 31054 34366 31106
rect 37762 31054 37774 31106
rect 37826 31054 37838 31106
rect 30270 31042 30322 31054
rect 8766 30994 8818 31006
rect 2818 30942 2830 30994
rect 2882 30942 2894 30994
rect 6626 30942 6638 30994
rect 6690 30942 6702 30994
rect 8530 30942 8542 30994
rect 8594 30942 8606 30994
rect 8766 30930 8818 30942
rect 8990 30994 9042 31006
rect 8990 30930 9042 30942
rect 9550 30994 9602 31006
rect 9550 30930 9602 30942
rect 9886 30994 9938 31006
rect 16046 30994 16098 31006
rect 10098 30942 10110 30994
rect 10162 30942 10174 30994
rect 13794 30942 13806 30994
rect 13858 30942 13870 30994
rect 9886 30930 9938 30942
rect 16046 30930 16098 30942
rect 16270 30994 16322 31006
rect 16270 30930 16322 30942
rect 16494 30994 16546 31006
rect 22654 30994 22706 31006
rect 29598 30994 29650 31006
rect 17602 30942 17614 30994
rect 17666 30942 17678 30994
rect 17826 30942 17838 30994
rect 17890 30942 17902 30994
rect 23650 30942 23662 30994
rect 23714 30942 23726 30994
rect 16494 30930 16546 30942
rect 22654 30930 22706 30942
rect 29598 30930 29650 30942
rect 30382 30994 30434 31006
rect 32062 30994 32114 31006
rect 31826 30942 31838 30994
rect 31890 30942 31902 30994
rect 30382 30930 30434 30942
rect 32062 30930 32114 30942
rect 32398 30994 32450 31006
rect 36542 30994 36594 31006
rect 33394 30942 33406 30994
rect 33458 30942 33470 30994
rect 35746 30942 35758 30994
rect 35810 30942 35822 30994
rect 36978 30942 36990 30994
rect 37042 30942 37054 30994
rect 37538 30942 37550 30994
rect 37602 30942 37614 30994
rect 32398 30930 32450 30942
rect 36542 30930 36594 30942
rect 24110 30882 24162 30894
rect 3602 30830 3614 30882
rect 3666 30830 3678 30882
rect 5730 30830 5742 30882
rect 5794 30830 5806 30882
rect 6402 30830 6414 30882
rect 6466 30830 6478 30882
rect 24110 30818 24162 30830
rect 32174 30882 32226 30894
rect 34066 30830 34078 30882
rect 34130 30830 34142 30882
rect 32174 30818 32226 30830
rect 10558 30770 10610 30782
rect 10558 30706 10610 30718
rect 18734 30770 18786 30782
rect 18734 30706 18786 30718
rect 30270 30770 30322 30782
rect 30270 30706 30322 30718
rect 1344 30602 39984 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 39984 30602
rect 1344 30516 39984 30550
rect 13918 30434 13970 30446
rect 13918 30370 13970 30382
rect 27806 30434 27858 30446
rect 27806 30370 27858 30382
rect 32174 30434 32226 30446
rect 32174 30370 32226 30382
rect 23662 30322 23714 30334
rect 27694 30322 27746 30334
rect 11778 30270 11790 30322
rect 11842 30270 11854 30322
rect 23986 30270 23998 30322
rect 24050 30270 24062 30322
rect 26450 30270 26462 30322
rect 26514 30270 26526 30322
rect 23662 30258 23714 30270
rect 27694 30258 27746 30270
rect 36318 30322 36370 30334
rect 36318 30258 36370 30270
rect 37326 30322 37378 30334
rect 37326 30258 37378 30270
rect 5966 30210 6018 30222
rect 5966 30146 6018 30158
rect 6414 30210 6466 30222
rect 8654 30210 8706 30222
rect 8082 30158 8094 30210
rect 8146 30158 8158 30210
rect 6414 30146 6466 30158
rect 8654 30146 8706 30158
rect 8766 30210 8818 30222
rect 8766 30146 8818 30158
rect 10222 30210 10274 30222
rect 14366 30210 14418 30222
rect 10546 30158 10558 30210
rect 10610 30158 10622 30210
rect 11666 30158 11678 30210
rect 11730 30158 11742 30210
rect 10222 30146 10274 30158
rect 14366 30146 14418 30158
rect 14926 30210 14978 30222
rect 14926 30146 14978 30158
rect 17054 30210 17106 30222
rect 17054 30146 17106 30158
rect 17502 30210 17554 30222
rect 17502 30146 17554 30158
rect 18398 30210 18450 30222
rect 27470 30210 27522 30222
rect 31166 30210 31218 30222
rect 24210 30158 24222 30210
rect 24274 30158 24286 30210
rect 26114 30158 26126 30210
rect 26178 30158 26190 30210
rect 29922 30158 29934 30210
rect 29986 30158 29998 30210
rect 30930 30158 30942 30210
rect 30994 30158 31006 30210
rect 18398 30146 18450 30158
rect 27470 30146 27522 30158
rect 31166 30146 31218 30158
rect 31390 30210 31442 30222
rect 31390 30146 31442 30158
rect 31502 30210 31554 30222
rect 36878 30210 36930 30222
rect 35858 30158 35870 30210
rect 35922 30158 35934 30210
rect 31502 30146 31554 30158
rect 36878 30146 36930 30158
rect 37550 30210 37602 30222
rect 37550 30146 37602 30158
rect 37662 30210 37714 30222
rect 37662 30146 37714 30158
rect 10782 30098 10834 30110
rect 10782 30034 10834 30046
rect 11230 30098 11282 30110
rect 11230 30034 11282 30046
rect 13694 30098 13746 30110
rect 13694 30034 13746 30046
rect 14478 30098 14530 30110
rect 14478 30034 14530 30046
rect 17390 30098 17442 30110
rect 17390 30034 17442 30046
rect 18174 30098 18226 30110
rect 18174 30034 18226 30046
rect 18734 30098 18786 30110
rect 18734 30034 18786 30046
rect 27022 30098 27074 30110
rect 27022 30034 27074 30046
rect 27358 30098 27410 30110
rect 31950 30098 32002 30110
rect 39230 30098 39282 30110
rect 30146 30046 30158 30098
rect 30210 30046 30222 30098
rect 38658 30046 38670 30098
rect 38722 30046 38734 30098
rect 27358 30034 27410 30046
rect 31950 30034 32002 30046
rect 39230 30034 39282 30046
rect 39342 30098 39394 30110
rect 39342 30034 39394 30046
rect 10894 29986 10946 29998
rect 6738 29934 6750 29986
rect 6802 29934 6814 29986
rect 10894 29922 10946 29934
rect 13806 29986 13858 29998
rect 13806 29922 13858 29934
rect 14254 29986 14306 29998
rect 14254 29922 14306 29934
rect 16718 29986 16770 29998
rect 16718 29922 16770 29934
rect 17166 29986 17218 29998
rect 17166 29922 17218 29934
rect 18398 29986 18450 29998
rect 18398 29922 18450 29934
rect 24894 29986 24946 29998
rect 24894 29922 24946 29934
rect 31278 29986 31330 29998
rect 36206 29986 36258 29998
rect 32498 29934 32510 29986
rect 32562 29934 32574 29986
rect 31278 29922 31330 29934
rect 36206 29922 36258 29934
rect 36430 29986 36482 29998
rect 36430 29922 36482 29934
rect 39006 29986 39058 29998
rect 39006 29922 39058 29934
rect 1344 29818 39984 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 39984 29818
rect 1344 29732 39984 29766
rect 5182 29650 5234 29662
rect 5182 29586 5234 29598
rect 10446 29650 10498 29662
rect 10446 29586 10498 29598
rect 10558 29650 10610 29662
rect 10558 29586 10610 29598
rect 11342 29650 11394 29662
rect 11342 29586 11394 29598
rect 13918 29650 13970 29662
rect 13918 29586 13970 29598
rect 14478 29650 14530 29662
rect 14478 29586 14530 29598
rect 17390 29650 17442 29662
rect 17390 29586 17442 29598
rect 26798 29650 26850 29662
rect 26798 29586 26850 29598
rect 28254 29650 28306 29662
rect 28254 29586 28306 29598
rect 31390 29650 31442 29662
rect 31390 29586 31442 29598
rect 36878 29650 36930 29662
rect 36878 29586 36930 29598
rect 36990 29650 37042 29662
rect 36990 29586 37042 29598
rect 11566 29538 11618 29550
rect 11566 29474 11618 29486
rect 17614 29538 17666 29550
rect 17614 29474 17666 29486
rect 17726 29538 17778 29550
rect 17726 29474 17778 29486
rect 18174 29538 18226 29550
rect 18174 29474 18226 29486
rect 19070 29538 19122 29550
rect 19070 29474 19122 29486
rect 19182 29538 19234 29550
rect 26462 29538 26514 29550
rect 26338 29486 26350 29538
rect 26402 29486 26414 29538
rect 19182 29474 19234 29486
rect 26462 29474 26514 29486
rect 26574 29538 26626 29550
rect 26574 29474 26626 29486
rect 26686 29538 26738 29550
rect 26686 29474 26738 29486
rect 28366 29538 28418 29550
rect 28366 29474 28418 29486
rect 31166 29538 31218 29550
rect 31166 29474 31218 29486
rect 37774 29538 37826 29550
rect 37774 29474 37826 29486
rect 37998 29538 38050 29550
rect 37998 29474 38050 29486
rect 10334 29426 10386 29438
rect 1922 29374 1934 29426
rect 1986 29374 1998 29426
rect 10098 29374 10110 29426
rect 10162 29374 10174 29426
rect 10334 29362 10386 29374
rect 10670 29426 10722 29438
rect 10670 29362 10722 29374
rect 11006 29426 11058 29438
rect 11006 29362 11058 29374
rect 14030 29426 14082 29438
rect 14030 29362 14082 29374
rect 14254 29426 14306 29438
rect 14254 29362 14306 29374
rect 14590 29426 14642 29438
rect 14590 29362 14642 29374
rect 19406 29426 19458 29438
rect 23998 29426 24050 29438
rect 20626 29374 20638 29426
rect 20690 29374 20702 29426
rect 19406 29362 19458 29374
rect 23998 29362 24050 29374
rect 27134 29426 27186 29438
rect 27134 29362 27186 29374
rect 27358 29426 27410 29438
rect 27358 29362 27410 29374
rect 27918 29426 27970 29438
rect 27918 29362 27970 29374
rect 28478 29426 28530 29438
rect 28478 29362 28530 29374
rect 30942 29426 30994 29438
rect 30942 29362 30994 29374
rect 31614 29426 31666 29438
rect 31614 29362 31666 29374
rect 36766 29426 36818 29438
rect 36766 29362 36818 29374
rect 37438 29426 37490 29438
rect 37438 29362 37490 29374
rect 30606 29314 30658 29326
rect 2594 29262 2606 29314
rect 2658 29262 2670 29314
rect 4722 29262 4734 29314
rect 4786 29262 4798 29314
rect 21298 29262 21310 29314
rect 21362 29262 21374 29314
rect 23426 29262 23438 29314
rect 23490 29262 23502 29314
rect 37650 29262 37662 29314
rect 37714 29262 37726 29314
rect 30606 29250 30658 29262
rect 11678 29202 11730 29214
rect 11678 29138 11730 29150
rect 13918 29202 13970 29214
rect 27682 29150 27694 29202
rect 27746 29150 27758 29202
rect 13918 29138 13970 29150
rect 1344 29034 39984 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 39984 29034
rect 1344 28948 39984 28982
rect 10446 28866 10498 28878
rect 10446 28802 10498 28814
rect 11006 28866 11058 28878
rect 11006 28802 11058 28814
rect 11790 28866 11842 28878
rect 11790 28802 11842 28814
rect 29822 28866 29874 28878
rect 29822 28802 29874 28814
rect 32510 28866 32562 28878
rect 32510 28802 32562 28814
rect 8542 28754 8594 28766
rect 8542 28690 8594 28702
rect 9438 28754 9490 28766
rect 9438 28690 9490 28702
rect 10670 28754 10722 28766
rect 10670 28690 10722 28702
rect 11566 28754 11618 28766
rect 11566 28690 11618 28702
rect 13694 28754 13746 28766
rect 31166 28754 31218 28766
rect 22754 28702 22766 28754
rect 22818 28702 22830 28754
rect 13694 28690 13746 28702
rect 31166 28690 31218 28702
rect 33406 28754 33458 28766
rect 33406 28690 33458 28702
rect 7982 28642 8034 28654
rect 7982 28578 8034 28590
rect 8430 28642 8482 28654
rect 8430 28578 8482 28590
rect 8654 28642 8706 28654
rect 10894 28642 10946 28654
rect 9202 28590 9214 28642
rect 9266 28590 9278 28642
rect 9538 28590 9550 28642
rect 9602 28590 9614 28642
rect 10210 28590 10222 28642
rect 10274 28590 10286 28642
rect 8654 28578 8706 28590
rect 10894 28578 10946 28590
rect 12014 28642 12066 28654
rect 12014 28578 12066 28590
rect 12126 28642 12178 28654
rect 12126 28578 12178 28590
rect 13470 28642 13522 28654
rect 13470 28578 13522 28590
rect 13918 28642 13970 28654
rect 13918 28578 13970 28590
rect 14030 28642 14082 28654
rect 14814 28642 14866 28654
rect 14354 28590 14366 28642
rect 14418 28590 14430 28642
rect 14030 28578 14082 28590
rect 14814 28578 14866 28590
rect 20190 28642 20242 28654
rect 20190 28578 20242 28590
rect 20750 28642 20802 28654
rect 20750 28578 20802 28590
rect 27470 28642 27522 28654
rect 28130 28590 28142 28642
rect 28194 28590 28206 28642
rect 28354 28590 28366 28642
rect 28418 28590 28430 28642
rect 31378 28590 31390 28642
rect 31442 28590 31454 28642
rect 31602 28590 31614 28642
rect 31666 28590 31678 28642
rect 32834 28590 32846 28642
rect 32898 28590 32910 28642
rect 27470 28578 27522 28590
rect 8990 28530 9042 28542
rect 8990 28466 9042 28478
rect 12350 28530 12402 28542
rect 27134 28530 27186 28542
rect 20402 28478 20414 28530
rect 20466 28478 20478 28530
rect 23762 28478 23774 28530
rect 23826 28478 23838 28530
rect 12350 28466 12402 28478
rect 27134 28466 27186 28478
rect 28702 28530 28754 28542
rect 28702 28466 28754 28478
rect 29710 28530 29762 28542
rect 29710 28466 29762 28478
rect 30830 28530 30882 28542
rect 30830 28466 30882 28478
rect 9774 28418 9826 28430
rect 26798 28418 26850 28430
rect 14018 28366 14030 28418
rect 14082 28366 14094 28418
rect 9774 28354 9826 28366
rect 26798 28354 26850 28366
rect 26910 28418 26962 28430
rect 26910 28354 26962 28366
rect 28590 28418 28642 28430
rect 28590 28354 28642 28366
rect 29822 28418 29874 28430
rect 29822 28354 29874 28366
rect 30494 28418 30546 28430
rect 30494 28354 30546 28366
rect 32622 28418 32674 28430
rect 32622 28354 32674 28366
rect 1344 28250 39984 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 39984 28250
rect 1344 28164 39984 28198
rect 8990 28082 9042 28094
rect 8990 28018 9042 28030
rect 11230 28082 11282 28094
rect 11230 28018 11282 28030
rect 15374 28082 15426 28094
rect 15374 28018 15426 28030
rect 21758 28082 21810 28094
rect 21758 28018 21810 28030
rect 22654 28082 22706 28094
rect 22654 28018 22706 28030
rect 8542 27970 8594 27982
rect 8542 27906 8594 27918
rect 10334 27970 10386 27982
rect 10334 27906 10386 27918
rect 21646 27970 21698 27982
rect 21646 27906 21698 27918
rect 21982 27970 22034 27982
rect 21982 27906 22034 27918
rect 23102 27970 23154 27982
rect 37214 27970 37266 27982
rect 33618 27918 33630 27970
rect 33682 27918 33694 27970
rect 23102 27906 23154 27918
rect 37214 27906 37266 27918
rect 8430 27858 8482 27870
rect 3826 27806 3838 27858
rect 3890 27806 3902 27858
rect 7858 27806 7870 27858
rect 7922 27806 7934 27858
rect 8430 27794 8482 27806
rect 10446 27858 10498 27870
rect 10446 27794 10498 27806
rect 10894 27858 10946 27870
rect 10894 27794 10946 27806
rect 22206 27858 22258 27870
rect 22206 27794 22258 27806
rect 26910 27858 26962 27870
rect 28242 27806 28254 27858
rect 28306 27806 28318 27858
rect 33394 27806 33406 27858
rect 33458 27806 33470 27858
rect 37650 27806 37662 27858
rect 37714 27806 37726 27858
rect 26910 27794 26962 27806
rect 6750 27746 6802 27758
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 6750 27682 6802 27694
rect 26238 27746 26290 27758
rect 35534 27746 35586 27758
rect 31826 27694 31838 27746
rect 31890 27694 31902 27746
rect 38098 27694 38110 27746
rect 38162 27694 38174 27746
rect 26238 27682 26290 27694
rect 35534 27682 35586 27694
rect 11118 27634 11170 27646
rect 15026 27582 15038 27634
rect 15090 27631 15102 27634
rect 15362 27631 15374 27634
rect 15090 27585 15374 27631
rect 15090 27582 15102 27585
rect 15362 27582 15374 27585
rect 15426 27582 15438 27634
rect 22306 27582 22318 27634
rect 22370 27631 22382 27634
rect 22866 27631 22878 27634
rect 22370 27585 22878 27631
rect 22370 27582 22382 27585
rect 22866 27582 22878 27585
rect 22930 27582 22942 27634
rect 11118 27570 11170 27582
rect 1344 27466 39984 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 39984 27466
rect 1344 27380 39984 27414
rect 8878 27186 8930 27198
rect 10446 27186 10498 27198
rect 4610 27134 4622 27186
rect 4674 27134 4686 27186
rect 9762 27134 9774 27186
rect 9826 27134 9838 27186
rect 8878 27122 8930 27134
rect 10446 27122 10498 27134
rect 11118 27186 11170 27198
rect 30158 27186 30210 27198
rect 35198 27186 35250 27198
rect 11890 27134 11902 27186
rect 11954 27134 11966 27186
rect 18834 27134 18846 27186
rect 18898 27134 18910 27186
rect 25890 27134 25902 27186
rect 25954 27134 25966 27186
rect 26674 27134 26686 27186
rect 26738 27134 26750 27186
rect 29362 27134 29374 27186
rect 29426 27134 29438 27186
rect 31826 27134 31838 27186
rect 31890 27134 31902 27186
rect 33954 27134 33966 27186
rect 34018 27134 34030 27186
rect 37314 27134 37326 27186
rect 37378 27134 37390 27186
rect 11118 27122 11170 27134
rect 30158 27122 30210 27134
rect 35198 27122 35250 27134
rect 13470 27074 13522 27086
rect 35870 27074 35922 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 9314 27022 9326 27074
rect 9378 27022 9390 27074
rect 11554 27022 11566 27074
rect 11618 27022 11630 27074
rect 15026 27022 15038 27074
rect 15090 27022 15102 27074
rect 16034 27022 16046 27074
rect 16098 27022 16110 27074
rect 25218 27022 25230 27074
rect 25282 27022 25294 27074
rect 26786 27022 26798 27074
rect 26850 27022 26862 27074
rect 29474 27022 29486 27074
rect 29538 27022 29550 27074
rect 34738 27022 34750 27074
rect 34802 27022 34814 27074
rect 13470 27010 13522 27022
rect 35870 27010 35922 27022
rect 35982 27074 36034 27086
rect 35982 27010 36034 27022
rect 36094 27074 36146 27086
rect 38334 27074 38386 27086
rect 37426 27022 37438 27074
rect 37490 27022 37502 27074
rect 39218 27022 39230 27074
rect 39282 27022 39294 27074
rect 36094 27010 36146 27022
rect 38334 27010 38386 27022
rect 5070 26962 5122 26974
rect 2482 26910 2494 26962
rect 2546 26910 2558 26962
rect 5070 26898 5122 26910
rect 7198 26962 7250 26974
rect 26126 26962 26178 26974
rect 13794 26910 13806 26962
rect 13858 26910 13870 26962
rect 14802 26910 14814 26962
rect 14866 26910 14878 26962
rect 16706 26910 16718 26962
rect 16770 26910 16782 26962
rect 7198 26898 7250 26910
rect 26126 26898 26178 26910
rect 27470 26962 27522 26974
rect 27470 26898 27522 26910
rect 31502 26962 31554 26974
rect 31502 26898 31554 26910
rect 36206 26962 36258 26974
rect 36206 26898 36258 26910
rect 36430 26962 36482 26974
rect 36430 26898 36482 26910
rect 36990 26962 37042 26974
rect 36990 26898 37042 26910
rect 38558 26962 38610 26974
rect 38994 26910 39006 26962
rect 39058 26910 39070 26962
rect 38558 26898 38610 26910
rect 15598 26850 15650 26862
rect 15598 26786 15650 26798
rect 38446 26850 38498 26862
rect 38446 26786 38498 26798
rect 1344 26682 39984 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 39984 26682
rect 1344 26596 39984 26630
rect 27246 26514 27298 26526
rect 27246 26450 27298 26462
rect 27470 26514 27522 26526
rect 27470 26450 27522 26462
rect 27918 26514 27970 26526
rect 27918 26450 27970 26462
rect 34638 26514 34690 26526
rect 34638 26450 34690 26462
rect 34974 26514 35026 26526
rect 35870 26514 35922 26526
rect 35298 26462 35310 26514
rect 35362 26462 35374 26514
rect 34974 26450 35026 26462
rect 35870 26450 35922 26462
rect 27806 26402 27858 26414
rect 6626 26350 6638 26402
rect 6690 26350 6702 26402
rect 37426 26350 37438 26402
rect 37490 26350 37502 26402
rect 27806 26338 27858 26350
rect 28142 26290 28194 26302
rect 6402 26238 6414 26290
rect 6466 26238 6478 26290
rect 13010 26238 13022 26290
rect 13074 26238 13086 26290
rect 20066 26238 20078 26290
rect 20130 26238 20142 26290
rect 25442 26238 25454 26290
rect 25506 26238 25518 26290
rect 26786 26238 26798 26290
rect 26850 26238 26862 26290
rect 27010 26238 27022 26290
rect 27074 26238 27086 26290
rect 28142 26226 28194 26238
rect 28926 26290 28978 26302
rect 28926 26226 28978 26238
rect 30718 26290 30770 26302
rect 36206 26290 36258 26302
rect 31154 26238 31166 26290
rect 31218 26238 31230 26290
rect 30718 26226 30770 26238
rect 36206 26226 36258 26238
rect 36318 26290 36370 26302
rect 36754 26238 36766 26290
rect 36818 26238 36830 26290
rect 36318 26226 36370 26238
rect 17502 26178 17554 26190
rect 23326 26178 23378 26190
rect 29150 26178 29202 26190
rect 16258 26126 16270 26178
rect 16322 26126 16334 26178
rect 20738 26126 20750 26178
rect 20802 26126 20814 26178
rect 22866 26126 22878 26178
rect 22930 26126 22942 26178
rect 25778 26126 25790 26178
rect 25842 26126 25854 26178
rect 27234 26126 27246 26178
rect 27298 26126 27310 26178
rect 17502 26114 17554 26126
rect 23326 26114 23378 26126
rect 29150 26114 29202 26126
rect 29710 26178 29762 26190
rect 31378 26126 31390 26178
rect 31442 26126 31454 26178
rect 39554 26126 39566 26178
rect 39618 26126 39630 26178
rect 29710 26114 29762 26126
rect 28254 26066 28306 26078
rect 26114 26014 26126 26066
rect 26178 26014 26190 26066
rect 28254 26002 28306 26014
rect 28702 26066 28754 26078
rect 28702 26002 28754 26014
rect 1344 25898 39984 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 39984 25898
rect 1344 25812 39984 25846
rect 3166 25730 3218 25742
rect 3166 25666 3218 25678
rect 26238 25618 26290 25630
rect 13458 25566 13470 25618
rect 13522 25566 13534 25618
rect 15586 25566 15598 25618
rect 15650 25566 15662 25618
rect 20738 25566 20750 25618
rect 20802 25566 20814 25618
rect 30146 25566 30158 25618
rect 30210 25566 30222 25618
rect 26238 25554 26290 25566
rect 26126 25506 26178 25518
rect 7298 25454 7310 25506
rect 7362 25454 7374 25506
rect 16258 25454 16270 25506
rect 16322 25454 16334 25506
rect 17938 25454 17950 25506
rect 18002 25454 18014 25506
rect 25778 25454 25790 25506
rect 25842 25454 25854 25506
rect 27234 25454 27246 25506
rect 27298 25454 27310 25506
rect 27682 25454 27694 25506
rect 27746 25454 27758 25506
rect 30034 25454 30046 25506
rect 30098 25454 30110 25506
rect 26126 25442 26178 25454
rect 3502 25394 3554 25406
rect 29374 25394 29426 25406
rect 7522 25342 7534 25394
rect 7586 25342 7598 25394
rect 7970 25342 7982 25394
rect 8034 25342 8046 25394
rect 18610 25342 18622 25394
rect 18674 25342 18686 25394
rect 26674 25342 26686 25394
rect 26738 25342 26750 25394
rect 28354 25342 28366 25394
rect 28418 25342 28430 25394
rect 3502 25330 3554 25342
rect 29374 25330 29426 25342
rect 3278 25282 3330 25294
rect 16830 25282 16882 25294
rect 8194 25230 8206 25282
rect 8258 25230 8270 25282
rect 3278 25218 3330 25230
rect 16830 25218 16882 25230
rect 17502 25282 17554 25294
rect 17502 25218 17554 25230
rect 22766 25282 22818 25294
rect 27234 25230 27246 25282
rect 27298 25230 27310 25282
rect 22766 25218 22818 25230
rect 1344 25114 39984 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 39984 25114
rect 1344 25028 39984 25062
rect 2382 24946 2434 24958
rect 22082 24894 22094 24946
rect 22146 24894 22158 24946
rect 2382 24882 2434 24894
rect 2270 24834 2322 24846
rect 2270 24770 2322 24782
rect 4286 24834 4338 24846
rect 6862 24834 6914 24846
rect 5954 24782 5966 24834
rect 6018 24782 6030 24834
rect 6514 24782 6526 24834
rect 6578 24782 6590 24834
rect 4286 24770 4338 24782
rect 6862 24770 6914 24782
rect 27806 24834 27858 24846
rect 27806 24770 27858 24782
rect 27918 24834 27970 24846
rect 27918 24770 27970 24782
rect 28142 24834 28194 24846
rect 28142 24770 28194 24782
rect 28366 24834 28418 24846
rect 28366 24770 28418 24782
rect 28926 24834 28978 24846
rect 28926 24770 28978 24782
rect 29374 24834 29426 24846
rect 29374 24770 29426 24782
rect 2494 24722 2546 24734
rect 2494 24658 2546 24670
rect 2830 24722 2882 24734
rect 4398 24722 4450 24734
rect 18286 24722 18338 24734
rect 3490 24670 3502 24722
rect 3554 24670 3566 24722
rect 4946 24670 4958 24722
rect 5010 24670 5022 24722
rect 5730 24670 5742 24722
rect 5794 24670 5806 24722
rect 2830 24658 2882 24670
rect 4398 24658 4450 24670
rect 18286 24658 18338 24670
rect 18846 24722 18898 24734
rect 18846 24658 18898 24670
rect 19294 24722 19346 24734
rect 19294 24658 19346 24670
rect 22430 24722 22482 24734
rect 24670 24722 24722 24734
rect 26238 24722 26290 24734
rect 22866 24670 22878 24722
rect 22930 24670 22942 24722
rect 25554 24670 25566 24722
rect 25618 24670 25630 24722
rect 22430 24658 22482 24670
rect 24670 24658 24722 24670
rect 26238 24658 26290 24670
rect 27358 24722 27410 24734
rect 28590 24722 28642 24734
rect 29710 24722 29762 24734
rect 37102 24722 37154 24734
rect 27570 24670 27582 24722
rect 27634 24670 27646 24722
rect 29138 24670 29150 24722
rect 29202 24670 29214 24722
rect 30034 24670 30046 24722
rect 30098 24670 30110 24722
rect 36082 24670 36094 24722
rect 36146 24670 36158 24722
rect 27358 24658 27410 24670
rect 28590 24658 28642 24670
rect 29710 24658 29762 24670
rect 37102 24658 37154 24670
rect 23326 24610 23378 24622
rect 29038 24610 29090 24622
rect 3602 24558 3614 24610
rect 3666 24558 3678 24610
rect 25778 24558 25790 24610
rect 25842 24558 25854 24610
rect 23326 24546 23378 24558
rect 29038 24546 29090 24558
rect 29822 24610 29874 24622
rect 36766 24610 36818 24622
rect 35858 24558 35870 24610
rect 35922 24558 35934 24610
rect 29822 24546 29874 24558
rect 36766 24546 36818 24558
rect 37662 24610 37714 24622
rect 37662 24546 37714 24558
rect 27022 24498 27074 24510
rect 27022 24434 27074 24446
rect 27134 24498 27186 24510
rect 27134 24434 27186 24446
rect 1344 24330 39984 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 39984 24330
rect 1344 24244 39984 24278
rect 15250 24110 15262 24162
rect 15314 24159 15326 24162
rect 15698 24159 15710 24162
rect 15314 24113 15710 24159
rect 15314 24110 15326 24113
rect 15698 24110 15710 24113
rect 15762 24110 15774 24162
rect 12798 24050 12850 24062
rect 5618 23998 5630 24050
rect 5682 23998 5694 24050
rect 11330 23998 11342 24050
rect 11394 23998 11406 24050
rect 12798 23986 12850 23998
rect 15262 24050 15314 24062
rect 15262 23986 15314 23998
rect 15710 24050 15762 24062
rect 35982 24050 36034 24062
rect 18946 23998 18958 24050
rect 19010 23998 19022 24050
rect 24546 23998 24558 24050
rect 24610 23998 24622 24050
rect 35186 23998 35198 24050
rect 35250 23998 35262 24050
rect 15710 23986 15762 23998
rect 35982 23986 36034 23998
rect 36430 24050 36482 24062
rect 37538 23998 37550 24050
rect 37602 23998 37614 24050
rect 36430 23986 36482 23998
rect 3726 23938 3778 23950
rect 3726 23874 3778 23886
rect 4062 23938 4114 23950
rect 4062 23874 4114 23886
rect 4398 23938 4450 23950
rect 4398 23874 4450 23886
rect 4622 23938 4674 23950
rect 11902 23938 11954 23950
rect 25006 23938 25058 23950
rect 4834 23886 4846 23938
rect 4898 23886 4910 23938
rect 8418 23886 8430 23938
rect 8482 23886 8494 23938
rect 16034 23886 16046 23938
rect 16098 23886 16110 23938
rect 21746 23886 21758 23938
rect 21810 23886 21822 23938
rect 4622 23874 4674 23886
rect 11902 23874 11954 23886
rect 25006 23874 25058 23886
rect 26574 23938 26626 23950
rect 26574 23874 26626 23886
rect 31950 23938 32002 23950
rect 37102 23938 37154 23950
rect 32274 23886 32286 23938
rect 32338 23886 32350 23938
rect 31950 23874 32002 23886
rect 37102 23874 37154 23886
rect 37438 23938 37490 23950
rect 37438 23874 37490 23886
rect 5966 23826 6018 23838
rect 5966 23762 6018 23774
rect 7646 23826 7698 23838
rect 7646 23762 7698 23774
rect 7870 23826 7922 23838
rect 13694 23826 13746 23838
rect 26686 23826 26738 23838
rect 9090 23774 9102 23826
rect 9154 23774 9166 23826
rect 16818 23774 16830 23826
rect 16882 23774 16894 23826
rect 22418 23774 22430 23826
rect 22482 23774 22494 23826
rect 7870 23762 7922 23774
rect 13694 23762 13746 23774
rect 26686 23762 26738 23774
rect 26910 23826 26962 23838
rect 37550 23826 37602 23838
rect 33058 23774 33070 23826
rect 33122 23774 33134 23826
rect 26910 23762 26962 23774
rect 37550 23762 37602 23774
rect 3838 23714 3890 23726
rect 3838 23650 3890 23662
rect 4734 23714 4786 23726
rect 4734 23650 4786 23662
rect 5742 23714 5794 23726
rect 5742 23650 5794 23662
rect 7758 23714 7810 23726
rect 7758 23650 7810 23662
rect 12910 23714 12962 23726
rect 12910 23650 12962 23662
rect 13918 23714 13970 23726
rect 13918 23650 13970 23662
rect 14030 23714 14082 23726
rect 14030 23650 14082 23662
rect 14142 23714 14194 23726
rect 14142 23650 14194 23662
rect 19518 23714 19570 23726
rect 19518 23650 19570 23662
rect 31390 23714 31442 23726
rect 31390 23650 31442 23662
rect 37214 23714 37266 23726
rect 37214 23650 37266 23662
rect 1344 23546 39984 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 39984 23546
rect 1344 23460 39984 23494
rect 16270 23378 16322 23390
rect 4722 23326 4734 23378
rect 4786 23326 4798 23378
rect 16270 23314 16322 23326
rect 17502 23378 17554 23390
rect 17502 23314 17554 23326
rect 18622 23378 18674 23390
rect 18622 23314 18674 23326
rect 19518 23378 19570 23390
rect 19518 23314 19570 23326
rect 22878 23378 22930 23390
rect 22878 23314 22930 23326
rect 27582 23378 27634 23390
rect 27582 23314 27634 23326
rect 31502 23378 31554 23390
rect 31502 23314 31554 23326
rect 6862 23266 6914 23278
rect 3154 23214 3166 23266
rect 3218 23214 3230 23266
rect 6862 23202 6914 23214
rect 8430 23266 8482 23278
rect 8430 23202 8482 23214
rect 16158 23266 16210 23278
rect 16158 23202 16210 23214
rect 19070 23266 19122 23278
rect 19070 23202 19122 23214
rect 22542 23266 22594 23278
rect 22542 23202 22594 23214
rect 26910 23266 26962 23278
rect 26910 23202 26962 23214
rect 31278 23266 31330 23278
rect 35410 23214 35422 23266
rect 35474 23214 35486 23266
rect 37090 23214 37102 23266
rect 37154 23214 37166 23266
rect 31278 23202 31330 23214
rect 3502 23154 3554 23166
rect 3502 23090 3554 23102
rect 5294 23154 5346 23166
rect 5294 23090 5346 23102
rect 7198 23154 7250 23166
rect 7198 23090 7250 23102
rect 7982 23154 8034 23166
rect 15598 23154 15650 23166
rect 17390 23154 17442 23166
rect 15250 23102 15262 23154
rect 15314 23102 15326 23154
rect 15922 23102 15934 23154
rect 15986 23102 15998 23154
rect 7982 23090 8034 23102
rect 15598 23090 15650 23102
rect 17390 23090 17442 23102
rect 17726 23154 17778 23166
rect 18510 23154 18562 23166
rect 18162 23102 18174 23154
rect 18226 23102 18238 23154
rect 17726 23090 17778 23102
rect 18510 23090 18562 23102
rect 18846 23154 18898 23166
rect 18846 23090 18898 23102
rect 19406 23154 19458 23166
rect 19406 23090 19458 23102
rect 19630 23154 19682 23166
rect 22766 23154 22818 23166
rect 19954 23102 19966 23154
rect 20018 23102 20030 23154
rect 19630 23090 19682 23102
rect 22766 23090 22818 23102
rect 22990 23154 23042 23166
rect 22990 23090 23042 23102
rect 27246 23154 27298 23166
rect 31166 23154 31218 23166
rect 27682 23102 27694 23154
rect 27746 23102 27758 23154
rect 28578 23102 28590 23154
rect 28642 23102 28654 23154
rect 27246 23090 27298 23102
rect 31166 23090 31218 23102
rect 31614 23154 31666 23166
rect 31614 23090 31666 23102
rect 32062 23154 32114 23166
rect 32062 23090 32114 23102
rect 32286 23154 32338 23166
rect 38894 23154 38946 23166
rect 37314 23102 37326 23154
rect 37378 23102 37390 23154
rect 38210 23102 38222 23154
rect 38274 23102 38286 23154
rect 38546 23102 38558 23154
rect 38610 23102 38622 23154
rect 32286 23090 32338 23102
rect 38894 23090 38946 23102
rect 16830 23042 16882 23054
rect 12450 22990 12462 23042
rect 12514 22990 12526 23042
rect 14578 22990 14590 23042
rect 14642 22990 14654 23042
rect 16830 22978 16882 22990
rect 20414 23042 20466 23054
rect 20414 22978 20466 22990
rect 22094 23042 22146 23054
rect 22094 22978 22146 22990
rect 23438 23042 23490 23054
rect 23438 22978 23490 22990
rect 23886 23042 23938 23054
rect 30382 23042 30434 23054
rect 28466 22990 28478 23042
rect 28530 22990 28542 23042
rect 23886 22978 23938 22990
rect 30382 22978 30434 22990
rect 30830 23042 30882 23054
rect 30830 22978 30882 22990
rect 31838 23042 31890 23054
rect 39118 23042 39170 23054
rect 34066 22990 34078 23042
rect 34130 22990 34142 23042
rect 37426 22990 37438 23042
rect 37490 22990 37502 23042
rect 31838 22978 31890 22990
rect 39118 22978 39170 22990
rect 5070 22930 5122 22942
rect 5070 22866 5122 22878
rect 8094 22930 8146 22942
rect 8094 22866 8146 22878
rect 8318 22930 8370 22942
rect 27470 22930 27522 22942
rect 17938 22878 17950 22930
rect 18002 22878 18014 22930
rect 8318 22866 8370 22878
rect 27470 22866 27522 22878
rect 28254 22930 28306 22942
rect 28254 22866 28306 22878
rect 1344 22762 39984 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 39984 22762
rect 1344 22676 39984 22710
rect 7646 22594 7698 22606
rect 7646 22530 7698 22542
rect 14030 22594 14082 22606
rect 14030 22530 14082 22542
rect 30494 22594 30546 22606
rect 30494 22530 30546 22542
rect 8206 22482 8258 22494
rect 8206 22418 8258 22430
rect 14478 22482 14530 22494
rect 14478 22418 14530 22430
rect 16942 22482 16994 22494
rect 16942 22418 16994 22430
rect 27694 22482 27746 22494
rect 27694 22418 27746 22430
rect 30270 22482 30322 22494
rect 36990 22482 37042 22494
rect 35746 22430 35758 22482
rect 35810 22430 35822 22482
rect 37314 22430 37326 22482
rect 37378 22430 37390 22482
rect 30270 22418 30322 22430
rect 36990 22418 37042 22430
rect 5854 22370 5906 22382
rect 5854 22306 5906 22318
rect 6302 22370 6354 22382
rect 6302 22306 6354 22318
rect 6750 22370 6802 22382
rect 6750 22306 6802 22318
rect 6974 22370 7026 22382
rect 6974 22306 7026 22318
rect 7422 22370 7474 22382
rect 7422 22306 7474 22318
rect 7982 22370 8034 22382
rect 7982 22306 8034 22318
rect 9886 22370 9938 22382
rect 15150 22370 15202 22382
rect 10322 22318 10334 22370
rect 10386 22318 10398 22370
rect 13458 22318 13470 22370
rect 13522 22318 13534 22370
rect 13682 22318 13694 22370
rect 13746 22318 13758 22370
rect 14242 22318 14254 22370
rect 14306 22318 14318 22370
rect 9886 22306 9938 22318
rect 15150 22306 15202 22318
rect 15710 22370 15762 22382
rect 15710 22306 15762 22318
rect 16046 22370 16098 22382
rect 16046 22306 16098 22318
rect 17950 22370 18002 22382
rect 17950 22306 18002 22318
rect 18286 22370 18338 22382
rect 29262 22370 29314 22382
rect 18946 22318 18958 22370
rect 19010 22318 19022 22370
rect 20066 22318 20078 22370
rect 20130 22318 20142 22370
rect 18286 22306 18338 22318
rect 29262 22306 29314 22318
rect 29934 22370 29986 22382
rect 29934 22306 29986 22318
rect 30046 22370 30098 22382
rect 30046 22306 30098 22318
rect 32174 22370 32226 22382
rect 36430 22370 36482 22382
rect 32834 22318 32846 22370
rect 32898 22318 32910 22370
rect 37426 22318 37438 22370
rect 37490 22318 37502 22370
rect 32174 22306 32226 22318
rect 36430 22306 36482 22318
rect 5966 22258 6018 22270
rect 9998 22258 10050 22270
rect 8866 22206 8878 22258
rect 8930 22206 8942 22258
rect 5966 22194 6018 22206
rect 9998 22194 10050 22206
rect 10110 22258 10162 22270
rect 10110 22194 10162 22206
rect 10782 22258 10834 22270
rect 10782 22194 10834 22206
rect 14590 22258 14642 22270
rect 14590 22194 14642 22206
rect 15486 22258 15538 22270
rect 15486 22194 15538 22206
rect 15598 22258 15650 22270
rect 19854 22258 19906 22270
rect 29374 22258 29426 22270
rect 19058 22206 19070 22258
rect 19122 22206 19134 22258
rect 20402 22206 20414 22258
rect 20466 22206 20478 22258
rect 15598 22194 15650 22206
rect 19854 22194 19906 22206
rect 29374 22194 29426 22206
rect 31950 22258 32002 22270
rect 31950 22194 32002 22206
rect 32510 22258 32562 22270
rect 33618 22206 33630 22258
rect 33682 22206 33694 22258
rect 36082 22206 36094 22258
rect 36146 22206 36158 22258
rect 32510 22194 32562 22206
rect 6190 22146 6242 22158
rect 6190 22082 6242 22094
rect 6862 22146 6914 22158
rect 6862 22082 6914 22094
rect 7310 22146 7362 22158
rect 7310 22082 7362 22094
rect 8542 22146 8594 22158
rect 8542 22082 8594 22094
rect 13918 22146 13970 22158
rect 13918 22082 13970 22094
rect 16606 22146 16658 22158
rect 16606 22082 16658 22094
rect 17838 22146 17890 22158
rect 17838 22082 17890 22094
rect 18174 22146 18226 22158
rect 20750 22146 20802 22158
rect 18946 22094 18958 22146
rect 19010 22094 19022 22146
rect 18174 22082 18226 22094
rect 20750 22082 20802 22094
rect 28254 22146 28306 22158
rect 28254 22082 28306 22094
rect 29822 22146 29874 22158
rect 29822 22082 29874 22094
rect 30942 22146 30994 22158
rect 30942 22082 30994 22094
rect 31502 22146 31554 22158
rect 31502 22082 31554 22094
rect 31726 22146 31778 22158
rect 31726 22082 31778 22094
rect 31838 22146 31890 22158
rect 31838 22082 31890 22094
rect 32398 22146 32450 22158
rect 32398 22082 32450 22094
rect 1344 21978 39984 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 39984 21978
rect 1344 21892 39984 21926
rect 8430 21810 8482 21822
rect 8430 21746 8482 21758
rect 14702 21810 14754 21822
rect 14702 21746 14754 21758
rect 18734 21810 18786 21822
rect 18734 21746 18786 21758
rect 25342 21810 25394 21822
rect 25342 21746 25394 21758
rect 32622 21810 32674 21822
rect 32622 21746 32674 21758
rect 8654 21698 8706 21710
rect 7746 21646 7758 21698
rect 7810 21646 7822 21698
rect 8654 21634 8706 21646
rect 9550 21698 9602 21710
rect 9550 21634 9602 21646
rect 9774 21698 9826 21710
rect 31838 21698 31890 21710
rect 14354 21646 14366 21698
rect 14418 21646 14430 21698
rect 26674 21646 26686 21698
rect 26738 21646 26750 21698
rect 27794 21646 27806 21698
rect 27858 21646 27870 21698
rect 33170 21646 33182 21698
rect 33234 21646 33246 21698
rect 9774 21634 9826 21646
rect 31838 21634 31890 21646
rect 8206 21586 8258 21598
rect 3714 21534 3726 21586
rect 3778 21534 3790 21586
rect 5058 21534 5070 21586
rect 5122 21534 5134 21586
rect 6402 21534 6414 21586
rect 6466 21534 6478 21586
rect 6962 21534 6974 21586
rect 7026 21534 7038 21586
rect 7522 21534 7534 21586
rect 7586 21534 7598 21586
rect 8206 21522 8258 21534
rect 8878 21586 8930 21598
rect 14590 21586 14642 21598
rect 18510 21586 18562 21598
rect 13458 21534 13470 21586
rect 13522 21534 13534 21586
rect 13794 21534 13806 21586
rect 13858 21534 13870 21586
rect 14914 21534 14926 21586
rect 14978 21534 14990 21586
rect 15138 21534 15150 21586
rect 15202 21534 15214 21586
rect 8878 21522 8930 21534
rect 14590 21522 14642 21534
rect 18510 21522 18562 21534
rect 18846 21586 18898 21598
rect 18846 21522 18898 21534
rect 19070 21586 19122 21598
rect 25902 21586 25954 21598
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 19070 21522 19122 21534
rect 25902 21522 25954 21534
rect 26350 21586 26402 21598
rect 27010 21534 27022 21586
rect 27074 21534 27086 21586
rect 31154 21534 31166 21586
rect 31218 21534 31230 21586
rect 36642 21534 36654 21586
rect 36706 21534 36718 21586
rect 26350 21522 26402 21534
rect 3054 21474 3106 21486
rect 5406 21474 5458 21486
rect 15598 21474 15650 21486
rect 30494 21474 30546 21486
rect 36430 21474 36482 21486
rect 3938 21422 3950 21474
rect 4002 21422 4014 21474
rect 7858 21422 7870 21474
rect 7922 21422 7934 21474
rect 9874 21422 9886 21474
rect 9938 21422 9950 21474
rect 13906 21422 13918 21474
rect 13970 21422 13982 21474
rect 22978 21422 22990 21474
rect 23042 21422 23054 21474
rect 29922 21422 29934 21474
rect 29986 21422 29998 21474
rect 31378 21422 31390 21474
rect 31442 21422 31454 21474
rect 34290 21422 34302 21474
rect 34354 21422 34366 21474
rect 37426 21422 37438 21474
rect 37490 21422 37502 21474
rect 39554 21422 39566 21474
rect 39618 21422 39630 21474
rect 3054 21410 3106 21422
rect 5406 21410 5458 21422
rect 15598 21410 15650 21422
rect 30494 21410 30546 21422
rect 36430 21410 36482 21422
rect 1344 21194 39984 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 39984 21194
rect 1344 21108 39984 21142
rect 11566 21026 11618 21038
rect 19630 21026 19682 21038
rect 9538 20974 9550 21026
rect 9602 20974 9614 21026
rect 18834 20974 18846 21026
rect 18898 21023 18910 21026
rect 19394 21023 19406 21026
rect 18898 20977 19406 21023
rect 18898 20974 18910 20977
rect 19394 20974 19406 20977
rect 19458 20974 19470 21026
rect 11566 20962 11618 20974
rect 19630 20962 19682 20974
rect 19966 21026 20018 21038
rect 19966 20962 20018 20974
rect 37438 21026 37490 21038
rect 37438 20962 37490 20974
rect 7422 20914 7474 20926
rect 4610 20862 4622 20914
rect 4674 20862 4686 20914
rect 7422 20850 7474 20862
rect 7646 20914 7698 20926
rect 7646 20850 7698 20862
rect 18846 20914 18898 20926
rect 32286 20914 32338 20926
rect 25666 20862 25678 20914
rect 25730 20862 25742 20914
rect 31826 20862 31838 20914
rect 31890 20862 31902 20914
rect 18846 20850 18898 20862
rect 32286 20850 32338 20862
rect 33070 20914 33122 20926
rect 33070 20850 33122 20862
rect 37550 20914 37602 20926
rect 37550 20850 37602 20862
rect 7870 20802 7922 20814
rect 1810 20750 1822 20802
rect 1874 20750 1886 20802
rect 7870 20738 7922 20750
rect 8654 20802 8706 20814
rect 8654 20738 8706 20750
rect 10446 20802 10498 20814
rect 10446 20738 10498 20750
rect 19742 20802 19794 20814
rect 19742 20738 19794 20750
rect 20078 20802 20130 20814
rect 26350 20802 26402 20814
rect 22866 20750 22878 20802
rect 22930 20750 22942 20802
rect 20078 20738 20130 20750
rect 26350 20738 26402 20750
rect 26798 20802 26850 20814
rect 26798 20738 26850 20750
rect 27246 20802 27298 20814
rect 27246 20738 27298 20750
rect 27694 20802 27746 20814
rect 33406 20802 33458 20814
rect 31602 20750 31614 20802
rect 31666 20750 31678 20802
rect 37762 20750 37774 20802
rect 37826 20750 37838 20802
rect 27694 20738 27746 20750
rect 33406 20738 33458 20750
rect 8318 20690 8370 20702
rect 11678 20690 11730 20702
rect 21646 20690 21698 20702
rect 27582 20690 27634 20702
rect 2482 20638 2494 20690
rect 2546 20638 2558 20690
rect 9650 20638 9662 20690
rect 9714 20638 9726 20690
rect 10098 20638 10110 20690
rect 10162 20638 10174 20690
rect 15026 20638 15038 20690
rect 15090 20638 15102 20690
rect 23538 20638 23550 20690
rect 23602 20638 23614 20690
rect 26002 20638 26014 20690
rect 26066 20638 26078 20690
rect 8318 20626 8370 20638
rect 11678 20626 11730 20638
rect 21646 20626 21698 20638
rect 27582 20626 27634 20638
rect 28254 20690 28306 20702
rect 28254 20626 28306 20638
rect 5070 20578 5122 20590
rect 11230 20578 11282 20590
rect 7074 20526 7086 20578
rect 7138 20526 7150 20578
rect 5070 20514 5122 20526
rect 11230 20514 11282 20526
rect 11566 20578 11618 20590
rect 11566 20514 11618 20526
rect 14702 20578 14754 20590
rect 14702 20514 14754 20526
rect 19294 20578 19346 20590
rect 19294 20514 19346 20526
rect 21310 20578 21362 20590
rect 21310 20514 21362 20526
rect 27470 20578 27522 20590
rect 27470 20514 27522 20526
rect 30494 20578 30546 20590
rect 37102 20578 37154 20590
rect 33730 20526 33742 20578
rect 33794 20526 33806 20578
rect 30494 20514 30546 20526
rect 37102 20514 37154 20526
rect 1344 20410 39984 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 39984 20410
rect 1344 20324 39984 20358
rect 8654 20242 8706 20254
rect 5842 20190 5854 20242
rect 5906 20190 5918 20242
rect 14130 20190 14142 20242
rect 14194 20190 14206 20242
rect 8654 20178 8706 20190
rect 2942 20130 2994 20142
rect 2942 20066 2994 20078
rect 3166 20130 3218 20142
rect 3166 20066 3218 20078
rect 6414 20130 6466 20142
rect 6414 20066 6466 20078
rect 9550 20130 9602 20142
rect 12686 20130 12738 20142
rect 10770 20078 10782 20130
rect 10834 20078 10846 20130
rect 9550 20066 9602 20078
rect 12686 20066 12738 20078
rect 15150 20130 15202 20142
rect 15150 20066 15202 20078
rect 15486 20130 15538 20142
rect 15486 20066 15538 20078
rect 16382 20130 16434 20142
rect 17390 20130 17442 20142
rect 21534 20130 21586 20142
rect 16706 20078 16718 20130
rect 16770 20078 16782 20130
rect 20514 20078 20526 20130
rect 20578 20078 20590 20130
rect 16382 20066 16434 20078
rect 17390 20066 17442 20078
rect 21534 20066 21586 20078
rect 26910 20130 26962 20142
rect 26910 20066 26962 20078
rect 27022 20130 27074 20142
rect 27022 20066 27074 20078
rect 28030 20130 28082 20142
rect 35970 20078 35982 20130
rect 36034 20078 36046 20130
rect 28030 20066 28082 20078
rect 6302 20018 6354 20030
rect 6302 19954 6354 19966
rect 6526 20018 6578 20030
rect 9774 20018 9826 20030
rect 8418 19966 8430 20018
rect 8482 19966 8494 20018
rect 6526 19954 6578 19966
rect 9774 19954 9826 19966
rect 12238 20018 12290 20030
rect 12238 19954 12290 19966
rect 12798 20018 12850 20030
rect 14478 20018 14530 20030
rect 13346 19966 13358 20018
rect 13410 19966 13422 20018
rect 12798 19954 12850 19966
rect 14478 19954 14530 19966
rect 14814 20018 14866 20030
rect 19406 20018 19458 20030
rect 19966 20018 20018 20030
rect 15922 19966 15934 20018
rect 15986 19966 15998 20018
rect 18946 19966 18958 20018
rect 19010 19966 19022 20018
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 14814 19954 14866 19966
rect 19406 19954 19458 19966
rect 19966 19954 20018 19966
rect 20078 20018 20130 20030
rect 23774 20018 23826 20030
rect 22082 19966 22094 20018
rect 22146 19966 22158 20018
rect 23090 19966 23102 20018
rect 23154 19966 23166 20018
rect 20078 19954 20130 19966
rect 23774 19954 23826 19966
rect 24222 20018 24274 20030
rect 24222 19954 24274 19966
rect 24446 20018 24498 20030
rect 24446 19954 24498 19966
rect 25902 20018 25954 20030
rect 25902 19954 25954 19966
rect 26126 20018 26178 20030
rect 26126 19954 26178 19966
rect 26350 20018 26402 20030
rect 28590 20018 28642 20030
rect 26674 19966 26686 20018
rect 26738 19966 26750 20018
rect 35746 19966 35758 20018
rect 35810 19966 35822 20018
rect 26350 19954 26402 19966
rect 28590 19954 28642 19966
rect 4286 19906 4338 19918
rect 2818 19854 2830 19906
rect 2882 19854 2894 19906
rect 4286 19842 4338 19854
rect 12462 19906 12514 19918
rect 12462 19842 12514 19854
rect 13806 19906 13858 19918
rect 21198 19906 21250 19918
rect 17826 19854 17838 19906
rect 17890 19854 17902 19906
rect 13806 19842 13858 19854
rect 21198 19842 21250 19854
rect 21646 19906 21698 19918
rect 21646 19842 21698 19854
rect 21870 19906 21922 19918
rect 23998 19906 24050 19918
rect 22642 19854 22654 19906
rect 22706 19854 22718 19906
rect 28130 19854 28142 19906
rect 28194 19854 28206 19906
rect 21870 19842 21922 19854
rect 23998 19842 24050 19854
rect 9998 19794 10050 19806
rect 9998 19730 10050 19742
rect 10222 19794 10274 19806
rect 25454 19794 25506 19806
rect 27806 19794 27858 19806
rect 23202 19742 23214 19794
rect 23266 19742 23278 19794
rect 27458 19742 27470 19794
rect 27522 19742 27534 19794
rect 10222 19730 10274 19742
rect 25454 19730 25506 19742
rect 27806 19730 27858 19742
rect 1344 19626 39984 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 39984 19626
rect 1344 19540 39984 19574
rect 3838 19458 3890 19470
rect 13694 19458 13746 19470
rect 23214 19458 23266 19470
rect 5618 19406 5630 19458
rect 5682 19406 5694 19458
rect 22082 19406 22094 19458
rect 22146 19406 22158 19458
rect 3838 19394 3890 19406
rect 13694 19394 13746 19406
rect 23214 19394 23266 19406
rect 26350 19458 26402 19470
rect 31502 19458 31554 19470
rect 31154 19406 31166 19458
rect 31218 19406 31230 19458
rect 26350 19394 26402 19406
rect 31502 19394 31554 19406
rect 33406 19458 33458 19470
rect 33406 19394 33458 19406
rect 15934 19346 15986 19358
rect 26798 19346 26850 19358
rect 14578 19294 14590 19346
rect 14642 19294 14654 19346
rect 20626 19294 20638 19346
rect 20690 19294 20702 19346
rect 23426 19294 23438 19346
rect 23490 19294 23502 19346
rect 15934 19282 15986 19294
rect 26798 19282 26850 19294
rect 37550 19346 37602 19358
rect 37550 19282 37602 19294
rect 3614 19234 3666 19246
rect 5070 19234 5122 19246
rect 4050 19182 4062 19234
rect 4114 19182 4126 19234
rect 3614 19170 3666 19182
rect 5070 19170 5122 19182
rect 5966 19234 6018 19246
rect 5966 19170 6018 19182
rect 6190 19234 6242 19246
rect 13470 19234 13522 19246
rect 9090 19182 9102 19234
rect 9154 19182 9166 19234
rect 11106 19182 11118 19234
rect 11170 19182 11182 19234
rect 6190 19170 6242 19182
rect 13470 19170 13522 19182
rect 14254 19234 14306 19246
rect 14254 19170 14306 19182
rect 17054 19234 17106 19246
rect 27022 19234 27074 19246
rect 21298 19182 21310 19234
rect 21362 19182 21374 19234
rect 23538 19182 23550 19234
rect 23602 19182 23614 19234
rect 17054 19170 17106 19182
rect 27022 19170 27074 19182
rect 27246 19234 27298 19246
rect 27246 19170 27298 19182
rect 31726 19234 31778 19246
rect 31726 19170 31778 19182
rect 32062 19234 32114 19246
rect 32062 19170 32114 19182
rect 32174 19234 32226 19246
rect 37326 19234 37378 19246
rect 32498 19182 32510 19234
rect 32562 19182 32574 19234
rect 33394 19182 33406 19234
rect 33458 19182 33470 19234
rect 32174 19170 32226 19182
rect 37326 19170 37378 19182
rect 3502 19122 3554 19134
rect 14814 19122 14866 19134
rect 4722 19070 4734 19122
rect 4786 19070 4798 19122
rect 9202 19070 9214 19122
rect 9266 19070 9278 19122
rect 12898 19070 12910 19122
rect 12962 19070 12974 19122
rect 3502 19058 3554 19070
rect 14814 19058 14866 19070
rect 19630 19122 19682 19134
rect 19630 19058 19682 19070
rect 21534 19122 21586 19134
rect 21534 19058 21586 19070
rect 21646 19122 21698 19134
rect 33742 19122 33794 19134
rect 22754 19070 22766 19122
rect 22818 19119 22830 19122
rect 23090 19119 23102 19122
rect 22818 19073 23102 19119
rect 22818 19070 22830 19073
rect 23090 19070 23102 19073
rect 23154 19070 23166 19122
rect 21646 19058 21698 19070
rect 33742 19058 33794 19070
rect 36206 19122 36258 19134
rect 36206 19058 36258 19070
rect 36318 19122 36370 19134
rect 36318 19058 36370 19070
rect 14590 19010 14642 19022
rect 12786 18958 12798 19010
rect 12850 18958 12862 19010
rect 14018 18958 14030 19010
rect 14082 18958 14094 19010
rect 14590 18946 14642 18958
rect 15150 19010 15202 19022
rect 20190 19010 20242 19022
rect 15474 18958 15486 19010
rect 15538 18958 15550 19010
rect 17378 18958 17390 19010
rect 17442 18958 17454 19010
rect 19282 18958 19294 19010
rect 19346 18958 19358 19010
rect 15150 18946 15202 18958
rect 20190 18946 20242 18958
rect 27694 19010 27746 19022
rect 27694 18946 27746 18958
rect 36542 19010 36594 19022
rect 36978 18958 36990 19010
rect 37042 18958 37054 19010
rect 36542 18946 36594 18958
rect 1344 18842 39984 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 39984 18842
rect 1344 18756 39984 18790
rect 4286 18674 4338 18686
rect 4286 18610 4338 18622
rect 14590 18674 14642 18686
rect 14590 18610 14642 18622
rect 18286 18674 18338 18686
rect 18286 18610 18338 18622
rect 19742 18674 19794 18686
rect 19742 18610 19794 18622
rect 31950 18674 32002 18686
rect 31950 18610 32002 18622
rect 33070 18674 33122 18686
rect 33070 18610 33122 18622
rect 38334 18674 38386 18686
rect 38334 18610 38386 18622
rect 19854 18562 19906 18574
rect 31726 18562 31778 18574
rect 36094 18562 36146 18574
rect 26450 18510 26462 18562
rect 26514 18510 26526 18562
rect 35746 18510 35758 18562
rect 35810 18510 35822 18562
rect 19854 18498 19906 18510
rect 31726 18498 31778 18510
rect 36094 18498 36146 18510
rect 38110 18562 38162 18574
rect 38110 18498 38162 18510
rect 18398 18450 18450 18462
rect 4498 18398 4510 18450
rect 4562 18398 4574 18450
rect 13682 18398 13694 18450
rect 13746 18398 13758 18450
rect 18398 18386 18450 18398
rect 18846 18450 18898 18462
rect 18846 18386 18898 18398
rect 26126 18450 26178 18462
rect 26126 18386 26178 18398
rect 32286 18450 32338 18462
rect 32286 18386 32338 18398
rect 33742 18450 33794 18462
rect 36318 18450 36370 18462
rect 38222 18450 38274 18462
rect 35858 18398 35870 18450
rect 35922 18398 35934 18450
rect 37090 18398 37102 18450
rect 37154 18398 37166 18450
rect 33742 18386 33794 18398
rect 36318 18386 36370 18398
rect 38222 18386 38274 18398
rect 14702 18338 14754 18350
rect 13906 18286 13918 18338
rect 13970 18286 13982 18338
rect 14702 18274 14754 18286
rect 33966 18338 34018 18350
rect 33966 18274 34018 18286
rect 34414 18338 34466 18350
rect 35970 18286 35982 18338
rect 36034 18286 36046 18338
rect 37538 18286 37550 18338
rect 37602 18286 37614 18338
rect 34414 18274 34466 18286
rect 4174 18226 4226 18238
rect 18286 18226 18338 18238
rect 14130 18174 14142 18226
rect 14194 18174 14206 18226
rect 4174 18162 4226 18174
rect 18286 18162 18338 18174
rect 19742 18226 19794 18238
rect 19742 18162 19794 18174
rect 31614 18226 31666 18238
rect 31614 18162 31666 18174
rect 33182 18226 33234 18238
rect 33182 18162 33234 18174
rect 33406 18226 33458 18238
rect 37202 18174 37214 18226
rect 37266 18174 37278 18226
rect 33406 18162 33458 18174
rect 1344 18058 39984 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 39984 18058
rect 1344 17972 39984 18006
rect 20178 17838 20190 17890
rect 20242 17838 20254 17890
rect 23426 17838 23438 17890
rect 23490 17838 23502 17890
rect 31266 17838 31278 17890
rect 31330 17887 31342 17890
rect 31602 17887 31614 17890
rect 31330 17841 31614 17887
rect 31330 17838 31342 17841
rect 31602 17838 31614 17841
rect 31666 17838 31678 17890
rect 5070 17778 5122 17790
rect 25118 17778 25170 17790
rect 2482 17726 2494 17778
rect 2546 17726 2558 17778
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 19058 17726 19070 17778
rect 19122 17726 19134 17778
rect 5070 17714 5122 17726
rect 25118 17714 25170 17726
rect 34750 17778 34802 17790
rect 34750 17714 34802 17726
rect 37102 17778 37154 17790
rect 37102 17714 37154 17726
rect 8766 17666 8818 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 5730 17614 5742 17666
rect 5794 17614 5806 17666
rect 8766 17602 8818 17614
rect 15822 17666 15874 17678
rect 19630 17666 19682 17678
rect 16146 17614 16158 17666
rect 16210 17614 16222 17666
rect 15822 17602 15874 17614
rect 19630 17602 19682 17614
rect 19742 17666 19794 17678
rect 19742 17602 19794 17614
rect 22542 17666 22594 17678
rect 23202 17614 23214 17666
rect 23266 17614 23278 17666
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 36978 17614 36990 17666
rect 37042 17614 37054 17666
rect 37202 17614 37214 17666
rect 37266 17614 37278 17666
rect 22542 17602 22594 17614
rect 5966 17554 6018 17566
rect 5966 17490 6018 17502
rect 8430 17554 8482 17566
rect 8430 17490 8482 17502
rect 8542 17554 8594 17566
rect 19518 17554 19570 17566
rect 23998 17554 24050 17566
rect 16930 17502 16942 17554
rect 16994 17502 17006 17554
rect 22866 17502 22878 17554
rect 22930 17502 22942 17554
rect 8542 17490 8594 17502
rect 19518 17490 19570 17502
rect 23998 17490 24050 17502
rect 24334 17554 24386 17566
rect 24334 17490 24386 17502
rect 24558 17554 24610 17566
rect 37438 17554 37490 17566
rect 32610 17502 32622 17554
rect 32674 17502 32686 17554
rect 24558 17490 24610 17502
rect 37438 17490 37490 17502
rect 37886 17554 37938 17566
rect 37886 17490 37938 17502
rect 37998 17554 38050 17566
rect 37998 17490 38050 17502
rect 24446 17442 24498 17454
rect 23650 17390 23662 17442
rect 23714 17390 23726 17442
rect 24446 17378 24498 17390
rect 31614 17442 31666 17454
rect 31614 17378 31666 17390
rect 37662 17442 37714 17454
rect 37662 17378 37714 17390
rect 1344 17274 39984 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 39984 17274
rect 1344 17188 39984 17222
rect 11678 17106 11730 17118
rect 11678 17042 11730 17054
rect 17614 17106 17666 17118
rect 17614 17042 17666 17054
rect 18846 17106 18898 17118
rect 18846 17042 18898 17054
rect 22878 17106 22930 17118
rect 22878 17042 22930 17054
rect 23438 17106 23490 17118
rect 23438 17042 23490 17054
rect 29934 17106 29986 17118
rect 29934 17042 29986 17054
rect 30494 17106 30546 17118
rect 30494 17042 30546 17054
rect 32062 17106 32114 17118
rect 36642 17054 36654 17106
rect 36706 17054 36718 17106
rect 32062 17042 32114 17054
rect 7310 16994 7362 17006
rect 7310 16930 7362 16942
rect 7646 16994 7698 17006
rect 7646 16930 7698 16942
rect 10558 16994 10610 17006
rect 10558 16930 10610 16942
rect 11118 16994 11170 17006
rect 11118 16930 11170 16942
rect 18398 16994 18450 17006
rect 18398 16930 18450 16942
rect 23214 16994 23266 17006
rect 23214 16930 23266 16942
rect 23550 16994 23602 17006
rect 23550 16930 23602 16942
rect 24558 16994 24610 17006
rect 30046 16994 30098 17006
rect 25218 16942 25230 16994
rect 25282 16942 25294 16994
rect 27458 16942 27470 16994
rect 27522 16942 27534 16994
rect 24558 16930 24610 16942
rect 30046 16930 30098 16942
rect 30942 16994 30994 17006
rect 31602 16942 31614 16994
rect 31666 16942 31678 16994
rect 35298 16942 35310 16994
rect 35362 16942 35374 16994
rect 30942 16930 30994 16942
rect 10446 16882 10498 16894
rect 17950 16882 18002 16894
rect 23662 16882 23714 16894
rect 25566 16882 25618 16894
rect 32174 16882 32226 16894
rect 10098 16830 10110 16882
rect 10162 16830 10174 16882
rect 17826 16830 17838 16882
rect 17890 16830 17902 16882
rect 18162 16830 18174 16882
rect 18226 16830 18238 16882
rect 24098 16830 24110 16882
rect 24162 16830 24174 16882
rect 24322 16830 24334 16882
rect 24386 16830 24398 16882
rect 26786 16830 26798 16882
rect 26850 16830 26862 16882
rect 31378 16830 31390 16882
rect 31442 16830 31454 16882
rect 10446 16818 10498 16830
rect 17950 16818 18002 16830
rect 23662 16818 23714 16830
rect 25566 16818 25618 16830
rect 32174 16818 32226 16830
rect 32958 16882 33010 16894
rect 32958 16818 33010 16830
rect 19294 16770 19346 16782
rect 37214 16770 37266 16782
rect 11218 16718 11230 16770
rect 11282 16718 11294 16770
rect 29586 16718 29598 16770
rect 29650 16718 29662 16770
rect 19294 16706 19346 16718
rect 37214 16706 37266 16718
rect 10894 16658 10946 16670
rect 10894 16594 10946 16606
rect 24222 16658 24274 16670
rect 24222 16594 24274 16606
rect 32062 16658 32114 16670
rect 32062 16594 32114 16606
rect 36990 16658 37042 16670
rect 36990 16594 37042 16606
rect 1344 16490 39984 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 39984 16490
rect 1344 16404 39984 16438
rect 6078 16322 6130 16334
rect 6078 16258 6130 16270
rect 6302 16322 6354 16334
rect 6302 16258 6354 16270
rect 7758 16322 7810 16334
rect 30046 16322 30098 16334
rect 22642 16270 22654 16322
rect 22706 16270 22718 16322
rect 7758 16258 7810 16270
rect 30046 16258 30098 16270
rect 3502 16210 3554 16222
rect 3502 16146 3554 16158
rect 9886 16210 9938 16222
rect 9886 16146 9938 16158
rect 10446 16210 10498 16222
rect 10446 16146 10498 16158
rect 12574 16210 12626 16222
rect 12574 16146 12626 16158
rect 15710 16210 15762 16222
rect 15710 16146 15762 16158
rect 18174 16210 18226 16222
rect 18174 16146 18226 16158
rect 18734 16210 18786 16222
rect 18734 16146 18786 16158
rect 19854 16210 19906 16222
rect 36990 16210 37042 16222
rect 31602 16158 31614 16210
rect 31666 16158 31678 16210
rect 33730 16158 33742 16210
rect 33794 16158 33806 16210
rect 19854 16146 19906 16158
rect 36990 16146 37042 16158
rect 5854 16098 5906 16110
rect 4274 16046 4286 16098
rect 4338 16046 4350 16098
rect 5854 16034 5906 16046
rect 6750 16098 6802 16110
rect 6750 16034 6802 16046
rect 7086 16098 7138 16110
rect 9774 16098 9826 16110
rect 9202 16046 9214 16098
rect 9266 16046 9278 16098
rect 7086 16034 7138 16046
rect 9774 16034 9826 16046
rect 23214 16098 23266 16110
rect 26686 16098 26738 16110
rect 28590 16098 28642 16110
rect 24434 16046 24446 16098
rect 24498 16046 24510 16098
rect 25554 16046 25566 16098
rect 25618 16046 25630 16098
rect 27010 16046 27022 16098
rect 27074 16046 27086 16098
rect 23214 16034 23266 16046
rect 26686 16034 26738 16046
rect 28590 16034 28642 16046
rect 30494 16098 30546 16110
rect 35534 16098 35586 16110
rect 37886 16098 37938 16110
rect 34402 16046 34414 16098
rect 34466 16046 34478 16098
rect 37426 16046 37438 16098
rect 37490 16046 37502 16098
rect 38546 16046 38558 16098
rect 38610 16046 38622 16098
rect 30494 16034 30546 16046
rect 35534 16034 35586 16046
rect 37886 16034 37938 16046
rect 3950 15986 4002 15998
rect 3950 15922 4002 15934
rect 5630 15986 5682 15998
rect 5630 15922 5682 15934
rect 7646 15986 7698 15998
rect 14366 15986 14418 15998
rect 13906 15934 13918 15986
rect 13970 15983 13982 15986
rect 14130 15983 14142 15986
rect 13970 15937 14142 15983
rect 13970 15934 13982 15937
rect 14130 15934 14142 15937
rect 14194 15934 14206 15986
rect 7646 15922 7698 15934
rect 14366 15922 14418 15934
rect 14590 15986 14642 15998
rect 14590 15922 14642 15934
rect 18622 15986 18674 15998
rect 18622 15922 18674 15934
rect 18846 15986 18898 15998
rect 18846 15922 18898 15934
rect 19294 15986 19346 15998
rect 19294 15922 19346 15934
rect 19406 15986 19458 15998
rect 19406 15922 19458 15934
rect 22430 15986 22482 15998
rect 22430 15922 22482 15934
rect 23102 15986 23154 15998
rect 23102 15922 23154 15934
rect 23326 15986 23378 15998
rect 27246 15986 27298 15998
rect 23874 15934 23886 15986
rect 23938 15934 23950 15986
rect 25442 15934 25454 15986
rect 25506 15934 25518 15986
rect 23326 15922 23378 15934
rect 27246 15922 27298 15934
rect 27806 15986 27858 15998
rect 27806 15922 27858 15934
rect 29934 15986 29986 15998
rect 35198 15986 35250 15998
rect 34850 15934 34862 15986
rect 34914 15934 34926 15986
rect 35858 15934 35870 15986
rect 35922 15934 35934 15986
rect 38322 15934 38334 15986
rect 38386 15934 38398 15986
rect 29934 15922 29986 15934
rect 35198 15922 35250 15934
rect 4062 15874 4114 15886
rect 4062 15810 4114 15822
rect 7422 15874 7474 15886
rect 7422 15810 7474 15822
rect 14478 15874 14530 15886
rect 14478 15810 14530 15822
rect 14926 15874 14978 15886
rect 19070 15874 19122 15886
rect 27358 15874 27410 15886
rect 15250 15822 15262 15874
rect 15314 15822 15326 15874
rect 23986 15822 23998 15874
rect 24050 15822 24062 15874
rect 14926 15810 14978 15822
rect 19070 15810 19122 15822
rect 27358 15810 27410 15822
rect 28030 15874 28082 15886
rect 28030 15810 28082 15822
rect 30046 15874 30098 15886
rect 30046 15810 30098 15822
rect 31054 15874 31106 15886
rect 31054 15810 31106 15822
rect 1344 15706 39984 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 39984 15706
rect 1344 15620 39984 15654
rect 6078 15538 6130 15550
rect 3602 15486 3614 15538
rect 3666 15486 3678 15538
rect 6078 15474 6130 15486
rect 7758 15538 7810 15550
rect 7758 15474 7810 15486
rect 16046 15538 16098 15550
rect 16046 15474 16098 15486
rect 17726 15538 17778 15550
rect 17726 15474 17778 15486
rect 17838 15538 17890 15550
rect 17838 15474 17890 15486
rect 19742 15538 19794 15550
rect 19742 15474 19794 15486
rect 20078 15538 20130 15550
rect 20078 15474 20130 15486
rect 20750 15538 20802 15550
rect 23438 15538 23490 15550
rect 23090 15486 23102 15538
rect 23154 15486 23166 15538
rect 20750 15474 20802 15486
rect 23438 15474 23490 15486
rect 24334 15538 24386 15550
rect 24334 15474 24386 15486
rect 30606 15538 30658 15550
rect 30606 15474 30658 15486
rect 31278 15538 31330 15550
rect 31278 15474 31330 15486
rect 32062 15538 32114 15550
rect 32062 15474 32114 15486
rect 36318 15538 36370 15550
rect 36318 15474 36370 15486
rect 4846 15426 4898 15438
rect 4846 15362 4898 15374
rect 5070 15426 5122 15438
rect 5070 15362 5122 15374
rect 5630 15426 5682 15438
rect 5630 15362 5682 15374
rect 6302 15426 6354 15438
rect 8990 15426 9042 15438
rect 19854 15426 19906 15438
rect 7186 15374 7198 15426
rect 7250 15374 7262 15426
rect 10322 15374 10334 15426
rect 10386 15374 10398 15426
rect 12002 15374 12014 15426
rect 12066 15374 12078 15426
rect 14802 15374 14814 15426
rect 14866 15374 14878 15426
rect 29586 15374 29598 15426
rect 29650 15374 29662 15426
rect 35298 15374 35310 15426
rect 35362 15374 35374 15426
rect 6302 15362 6354 15374
rect 8990 15362 9042 15374
rect 19854 15362 19906 15374
rect 2830 15314 2882 15326
rect 2830 15250 2882 15262
rect 3054 15314 3106 15326
rect 4062 15314 4114 15326
rect 3266 15262 3278 15314
rect 3330 15262 3342 15314
rect 3054 15250 3106 15262
rect 4062 15250 4114 15262
rect 4174 15314 4226 15326
rect 4622 15314 4674 15326
rect 4386 15262 4398 15314
rect 4450 15262 4462 15314
rect 4174 15250 4226 15262
rect 4622 15250 4674 15262
rect 5294 15314 5346 15326
rect 5294 15250 5346 15262
rect 5854 15314 5906 15326
rect 5854 15250 5906 15262
rect 6862 15314 6914 15326
rect 6862 15250 6914 15262
rect 6974 15314 7026 15326
rect 17614 15314 17666 15326
rect 7298 15262 7310 15314
rect 7362 15262 7374 15314
rect 8530 15262 8542 15314
rect 8594 15262 8606 15314
rect 11554 15262 11566 15314
rect 11618 15262 11630 15314
rect 15586 15262 15598 15314
rect 15650 15262 15662 15314
rect 6974 15250 7026 15262
rect 17614 15250 17666 15262
rect 17950 15314 18002 15326
rect 19070 15314 19122 15326
rect 18162 15262 18174 15314
rect 18226 15262 18238 15314
rect 17950 15250 18002 15262
rect 19070 15250 19122 15262
rect 19294 15314 19346 15326
rect 31950 15314 32002 15326
rect 20290 15262 20302 15314
rect 20354 15262 20366 15314
rect 29810 15262 29822 15314
rect 29874 15262 29886 15314
rect 19294 15250 19346 15262
rect 31950 15250 32002 15262
rect 32174 15314 32226 15326
rect 32174 15250 32226 15262
rect 32622 15314 32674 15326
rect 32622 15250 32674 15262
rect 32958 15314 33010 15326
rect 36642 15262 36654 15314
rect 36706 15262 36718 15314
rect 32958 15250 33010 15262
rect 10110 15202 10162 15214
rect 18398 15202 18450 15214
rect 8082 15150 8094 15202
rect 8146 15150 8158 15202
rect 12674 15150 12686 15202
rect 12738 15150 12750 15202
rect 10110 15138 10162 15150
rect 18398 15138 18450 15150
rect 19518 15202 19570 15214
rect 19518 15138 19570 15150
rect 23774 15202 23826 15214
rect 37426 15150 37438 15202
rect 37490 15150 37502 15202
rect 39554 15150 39566 15202
rect 39618 15150 39630 15202
rect 23774 15138 23826 15150
rect 2718 15090 2770 15102
rect 2718 15026 2770 15038
rect 6190 15090 6242 15102
rect 6190 15026 6242 15038
rect 18846 15090 18898 15102
rect 18846 15026 18898 15038
rect 1344 14922 39984 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 39984 14922
rect 1344 14836 39984 14870
rect 3502 14754 3554 14766
rect 3502 14690 3554 14702
rect 3726 14754 3778 14766
rect 3726 14690 3778 14702
rect 18622 14754 18674 14766
rect 18622 14690 18674 14702
rect 23886 14754 23938 14766
rect 23886 14690 23938 14702
rect 4510 14642 4562 14654
rect 4510 14578 4562 14590
rect 11566 14642 11618 14654
rect 11566 14578 11618 14590
rect 19854 14642 19906 14654
rect 19854 14578 19906 14590
rect 29598 14642 29650 14654
rect 29598 14578 29650 14590
rect 30494 14642 30546 14654
rect 30494 14578 30546 14590
rect 30942 14642 30994 14654
rect 30942 14578 30994 14590
rect 31726 14642 31778 14654
rect 31726 14578 31778 14590
rect 12126 14530 12178 14542
rect 3938 14478 3950 14530
rect 4002 14478 4014 14530
rect 4946 14478 4958 14530
rect 5010 14478 5022 14530
rect 6738 14478 6750 14530
rect 6802 14478 6814 14530
rect 12126 14466 12178 14478
rect 12462 14530 12514 14542
rect 12462 14466 12514 14478
rect 12574 14530 12626 14542
rect 12574 14466 12626 14478
rect 15150 14530 15202 14542
rect 15150 14466 15202 14478
rect 18734 14530 18786 14542
rect 18734 14466 18786 14478
rect 18958 14530 19010 14542
rect 19966 14530 20018 14542
rect 22542 14530 22594 14542
rect 19170 14478 19182 14530
rect 19234 14478 19246 14530
rect 19506 14478 19518 14530
rect 19570 14478 19582 14530
rect 20178 14478 20190 14530
rect 20242 14478 20254 14530
rect 18958 14466 19010 14478
rect 19966 14466 20018 14478
rect 22542 14466 22594 14478
rect 29934 14530 29986 14542
rect 29934 14466 29986 14478
rect 3390 14418 3442 14430
rect 5854 14418 5906 14430
rect 4722 14366 4734 14418
rect 4786 14366 4798 14418
rect 3390 14354 3442 14366
rect 5854 14354 5906 14366
rect 6190 14418 6242 14430
rect 6190 14354 6242 14366
rect 6526 14418 6578 14430
rect 6526 14354 6578 14366
rect 13582 14418 13634 14430
rect 13582 14354 13634 14366
rect 23774 14418 23826 14430
rect 23774 14354 23826 14366
rect 29486 14418 29538 14430
rect 29486 14354 29538 14366
rect 29710 14418 29762 14430
rect 29710 14354 29762 14366
rect 30606 14418 30658 14430
rect 30606 14354 30658 14366
rect 31166 14418 31218 14430
rect 37314 14366 37326 14418
rect 37378 14366 37390 14418
rect 31166 14354 31218 14366
rect 11454 14306 11506 14318
rect 11454 14242 11506 14254
rect 11678 14306 11730 14318
rect 11678 14242 11730 14254
rect 12350 14306 12402 14318
rect 12350 14242 12402 14254
rect 12798 14306 12850 14318
rect 12798 14242 12850 14254
rect 13470 14306 13522 14318
rect 13470 14242 13522 14254
rect 14590 14306 14642 14318
rect 14590 14242 14642 14254
rect 17614 14306 17666 14318
rect 17614 14242 17666 14254
rect 17950 14306 18002 14318
rect 19742 14306 19794 14318
rect 26014 14306 26066 14318
rect 18274 14254 18286 14306
rect 18338 14254 18350 14306
rect 22866 14254 22878 14306
rect 22930 14254 22942 14306
rect 17950 14242 18002 14254
rect 19742 14242 19794 14254
rect 26014 14242 26066 14254
rect 28590 14306 28642 14318
rect 28590 14242 28642 14254
rect 30382 14306 30434 14318
rect 30382 14242 30434 14254
rect 31054 14306 31106 14318
rect 31054 14242 31106 14254
rect 39678 14306 39730 14318
rect 39678 14242 39730 14254
rect 1344 14138 39984 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 39984 14138
rect 1344 14052 39984 14086
rect 9662 13970 9714 13982
rect 9662 13906 9714 13918
rect 16270 13970 16322 13982
rect 16270 13906 16322 13918
rect 17614 13970 17666 13982
rect 17614 13906 17666 13918
rect 18174 13970 18226 13982
rect 18174 13906 18226 13918
rect 18398 13970 18450 13982
rect 18398 13906 18450 13918
rect 19966 13970 20018 13982
rect 19966 13906 20018 13918
rect 26126 13970 26178 13982
rect 26126 13906 26178 13918
rect 33182 13970 33234 13982
rect 33182 13906 33234 13918
rect 37102 13970 37154 13982
rect 37102 13906 37154 13918
rect 37214 13970 37266 13982
rect 37214 13906 37266 13918
rect 37326 13970 37378 13982
rect 37326 13906 37378 13918
rect 19182 13858 19234 13870
rect 2594 13806 2606 13858
rect 2658 13806 2670 13858
rect 19182 13794 19234 13806
rect 19406 13858 19458 13870
rect 19406 13794 19458 13806
rect 25342 13858 25394 13870
rect 25342 13794 25394 13806
rect 25902 13858 25954 13870
rect 37438 13858 37490 13870
rect 31266 13806 31278 13858
rect 31330 13806 31342 13858
rect 35858 13806 35870 13858
rect 35922 13806 35934 13858
rect 25902 13794 25954 13806
rect 37438 13794 37490 13806
rect 37662 13858 37714 13870
rect 37662 13794 37714 13806
rect 38110 13858 38162 13870
rect 38110 13794 38162 13806
rect 38334 13858 38386 13870
rect 38334 13794 38386 13806
rect 38558 13858 38610 13870
rect 38558 13794 38610 13806
rect 38782 13858 38834 13870
rect 38782 13794 38834 13806
rect 17950 13746 18002 13758
rect 1922 13694 1934 13746
rect 1986 13694 1998 13746
rect 12002 13694 12014 13746
rect 12066 13694 12078 13746
rect 17950 13682 18002 13694
rect 18510 13746 18562 13758
rect 18510 13682 18562 13694
rect 25790 13746 25842 13758
rect 38894 13746 38946 13758
rect 26338 13694 26350 13746
rect 26402 13694 26414 13746
rect 25790 13682 25842 13694
rect 38894 13682 38946 13694
rect 5182 13634 5234 13646
rect 4722 13582 4734 13634
rect 4786 13582 4798 13634
rect 5182 13570 5234 13582
rect 9550 13634 9602 13646
rect 22654 13634 22706 13646
rect 39342 13634 39394 13646
rect 15026 13582 15038 13634
rect 15090 13582 15102 13634
rect 37986 13582 37998 13634
rect 38050 13582 38062 13634
rect 9550 13570 9602 13582
rect 22654 13570 22706 13582
rect 39342 13570 39394 13582
rect 19070 13522 19122 13534
rect 19070 13458 19122 13470
rect 22766 13522 22818 13534
rect 22766 13458 22818 13470
rect 25454 13522 25506 13534
rect 25454 13458 25506 13470
rect 33742 13522 33794 13534
rect 33742 13458 33794 13470
rect 1344 13354 39984 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 39984 13354
rect 1344 13268 39984 13302
rect 19742 13186 19794 13198
rect 19742 13122 19794 13134
rect 38446 13186 38498 13198
rect 38446 13122 38498 13134
rect 7198 13074 7250 13086
rect 29262 13074 29314 13086
rect 10658 13022 10670 13074
rect 10722 13022 10734 13074
rect 18722 13022 18734 13074
rect 18786 13022 18798 13074
rect 23426 13022 23438 13074
rect 23490 13022 23502 13074
rect 24882 13022 24894 13074
rect 24946 13022 24958 13074
rect 7198 13010 7250 13022
rect 29262 13010 29314 13022
rect 33182 13074 33234 13086
rect 33182 13010 33234 13022
rect 34414 13074 34466 13086
rect 34414 13010 34466 13022
rect 36430 13074 36482 13086
rect 37650 13022 37662 13074
rect 37714 13022 37726 13074
rect 36430 13010 36482 13022
rect 8094 12962 8146 12974
rect 8094 12898 8146 12910
rect 19070 12962 19122 12974
rect 19070 12898 19122 12910
rect 22318 12962 22370 12974
rect 23886 12962 23938 12974
rect 26014 12962 26066 12974
rect 27694 12962 27746 12974
rect 22754 12910 22766 12962
rect 22818 12910 22830 12962
rect 25218 12910 25230 12962
rect 25282 12910 25294 12962
rect 26226 12910 26238 12962
rect 26290 12910 26302 12962
rect 27122 12910 27134 12962
rect 27186 12910 27198 12962
rect 22318 12898 22370 12910
rect 23886 12898 23938 12910
rect 26014 12898 26066 12910
rect 27694 12898 27746 12910
rect 28142 12962 28194 12974
rect 28142 12898 28194 12910
rect 29486 12962 29538 12974
rect 29486 12898 29538 12910
rect 29934 12962 29986 12974
rect 29934 12898 29986 12910
rect 30942 12962 30994 12974
rect 30942 12898 30994 12910
rect 31390 12962 31442 12974
rect 31390 12898 31442 12910
rect 32398 12962 32450 12974
rect 32398 12898 32450 12910
rect 32622 12962 32674 12974
rect 32622 12898 32674 12910
rect 33294 12962 33346 12974
rect 34190 12962 34242 12974
rect 33618 12910 33630 12962
rect 33682 12910 33694 12962
rect 33294 12898 33346 12910
rect 34190 12898 34242 12910
rect 34862 12962 34914 12974
rect 37202 12910 37214 12962
rect 37266 12910 37278 12962
rect 34862 12898 34914 12910
rect 8206 12850 8258 12862
rect 19294 12850 19346 12862
rect 11106 12798 11118 12850
rect 11170 12798 11182 12850
rect 12562 12798 12574 12850
rect 12626 12798 12638 12850
rect 8206 12786 8258 12798
rect 19294 12786 19346 12798
rect 19630 12850 19682 12862
rect 25678 12850 25730 12862
rect 30046 12850 30098 12862
rect 22978 12798 22990 12850
rect 23042 12798 23054 12850
rect 27458 12798 27470 12850
rect 27522 12798 27534 12850
rect 28466 12798 28478 12850
rect 28530 12798 28542 12850
rect 19630 12786 19682 12798
rect 25678 12786 25730 12798
rect 30046 12786 30098 12798
rect 30718 12850 30770 12862
rect 30718 12786 30770 12798
rect 31614 12850 31666 12862
rect 31614 12786 31666 12798
rect 31950 12850 32002 12862
rect 31950 12786 32002 12798
rect 32174 12850 32226 12862
rect 32174 12786 32226 12798
rect 33966 12850 34018 12862
rect 33966 12786 34018 12798
rect 34526 12850 34578 12862
rect 34526 12786 34578 12798
rect 37774 12850 37826 12862
rect 37774 12786 37826 12798
rect 37998 12850 38050 12862
rect 37998 12786 38050 12798
rect 38334 12850 38386 12862
rect 38334 12786 38386 12798
rect 38446 12850 38498 12862
rect 38446 12786 38498 12798
rect 7310 12738 7362 12750
rect 7310 12674 7362 12686
rect 8430 12738 8482 12750
rect 18734 12738 18786 12750
rect 12450 12686 12462 12738
rect 12514 12686 12526 12738
rect 8430 12674 8482 12686
rect 18734 12674 18786 12686
rect 18846 12738 18898 12750
rect 18846 12674 18898 12686
rect 19742 12738 19794 12750
rect 19742 12674 19794 12686
rect 30158 12738 30210 12750
rect 30158 12674 30210 12686
rect 31166 12738 31218 12750
rect 31166 12674 31218 12686
rect 31726 12738 31778 12750
rect 31726 12674 31778 12686
rect 32398 12738 32450 12750
rect 32398 12674 32450 12686
rect 33070 12738 33122 12750
rect 33070 12674 33122 12686
rect 34974 12738 35026 12750
rect 34974 12674 35026 12686
rect 35198 12738 35250 12750
rect 36978 12686 36990 12738
rect 37042 12686 37054 12738
rect 35198 12674 35250 12686
rect 1344 12570 39984 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 39984 12570
rect 1344 12484 39984 12518
rect 5630 12402 5682 12414
rect 8094 12402 8146 12414
rect 6626 12350 6638 12402
rect 6690 12350 6702 12402
rect 5630 12338 5682 12350
rect 8094 12338 8146 12350
rect 8766 12402 8818 12414
rect 8766 12338 8818 12350
rect 18286 12402 18338 12414
rect 18286 12338 18338 12350
rect 19294 12402 19346 12414
rect 19294 12338 19346 12350
rect 19406 12402 19458 12414
rect 25790 12402 25842 12414
rect 33406 12402 33458 12414
rect 21410 12350 21422 12402
rect 21474 12350 21486 12402
rect 30258 12350 30270 12402
rect 30322 12350 30334 12402
rect 19406 12338 19458 12350
rect 25790 12338 25842 12350
rect 33406 12338 33458 12350
rect 33630 12402 33682 12414
rect 33630 12338 33682 12350
rect 33742 12402 33794 12414
rect 33742 12338 33794 12350
rect 34862 12402 34914 12414
rect 34862 12338 34914 12350
rect 37102 12402 37154 12414
rect 37102 12338 37154 12350
rect 12462 12290 12514 12302
rect 3042 12238 3054 12290
rect 3106 12238 3118 12290
rect 12462 12226 12514 12238
rect 17950 12290 18002 12302
rect 17950 12226 18002 12238
rect 25342 12290 25394 12302
rect 26238 12290 26290 12302
rect 29150 12290 29202 12302
rect 25554 12238 25566 12290
rect 25618 12238 25630 12290
rect 26562 12238 26574 12290
rect 26626 12238 26638 12290
rect 25342 12226 25394 12238
rect 26238 12226 26290 12238
rect 29150 12226 29202 12238
rect 34078 12290 34130 12302
rect 34078 12226 34130 12238
rect 35870 12290 35922 12302
rect 35870 12226 35922 12238
rect 37214 12290 37266 12302
rect 37538 12238 37550 12290
rect 37602 12238 37614 12290
rect 37214 12226 37266 12238
rect 6302 12178 6354 12190
rect 2258 12126 2270 12178
rect 2322 12126 2334 12178
rect 6302 12114 6354 12126
rect 7758 12178 7810 12190
rect 7758 12114 7810 12126
rect 8094 12178 8146 12190
rect 8094 12114 8146 12126
rect 8318 12178 8370 12190
rect 8318 12114 8370 12126
rect 8542 12178 8594 12190
rect 8542 12114 8594 12126
rect 8878 12178 8930 12190
rect 10446 12178 10498 12190
rect 18622 12178 18674 12190
rect 19070 12178 19122 12190
rect 19966 12178 20018 12190
rect 9986 12126 9998 12178
rect 10050 12126 10062 12178
rect 17602 12126 17614 12178
rect 17666 12126 17678 12178
rect 18274 12126 18286 12178
rect 18338 12126 18350 12178
rect 18834 12126 18846 12178
rect 18898 12126 18910 12178
rect 19618 12126 19630 12178
rect 19682 12126 19694 12178
rect 8878 12114 8930 12126
rect 10446 12114 10498 12126
rect 18622 12114 18674 12126
rect 19070 12114 19122 12126
rect 19966 12114 20018 12126
rect 21758 12178 21810 12190
rect 21758 12114 21810 12126
rect 22206 12178 22258 12190
rect 22206 12114 22258 12126
rect 25790 12178 25842 12190
rect 25790 12114 25842 12126
rect 26014 12178 26066 12190
rect 36990 12178 37042 12190
rect 28130 12126 28142 12178
rect 28194 12126 28206 12178
rect 28578 12126 28590 12178
rect 28642 12126 28654 12178
rect 33170 12126 33182 12178
rect 33234 12126 33246 12178
rect 35074 12126 35086 12178
rect 35138 12126 35150 12178
rect 36194 12126 36206 12178
rect 36258 12126 36270 12178
rect 37426 12126 37438 12178
rect 37490 12126 37502 12178
rect 26014 12114 26066 12126
rect 36990 12114 37042 12126
rect 9550 12066 9602 12078
rect 17838 12066 17890 12078
rect 5170 12014 5182 12066
rect 5234 12014 5246 12066
rect 5394 12014 5406 12066
rect 5458 12014 5470 12066
rect 12562 12014 12574 12066
rect 12626 12014 12638 12066
rect 5409 11951 5455 12014
rect 9550 12002 9602 12014
rect 17838 12002 17890 12014
rect 24782 12066 24834 12078
rect 33954 12014 33966 12066
rect 34018 12014 34030 12066
rect 24782 12002 24834 12014
rect 12238 11954 12290 11966
rect 5842 11951 5854 11954
rect 5409 11905 5854 11951
rect 5842 11902 5854 11905
rect 5906 11951 5918 11954
rect 6066 11951 6078 11954
rect 5906 11905 6078 11951
rect 5906 11902 5918 11905
rect 6066 11902 6078 11905
rect 6130 11902 6142 11954
rect 7298 11902 7310 11954
rect 7362 11951 7374 11954
rect 7634 11951 7646 11954
rect 7362 11905 7646 11951
rect 7362 11902 7374 11905
rect 7634 11902 7646 11905
rect 7698 11902 7710 11954
rect 12238 11890 12290 11902
rect 34302 11954 34354 11966
rect 34302 11890 34354 11902
rect 36206 11954 36258 11966
rect 36206 11890 36258 11902
rect 1344 11786 39984 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 39984 11786
rect 1344 11700 39984 11734
rect 6414 11618 6466 11630
rect 6414 11554 6466 11566
rect 7422 11618 7474 11630
rect 22206 11618 22258 11630
rect 18834 11566 18846 11618
rect 18898 11566 18910 11618
rect 7422 11554 7474 11566
rect 22206 11554 22258 11566
rect 28254 11618 28306 11630
rect 28254 11554 28306 11566
rect 37886 11618 37938 11630
rect 37886 11554 37938 11566
rect 7310 11506 7362 11518
rect 29262 11506 29314 11518
rect 36430 11506 36482 11518
rect 13682 11454 13694 11506
rect 13746 11454 13758 11506
rect 15810 11454 15822 11506
rect 15874 11454 15886 11506
rect 22418 11454 22430 11506
rect 22482 11454 22494 11506
rect 32610 11454 32622 11506
rect 32674 11454 32686 11506
rect 7310 11442 7362 11454
rect 29262 11442 29314 11454
rect 36430 11442 36482 11454
rect 37102 11506 37154 11518
rect 37102 11442 37154 11454
rect 5854 11394 5906 11406
rect 11454 11394 11506 11406
rect 6738 11342 6750 11394
rect 6802 11342 6814 11394
rect 8642 11342 8654 11394
rect 8706 11342 8718 11394
rect 9538 11342 9550 11394
rect 9602 11342 9614 11394
rect 5854 11330 5906 11342
rect 11454 11330 11506 11342
rect 11790 11394 11842 11406
rect 12574 11394 12626 11406
rect 17726 11394 17778 11406
rect 19070 11394 19122 11406
rect 12002 11342 12014 11394
rect 12066 11342 12078 11394
rect 16594 11342 16606 11394
rect 16658 11342 16670 11394
rect 18610 11342 18622 11394
rect 18674 11342 18686 11394
rect 11790 11330 11842 11342
rect 12574 11330 12626 11342
rect 17726 11330 17778 11342
rect 19070 11330 19122 11342
rect 19406 11394 19458 11406
rect 19406 11330 19458 11342
rect 19630 11394 19682 11406
rect 19630 11330 19682 11342
rect 19966 11394 20018 11406
rect 19966 11330 20018 11342
rect 20750 11394 20802 11406
rect 23214 11394 23266 11406
rect 21858 11342 21870 11394
rect 21922 11342 21934 11394
rect 25778 11342 25790 11394
rect 25842 11342 25854 11394
rect 26674 11342 26686 11394
rect 26738 11342 26750 11394
rect 27458 11342 27470 11394
rect 27522 11342 27534 11394
rect 20750 11330 20802 11342
rect 23214 11330 23266 11342
rect 5966 11282 6018 11294
rect 11566 11282 11618 11294
rect 8082 11230 8094 11282
rect 8146 11230 8158 11282
rect 5966 11218 6018 11230
rect 11566 11218 11618 11230
rect 17950 11282 18002 11294
rect 17950 11218 18002 11230
rect 21646 11282 21698 11294
rect 22878 11282 22930 11294
rect 22754 11230 22766 11282
rect 22818 11230 22830 11282
rect 21646 11218 21698 11230
rect 22878 11218 22930 11230
rect 22990 11282 23042 11294
rect 22990 11218 23042 11230
rect 23662 11282 23714 11294
rect 28366 11282 28418 11294
rect 26562 11230 26574 11282
rect 26626 11230 26638 11282
rect 27346 11230 27358 11282
rect 27410 11230 27422 11282
rect 23662 11218 23714 11230
rect 28366 11218 28418 11230
rect 31726 11282 31778 11294
rect 31726 11218 31778 11230
rect 32286 11282 32338 11294
rect 38110 11282 38162 11294
rect 35522 11230 35534 11282
rect 35586 11230 35598 11282
rect 32286 11218 32338 11230
rect 38110 11218 38162 11230
rect 38558 11282 38610 11294
rect 38558 11218 38610 11230
rect 38670 11282 38722 11294
rect 38670 11218 38722 11230
rect 6190 11170 6242 11182
rect 6190 11106 6242 11118
rect 6526 11170 6578 11182
rect 6526 11106 6578 11118
rect 7198 11170 7250 11182
rect 12350 11170 12402 11182
rect 9650 11118 9662 11170
rect 9714 11118 9726 11170
rect 7198 11106 7250 11118
rect 12350 11106 12402 11118
rect 12462 11170 12514 11182
rect 12462 11106 12514 11118
rect 17054 11170 17106 11182
rect 17054 11106 17106 11118
rect 17838 11170 17890 11182
rect 17838 11106 17890 11118
rect 18174 11170 18226 11182
rect 19854 11170 19906 11182
rect 18946 11118 18958 11170
rect 19010 11118 19022 11170
rect 18174 11106 18226 11118
rect 19854 11106 19906 11118
rect 22094 11170 22146 11182
rect 22094 11106 22146 11118
rect 25230 11170 25282 11182
rect 25230 11106 25282 11118
rect 31838 11170 31890 11182
rect 31838 11106 31890 11118
rect 32062 11170 32114 11182
rect 32062 11106 32114 11118
rect 32510 11170 32562 11182
rect 32510 11106 32562 11118
rect 35870 11170 35922 11182
rect 35870 11106 35922 11118
rect 36990 11170 37042 11182
rect 36990 11106 37042 11118
rect 37214 11170 37266 11182
rect 37214 11106 37266 11118
rect 37438 11170 37490 11182
rect 37438 11106 37490 11118
rect 37998 11170 38050 11182
rect 37998 11106 38050 11118
rect 38894 11170 38946 11182
rect 38894 11106 38946 11118
rect 1344 11002 39984 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 39984 11002
rect 1344 10916 39984 10950
rect 7086 10834 7138 10846
rect 7086 10770 7138 10782
rect 7310 10834 7362 10846
rect 7310 10770 7362 10782
rect 8206 10834 8258 10846
rect 8206 10770 8258 10782
rect 18846 10834 18898 10846
rect 18846 10770 18898 10782
rect 19070 10834 19122 10846
rect 19070 10770 19122 10782
rect 19742 10834 19794 10846
rect 19742 10770 19794 10782
rect 20190 10834 20242 10846
rect 20190 10770 20242 10782
rect 29262 10834 29314 10846
rect 29262 10770 29314 10782
rect 35422 10834 35474 10846
rect 35422 10770 35474 10782
rect 37438 10834 37490 10846
rect 37438 10770 37490 10782
rect 37662 10834 37714 10846
rect 37662 10770 37714 10782
rect 38670 10834 38722 10846
rect 38670 10770 38722 10782
rect 7870 10722 7922 10734
rect 7870 10658 7922 10670
rect 7982 10722 8034 10734
rect 17950 10722 18002 10734
rect 16594 10670 16606 10722
rect 16658 10670 16670 10722
rect 7982 10658 8034 10670
rect 17950 10658 18002 10670
rect 18622 10722 18674 10734
rect 30158 10722 30210 10734
rect 28018 10670 28030 10722
rect 28082 10670 28094 10722
rect 18622 10658 18674 10670
rect 30158 10658 30210 10670
rect 33518 10722 33570 10734
rect 33518 10658 33570 10670
rect 38782 10722 38834 10734
rect 38782 10658 38834 10670
rect 7534 10610 7586 10622
rect 17726 10610 17778 10622
rect 13010 10558 13022 10610
rect 13074 10558 13086 10610
rect 7534 10546 7586 10558
rect 17726 10546 17778 10558
rect 18398 10610 18450 10622
rect 24558 10610 24610 10622
rect 21186 10558 21198 10610
rect 21250 10558 21262 10610
rect 18398 10546 18450 10558
rect 24558 10546 24610 10558
rect 26574 10610 26626 10622
rect 28590 10610 28642 10622
rect 27010 10558 27022 10610
rect 27074 10558 27086 10610
rect 27682 10558 27694 10610
rect 27746 10558 27758 10610
rect 26574 10546 26626 10558
rect 28590 10546 28642 10558
rect 29038 10610 29090 10622
rect 29038 10546 29090 10558
rect 29598 10610 29650 10622
rect 29598 10546 29650 10558
rect 29822 10610 29874 10622
rect 29822 10546 29874 10558
rect 31950 10610 32002 10622
rect 33070 10610 33122 10622
rect 32498 10558 32510 10610
rect 32562 10558 32574 10610
rect 31950 10546 32002 10558
rect 33070 10546 33122 10558
rect 33294 10610 33346 10622
rect 33294 10546 33346 10558
rect 33742 10610 33794 10622
rect 33742 10546 33794 10558
rect 34862 10610 34914 10622
rect 34862 10546 34914 10558
rect 35310 10610 35362 10622
rect 35310 10546 35362 10558
rect 35534 10610 35586 10622
rect 35534 10546 35586 10558
rect 36318 10610 36370 10622
rect 38558 10610 38610 10622
rect 36530 10558 36542 10610
rect 36594 10558 36606 10610
rect 37874 10558 37886 10610
rect 37938 10558 37950 10610
rect 38098 10558 38110 10610
rect 38162 10558 38174 10610
rect 39106 10558 39118 10610
rect 39170 10558 39182 10610
rect 36318 10546 36370 10558
rect 38558 10546 38610 10558
rect 7422 10498 7474 10510
rect 7422 10434 7474 10446
rect 18174 10498 18226 10510
rect 29150 10498 29202 10510
rect 21858 10446 21870 10498
rect 21922 10446 21934 10498
rect 23986 10446 23998 10498
rect 24050 10446 24062 10498
rect 28130 10446 28142 10498
rect 28194 10446 28206 10498
rect 18174 10434 18226 10446
rect 29150 10434 29202 10446
rect 30046 10498 30098 10510
rect 30046 10434 30098 10446
rect 33630 10498 33682 10510
rect 35970 10446 35982 10498
rect 36034 10446 36046 10498
rect 38210 10446 38222 10498
rect 38274 10446 38286 10498
rect 33630 10434 33682 10446
rect 18734 10386 18786 10398
rect 18734 10322 18786 10334
rect 32174 10386 32226 10398
rect 36978 10334 36990 10386
rect 37042 10334 37054 10386
rect 32174 10322 32226 10334
rect 1344 10218 39984 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 39984 10218
rect 1344 10132 39984 10166
rect 2830 10050 2882 10062
rect 2830 9986 2882 9998
rect 22318 10050 22370 10062
rect 22318 9986 22370 9998
rect 30494 10050 30546 10062
rect 30494 9986 30546 9998
rect 31726 10050 31778 10062
rect 31726 9986 31778 9998
rect 33518 10050 33570 10062
rect 33518 9986 33570 9998
rect 22430 9938 22482 9950
rect 23998 9938 24050 9950
rect 23090 9886 23102 9938
rect 23154 9886 23166 9938
rect 22430 9874 22482 9886
rect 23998 9874 24050 9886
rect 26350 9938 26402 9950
rect 26350 9874 26402 9886
rect 29486 9938 29538 9950
rect 32722 9886 32734 9938
rect 32786 9886 32798 9938
rect 29486 9874 29538 9886
rect 13582 9826 13634 9838
rect 3154 9774 3166 9826
rect 3218 9774 3230 9826
rect 8530 9774 8542 9826
rect 8594 9774 8606 9826
rect 9538 9774 9550 9826
rect 9602 9774 9614 9826
rect 13582 9762 13634 9774
rect 14142 9826 14194 9838
rect 14142 9762 14194 9774
rect 14254 9826 14306 9838
rect 14254 9762 14306 9774
rect 14702 9826 14754 9838
rect 26574 9826 26626 9838
rect 23538 9774 23550 9826
rect 23602 9774 23614 9826
rect 14702 9762 14754 9774
rect 26574 9762 26626 9774
rect 27022 9826 27074 9838
rect 27022 9762 27074 9774
rect 27582 9826 27634 9838
rect 27582 9762 27634 9774
rect 28254 9826 28306 9838
rect 29598 9826 29650 9838
rect 30718 9826 30770 9838
rect 29138 9774 29150 9826
rect 29202 9774 29214 9826
rect 29810 9774 29822 9826
rect 29874 9774 29886 9826
rect 28254 9762 28306 9774
rect 29598 9762 29650 9774
rect 30718 9762 30770 9774
rect 31278 9826 31330 9838
rect 31278 9762 31330 9774
rect 31838 9826 31890 9838
rect 31838 9762 31890 9774
rect 32398 9826 32450 9838
rect 37550 9826 37602 9838
rect 36978 9774 36990 9826
rect 37042 9774 37054 9826
rect 32398 9762 32450 9774
rect 37550 9762 37602 9774
rect 39230 9826 39282 9838
rect 39230 9762 39282 9774
rect 9998 9714 10050 9726
rect 18062 9714 18114 9726
rect 4050 9662 4062 9714
rect 4114 9662 4126 9714
rect 8306 9662 8318 9714
rect 8370 9662 8382 9714
rect 13906 9662 13918 9714
rect 13970 9662 13982 9714
rect 15026 9662 15038 9714
rect 15090 9662 15102 9714
rect 9998 9650 10050 9662
rect 18062 9650 18114 9662
rect 18398 9714 18450 9726
rect 27246 9714 27298 9726
rect 32174 9714 32226 9726
rect 19058 9662 19070 9714
rect 19122 9662 19134 9714
rect 27906 9662 27918 9714
rect 27970 9662 27982 9714
rect 28578 9662 28590 9714
rect 28642 9662 28654 9714
rect 18398 9650 18450 9662
rect 27246 9650 27298 9662
rect 32174 9650 32226 9662
rect 32622 9714 32674 9726
rect 39118 9714 39170 9726
rect 35634 9662 35646 9714
rect 35698 9662 35710 9714
rect 37986 9662 37998 9714
rect 38050 9662 38062 9714
rect 32622 9650 32674 9662
rect 39118 9650 39170 9662
rect 2942 9602 2994 9614
rect 2942 9538 2994 9550
rect 4398 9602 4450 9614
rect 4398 9538 4450 9550
rect 13358 9602 13410 9614
rect 13358 9538 13410 9550
rect 16942 9602 16994 9614
rect 16942 9538 16994 9550
rect 17390 9602 17442 9614
rect 17390 9538 17442 9550
rect 18734 9602 18786 9614
rect 18734 9538 18786 9550
rect 26798 9602 26850 9614
rect 26798 9538 26850 9550
rect 29374 9602 29426 9614
rect 31726 9602 31778 9614
rect 30146 9550 30158 9602
rect 30210 9550 30222 9602
rect 29374 9538 29426 9550
rect 31726 9538 31778 9550
rect 32734 9602 32786 9614
rect 32734 9538 32786 9550
rect 33294 9602 33346 9614
rect 33294 9538 33346 9550
rect 37214 9602 37266 9614
rect 37214 9538 37266 9550
rect 37326 9602 37378 9614
rect 37326 9538 37378 9550
rect 37438 9602 37490 9614
rect 37438 9538 37490 9550
rect 38334 9602 38386 9614
rect 38334 9538 38386 9550
rect 38894 9602 38946 9614
rect 38894 9538 38946 9550
rect 1344 9434 39984 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 39984 9434
rect 1344 9348 39984 9382
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 33630 9266 33682 9278
rect 33630 9202 33682 9214
rect 34302 9266 34354 9278
rect 34302 9202 34354 9214
rect 34526 9266 34578 9278
rect 34526 9202 34578 9214
rect 35758 9266 35810 9278
rect 35758 9202 35810 9214
rect 36318 9266 36370 9278
rect 38994 9214 39006 9266
rect 39058 9214 39070 9266
rect 36318 9202 36370 9214
rect 13918 9154 13970 9166
rect 31166 9154 31218 9166
rect 2482 9102 2494 9154
rect 2546 9102 2558 9154
rect 12226 9102 12238 9154
rect 12290 9102 12302 9154
rect 28690 9102 28702 9154
rect 28754 9102 28766 9154
rect 13918 9090 13970 9102
rect 31166 9090 31218 9102
rect 34078 9154 34130 9166
rect 34078 9090 34130 9102
rect 36990 9154 37042 9166
rect 37662 9154 37714 9166
rect 37314 9102 37326 9154
rect 37378 9102 37390 9154
rect 36990 9090 37042 9102
rect 37662 9090 37714 9102
rect 37998 9154 38050 9166
rect 37998 9090 38050 9102
rect 38334 9154 38386 9166
rect 38334 9090 38386 9102
rect 9438 9042 9490 9054
rect 1810 8990 1822 9042
rect 1874 8990 1886 9042
rect 9438 8978 9490 8990
rect 9886 9042 9938 9054
rect 9886 8978 9938 8990
rect 10110 9042 10162 9054
rect 24670 9042 24722 9054
rect 31278 9042 31330 9054
rect 13234 8990 13246 9042
rect 13298 8990 13310 9042
rect 25330 8990 25342 9042
rect 25394 8990 25406 9042
rect 10110 8978 10162 8990
rect 24670 8978 24722 8990
rect 31278 8978 31330 8990
rect 33070 9042 33122 9054
rect 33070 8978 33122 8990
rect 33518 9042 33570 9054
rect 33518 8978 33570 8990
rect 33742 9042 33794 9054
rect 33742 8978 33794 8990
rect 34638 9042 34690 9054
rect 34638 8978 34690 8990
rect 35870 9042 35922 9054
rect 35870 8978 35922 8990
rect 36206 9042 36258 9054
rect 38546 8990 38558 9042
rect 38610 8990 38622 9042
rect 39218 8990 39230 9042
rect 39282 8990 39294 9042
rect 36206 8978 36258 8990
rect 5070 8930 5122 8942
rect 31726 8930 31778 8942
rect 4610 8878 4622 8930
rect 4674 8878 4686 8930
rect 11778 8878 11790 8930
rect 11842 8878 11854 8930
rect 5070 8866 5122 8878
rect 31726 8866 31778 8878
rect 31166 8818 31218 8830
rect 31166 8754 31218 8766
rect 31614 8818 31666 8830
rect 31614 8754 31666 8766
rect 36318 8818 36370 8830
rect 36318 8754 36370 8766
rect 1344 8650 39984 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 39984 8650
rect 1344 8564 39984 8598
rect 13582 8482 13634 8494
rect 13582 8418 13634 8430
rect 34078 8482 34130 8494
rect 34078 8418 34130 8430
rect 12462 8370 12514 8382
rect 19854 8370 19906 8382
rect 3938 8318 3950 8370
rect 4002 8318 4014 8370
rect 16034 8318 16046 8370
rect 16098 8318 16110 8370
rect 16482 8318 16494 8370
rect 16546 8318 16558 8370
rect 18610 8318 18622 8370
rect 18674 8318 18686 8370
rect 12462 8306 12514 8318
rect 19854 8306 19906 8318
rect 29598 8370 29650 8382
rect 29598 8306 29650 8318
rect 30158 8370 30210 8382
rect 30158 8306 30210 8318
rect 31838 8370 31890 8382
rect 31838 8306 31890 8318
rect 37998 8370 38050 8382
rect 37998 8306 38050 8318
rect 12238 8258 12290 8270
rect 2370 8206 2382 8258
rect 2434 8206 2446 8258
rect 3714 8206 3726 8258
rect 3778 8206 3790 8258
rect 12238 8194 12290 8206
rect 12686 8258 12738 8270
rect 12686 8194 12738 8206
rect 13918 8258 13970 8270
rect 13918 8194 13970 8206
rect 15262 8258 15314 8270
rect 26238 8258 26290 8270
rect 15922 8206 15934 8258
rect 15986 8206 15998 8258
rect 19394 8206 19406 8258
rect 19458 8206 19470 8258
rect 15262 8194 15314 8206
rect 26238 8194 26290 8206
rect 29486 8258 29538 8270
rect 29486 8194 29538 8206
rect 29934 8258 29986 8270
rect 32622 8258 32674 8270
rect 30482 8206 30494 8258
rect 30546 8206 30558 8258
rect 31602 8206 31614 8258
rect 31666 8206 31678 8258
rect 29934 8194 29986 8206
rect 32622 8194 32674 8206
rect 33182 8258 33234 8270
rect 33182 8194 33234 8206
rect 33406 8258 33458 8270
rect 33406 8194 33458 8206
rect 33630 8258 33682 8270
rect 36542 8258 36594 8270
rect 34514 8206 34526 8258
rect 34578 8206 34590 8258
rect 33630 8194 33682 8206
rect 36542 8194 36594 8206
rect 37326 8258 37378 8270
rect 37326 8194 37378 8206
rect 37774 8258 37826 8270
rect 37774 8194 37826 8206
rect 38110 8258 38162 8270
rect 38882 8206 38894 8258
rect 38946 8206 38958 8258
rect 38110 8194 38162 8206
rect 2718 8146 2770 8158
rect 2718 8082 2770 8094
rect 3054 8146 3106 8158
rect 3054 8082 3106 8094
rect 5070 8146 5122 8158
rect 5070 8082 5122 8094
rect 5630 8146 5682 8158
rect 8878 8146 8930 8158
rect 5954 8094 5966 8146
rect 6018 8094 6030 8146
rect 5630 8082 5682 8094
rect 8878 8082 8930 8094
rect 12910 8146 12962 8158
rect 15150 8146 15202 8158
rect 14130 8094 14142 8146
rect 14194 8094 14206 8146
rect 14690 8094 14702 8146
rect 14754 8094 14766 8146
rect 12910 8082 12962 8094
rect 15150 8082 15202 8094
rect 15374 8146 15426 8158
rect 15374 8082 15426 8094
rect 29710 8146 29762 8158
rect 29710 8082 29762 8094
rect 31950 8146 32002 8158
rect 31950 8082 32002 8094
rect 32286 8146 32338 8158
rect 32286 8082 32338 8094
rect 32398 8146 32450 8158
rect 36206 8146 36258 8158
rect 34290 8094 34302 8146
rect 34354 8094 34366 8146
rect 32398 8082 32450 8094
rect 36206 8082 36258 8094
rect 36318 8146 36370 8158
rect 36318 8082 36370 8094
rect 36990 8146 37042 8158
rect 36990 8082 37042 8094
rect 37550 8146 37602 8158
rect 38994 8094 39006 8146
rect 39058 8094 39070 8146
rect 37550 8082 37602 8094
rect 2606 8034 2658 8046
rect 2606 7970 2658 7982
rect 4958 8034 5010 8046
rect 4958 7970 5010 7982
rect 8990 8034 9042 8046
rect 30718 8034 30770 8046
rect 26562 7982 26574 8034
rect 26626 7982 26638 8034
rect 8990 7970 9042 7982
rect 30718 7970 30770 7982
rect 30830 8034 30882 8046
rect 30830 7970 30882 7982
rect 30942 8034 30994 8046
rect 30942 7970 30994 7982
rect 31054 8034 31106 8046
rect 31054 7970 31106 7982
rect 37102 8034 37154 8046
rect 37102 7970 37154 7982
rect 38558 8034 38610 8046
rect 39218 7982 39230 8034
rect 39282 7982 39294 8034
rect 38558 7970 38610 7982
rect 1344 7866 39984 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 39984 7866
rect 1344 7780 39984 7814
rect 6638 7698 6690 7710
rect 6638 7634 6690 7646
rect 9662 7698 9714 7710
rect 9662 7634 9714 7646
rect 9886 7698 9938 7710
rect 9886 7634 9938 7646
rect 10558 7698 10610 7710
rect 10558 7634 10610 7646
rect 15822 7698 15874 7710
rect 15822 7634 15874 7646
rect 17726 7698 17778 7710
rect 17726 7634 17778 7646
rect 20750 7698 20802 7710
rect 20750 7634 20802 7646
rect 21422 7698 21474 7710
rect 29598 7698 29650 7710
rect 28578 7646 28590 7698
rect 28642 7646 28654 7698
rect 21422 7634 21474 7646
rect 29598 7634 29650 7646
rect 32174 7698 32226 7710
rect 32174 7634 32226 7646
rect 32398 7698 32450 7710
rect 32398 7634 32450 7646
rect 8094 7586 8146 7598
rect 2706 7534 2718 7586
rect 2770 7534 2782 7586
rect 8094 7522 8146 7534
rect 9774 7586 9826 7598
rect 9774 7522 9826 7534
rect 10670 7586 10722 7598
rect 10670 7522 10722 7534
rect 14478 7586 14530 7598
rect 24222 7586 24274 7598
rect 21746 7534 21758 7586
rect 21810 7534 21822 7586
rect 14478 7522 14530 7534
rect 24222 7522 24274 7534
rect 24446 7586 24498 7598
rect 24446 7522 24498 7534
rect 25678 7586 25730 7598
rect 25678 7522 25730 7534
rect 29038 7586 29090 7598
rect 29038 7522 29090 7534
rect 30158 7586 30210 7598
rect 30158 7522 30210 7534
rect 30830 7586 30882 7598
rect 35982 7586 36034 7598
rect 35634 7534 35646 7586
rect 35698 7534 35710 7586
rect 37650 7534 37662 7586
rect 37714 7534 37726 7586
rect 39218 7534 39230 7586
rect 39282 7534 39294 7586
rect 30830 7522 30882 7534
rect 35982 7522 36034 7534
rect 6750 7474 6802 7486
rect 7982 7474 8034 7486
rect 1922 7422 1934 7474
rect 1986 7422 1998 7474
rect 7298 7422 7310 7474
rect 7362 7422 7374 7474
rect 6750 7410 6802 7422
rect 7982 7410 8034 7422
rect 9998 7474 10050 7486
rect 13582 7474 13634 7486
rect 20974 7474 21026 7486
rect 10210 7422 10222 7474
rect 10274 7422 10286 7474
rect 13794 7422 13806 7474
rect 13858 7422 13870 7474
rect 9998 7410 10050 7422
rect 13582 7410 13634 7422
rect 20974 7410 21026 7422
rect 21086 7474 21138 7486
rect 21086 7410 21138 7422
rect 22094 7474 22146 7486
rect 22094 7410 22146 7422
rect 23774 7474 23826 7486
rect 23774 7410 23826 7422
rect 26126 7474 26178 7486
rect 26126 7410 26178 7422
rect 26350 7474 26402 7486
rect 27022 7474 27074 7486
rect 27918 7474 27970 7486
rect 29374 7474 29426 7486
rect 32510 7474 32562 7486
rect 26562 7422 26574 7474
rect 26626 7422 26638 7474
rect 27458 7422 27470 7474
rect 27522 7422 27534 7474
rect 28466 7422 28478 7474
rect 28530 7422 28542 7474
rect 28802 7422 28814 7474
rect 28866 7422 28878 7474
rect 31490 7422 31502 7474
rect 31554 7422 31566 7474
rect 26350 7410 26402 7422
rect 27022 7410 27074 7422
rect 27918 7410 27970 7422
rect 29374 7410 29426 7422
rect 32510 7410 32562 7422
rect 5294 7362 5346 7374
rect 4834 7310 4846 7362
rect 4898 7310 4910 7362
rect 5294 7298 5346 7310
rect 8654 7362 8706 7374
rect 28590 7362 28642 7374
rect 33854 7362 33906 7374
rect 22530 7310 22542 7362
rect 22594 7310 22606 7362
rect 29586 7310 29598 7362
rect 29650 7310 29662 7362
rect 31154 7310 31166 7362
rect 31218 7310 31230 7362
rect 8654 7298 8706 7310
rect 28590 7298 28642 7310
rect 33854 7298 33906 7310
rect 35310 7362 35362 7374
rect 36530 7310 36542 7362
rect 36594 7310 36606 7362
rect 38098 7310 38110 7362
rect 38162 7310 38174 7362
rect 35310 7298 35362 7310
rect 7310 7250 7362 7262
rect 7310 7186 7362 7198
rect 7646 7250 7698 7262
rect 7646 7186 7698 7198
rect 8094 7250 8146 7262
rect 8094 7186 8146 7198
rect 24110 7250 24162 7262
rect 24110 7186 24162 7198
rect 26014 7250 26066 7262
rect 26014 7186 26066 7198
rect 1344 7082 39984 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 39984 7082
rect 1344 6996 39984 7030
rect 29710 6914 29762 6926
rect 8978 6862 8990 6914
rect 9042 6911 9054 6914
rect 9762 6911 9774 6914
rect 9042 6865 9774 6911
rect 9042 6862 9054 6865
rect 9762 6862 9774 6865
rect 9826 6862 9838 6914
rect 29710 6850 29762 6862
rect 33294 6914 33346 6926
rect 33294 6850 33346 6862
rect 10558 6802 10610 6814
rect 36990 6802 37042 6814
rect 6850 6750 6862 6802
rect 6914 6750 6926 6802
rect 13682 6750 13694 6802
rect 13746 6750 13758 6802
rect 20738 6750 20750 6802
rect 20802 6750 20814 6802
rect 23538 6750 23550 6802
rect 23602 6750 23614 6802
rect 25666 6750 25678 6802
rect 25730 6750 25742 6802
rect 10558 6738 10610 6750
rect 36990 6738 37042 6750
rect 37102 6802 37154 6814
rect 38210 6750 38222 6802
rect 38274 6750 38286 6802
rect 37102 6738 37154 6750
rect 9326 6690 9378 6702
rect 7186 6638 7198 6690
rect 7250 6638 7262 6690
rect 9326 6626 9378 6638
rect 10334 6690 10386 6702
rect 10334 6626 10386 6638
rect 11230 6690 11282 6702
rect 11230 6626 11282 6638
rect 11678 6690 11730 6702
rect 14590 6690 14642 6702
rect 14130 6638 14142 6690
rect 14194 6638 14206 6690
rect 11678 6626 11730 6638
rect 14590 6626 14642 6638
rect 15374 6690 15426 6702
rect 16382 6690 16434 6702
rect 17054 6690 17106 6702
rect 34414 6690 34466 6702
rect 15586 6638 15598 6690
rect 15650 6638 15662 6690
rect 16706 6638 16718 6690
rect 16770 6638 16782 6690
rect 17826 6638 17838 6690
rect 17890 6638 17902 6690
rect 18610 6638 18622 6690
rect 18674 6638 18686 6690
rect 22866 6638 22878 6690
rect 22930 6638 22942 6690
rect 28130 6638 28142 6690
rect 28194 6638 28206 6690
rect 29362 6638 29374 6690
rect 29426 6638 29438 6690
rect 34738 6638 34750 6690
rect 34802 6638 34814 6690
rect 35746 6638 35758 6690
rect 35810 6638 35822 6690
rect 15374 6626 15426 6638
rect 16382 6626 16434 6638
rect 17054 6626 17106 6638
rect 34414 6626 34466 6638
rect 7758 6578 7810 6590
rect 15150 6578 15202 6590
rect 8418 6526 8430 6578
rect 8482 6526 8494 6578
rect 7758 6514 7810 6526
rect 15150 6514 15202 6526
rect 16942 6578 16994 6590
rect 29150 6578 29202 6590
rect 28354 6526 28366 6578
rect 28418 6526 28430 6578
rect 16942 6514 16994 6526
rect 29150 6514 29202 6526
rect 34302 6578 34354 6590
rect 37214 6578 37266 6590
rect 34850 6526 34862 6578
rect 34914 6526 34926 6578
rect 36306 6526 36318 6578
rect 36370 6526 36382 6578
rect 39106 6526 39118 6578
rect 39170 6526 39182 6578
rect 34302 6514 34354 6526
rect 37214 6514 37266 6526
rect 8094 6466 8146 6478
rect 8094 6402 8146 6414
rect 8878 6466 8930 6478
rect 10894 6466 10946 6478
rect 9986 6414 9998 6466
rect 10050 6414 10062 6466
rect 8878 6402 8930 6414
rect 10894 6402 10946 6414
rect 12686 6466 12738 6478
rect 12686 6402 12738 6414
rect 15038 6466 15090 6478
rect 15038 6402 15090 6414
rect 15262 6466 15314 6478
rect 26126 6466 26178 6478
rect 17490 6414 17502 6466
rect 17554 6414 17566 6466
rect 15262 6402 15314 6414
rect 26126 6402 26178 6414
rect 29598 6466 29650 6478
rect 29598 6402 29650 6414
rect 33406 6466 33458 6478
rect 33406 6402 33458 6414
rect 33518 6466 33570 6478
rect 37774 6466 37826 6478
rect 35858 6414 35870 6466
rect 35922 6414 35934 6466
rect 33518 6402 33570 6414
rect 37774 6402 37826 6414
rect 1344 6298 39984 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 39984 6298
rect 1344 6212 39984 6246
rect 4958 6130 5010 6142
rect 4958 6066 5010 6078
rect 5406 6130 5458 6142
rect 5406 6066 5458 6078
rect 10558 6130 10610 6142
rect 10558 6066 10610 6078
rect 11454 6130 11506 6142
rect 11454 6066 11506 6078
rect 12686 6130 12738 6142
rect 13918 6130 13970 6142
rect 13458 6078 13470 6130
rect 13522 6078 13534 6130
rect 12686 6066 12738 6078
rect 13918 6066 13970 6078
rect 16942 6130 16994 6142
rect 16942 6066 16994 6078
rect 18398 6130 18450 6142
rect 18398 6066 18450 6078
rect 22878 6130 22930 6142
rect 22878 6066 22930 6078
rect 24670 6130 24722 6142
rect 28242 6078 28254 6130
rect 28306 6078 28318 6130
rect 29250 6078 29262 6130
rect 29314 6078 29326 6130
rect 34178 6078 34190 6130
rect 34242 6078 34254 6130
rect 39106 6078 39118 6130
rect 39170 6078 39182 6130
rect 24670 6066 24722 6078
rect 5630 6018 5682 6030
rect 5630 5954 5682 5966
rect 5742 6018 5794 6030
rect 5742 5954 5794 5966
rect 11790 6018 11842 6030
rect 11790 5954 11842 5966
rect 14254 6018 14306 6030
rect 15822 6018 15874 6030
rect 15138 5966 15150 6018
rect 15202 5966 15214 6018
rect 14254 5954 14306 5966
rect 15822 5954 15874 5966
rect 25342 6018 25394 6030
rect 25342 5954 25394 5966
rect 25566 6018 25618 6030
rect 35746 5966 35758 6018
rect 35810 5966 35822 6018
rect 38322 5966 38334 6018
rect 38386 5966 38398 6018
rect 25566 5954 25618 5966
rect 10334 5906 10386 5918
rect 6066 5854 6078 5906
rect 6130 5854 6142 5906
rect 9650 5854 9662 5906
rect 9714 5854 9726 5906
rect 10334 5842 10386 5854
rect 11006 5906 11058 5918
rect 11006 5842 11058 5854
rect 13134 5906 13186 5918
rect 16158 5906 16210 5918
rect 15362 5854 15374 5906
rect 15426 5854 15438 5906
rect 13134 5842 13186 5854
rect 16158 5842 16210 5854
rect 16494 5906 16546 5918
rect 17838 5906 17890 5918
rect 22318 5906 22370 5918
rect 17378 5854 17390 5906
rect 17442 5854 17454 5906
rect 21858 5854 21870 5906
rect 21922 5854 21934 5906
rect 16494 5842 16546 5854
rect 17838 5842 17890 5854
rect 22318 5842 22370 5854
rect 28590 5906 28642 5918
rect 29026 5854 29038 5906
rect 29090 5854 29102 5906
rect 39330 5854 39342 5906
rect 39394 5854 39406 5906
rect 28590 5842 28642 5854
rect 9886 5794 9938 5806
rect 9886 5730 9938 5742
rect 10446 5794 10498 5806
rect 10446 5730 10498 5742
rect 12910 5794 12962 5806
rect 12910 5730 12962 5742
rect 16270 5794 16322 5806
rect 16270 5730 16322 5742
rect 17614 5794 17666 5806
rect 17614 5730 17666 5742
rect 21422 5794 21474 5806
rect 21422 5730 21474 5742
rect 32286 5794 32338 5806
rect 32286 5730 32338 5742
rect 33406 5794 33458 5806
rect 33406 5730 33458 5742
rect 33630 5794 33682 5806
rect 34514 5742 34526 5794
rect 34578 5742 34590 5794
rect 33630 5730 33682 5742
rect 7086 5682 7138 5694
rect 7086 5618 7138 5630
rect 9998 5682 10050 5694
rect 9998 5618 10050 5630
rect 14366 5682 14418 5694
rect 14366 5618 14418 5630
rect 17950 5682 18002 5694
rect 17950 5618 18002 5630
rect 25230 5682 25282 5694
rect 25230 5618 25282 5630
rect 33854 5682 33906 5694
rect 33854 5618 33906 5630
rect 36206 5682 36258 5694
rect 36206 5618 36258 5630
rect 1344 5514 39984 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 39984 5514
rect 1344 5428 39984 5462
rect 8878 5346 8930 5358
rect 8878 5282 8930 5294
rect 12798 5346 12850 5358
rect 12798 5282 12850 5294
rect 21646 5346 21698 5358
rect 21646 5282 21698 5294
rect 35870 5346 35922 5358
rect 35870 5282 35922 5294
rect 8990 5234 9042 5246
rect 17614 5234 17666 5246
rect 4722 5182 4734 5234
rect 4786 5182 4798 5234
rect 5618 5182 5630 5234
rect 5682 5182 5694 5234
rect 7746 5182 7758 5234
rect 7810 5182 7822 5234
rect 10322 5182 10334 5234
rect 10386 5182 10398 5234
rect 12450 5182 12462 5234
rect 12514 5182 12526 5234
rect 14130 5182 14142 5234
rect 14194 5182 14206 5234
rect 16258 5182 16270 5234
rect 16322 5182 16334 5234
rect 8990 5170 9042 5182
rect 17614 5170 17666 5182
rect 22094 5234 22146 5246
rect 27246 5234 27298 5246
rect 24658 5182 24670 5234
rect 24722 5182 24734 5234
rect 26786 5182 26798 5234
rect 26850 5182 26862 5234
rect 22094 5170 22146 5182
rect 27246 5170 27298 5182
rect 28590 5234 28642 5246
rect 39230 5234 39282 5246
rect 29250 5182 29262 5234
rect 29314 5182 29326 5234
rect 31378 5182 31390 5234
rect 31442 5182 31454 5234
rect 33394 5182 33406 5234
rect 33458 5182 33470 5234
rect 35522 5182 35534 5234
rect 35586 5182 35598 5234
rect 28590 5170 28642 5182
rect 39230 5170 39282 5182
rect 1922 5070 1934 5122
rect 1986 5070 1998 5122
rect 8530 5070 8542 5122
rect 8594 5070 8606 5122
rect 9202 5070 9214 5122
rect 9266 5070 9278 5122
rect 9538 5070 9550 5122
rect 9602 5070 9614 5122
rect 13570 5070 13582 5122
rect 13634 5070 13646 5122
rect 16930 5070 16942 5122
rect 16994 5070 17006 5122
rect 21298 5070 21310 5122
rect 21362 5070 21374 5122
rect 23874 5070 23886 5122
rect 23938 5070 23950 5122
rect 32050 5070 32062 5122
rect 32114 5070 32126 5122
rect 32610 5070 32622 5122
rect 32674 5070 32686 5122
rect 12910 5010 12962 5022
rect 2594 4958 2606 5010
rect 2658 4958 2670 5010
rect 12910 4946 12962 4958
rect 36094 5010 36146 5022
rect 37090 4958 37102 5010
rect 37154 4958 37166 5010
rect 36094 4946 36146 4958
rect 13806 4898 13858 4910
rect 13806 4834 13858 4846
rect 21534 4898 21586 4910
rect 21534 4834 21586 4846
rect 35982 4898 36034 4910
rect 35982 4834 36034 4846
rect 1344 4730 39984 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 39984 4730
rect 1344 4644 39984 4678
rect 3950 4562 4002 4574
rect 3950 4498 4002 4510
rect 4958 4562 5010 4574
rect 4958 4498 5010 4510
rect 5854 4562 5906 4574
rect 5854 4498 5906 4510
rect 5966 4562 6018 4574
rect 5966 4498 6018 4510
rect 22990 4562 23042 4574
rect 22990 4498 23042 4510
rect 29710 4562 29762 4574
rect 29710 4498 29762 4510
rect 32510 4562 32562 4574
rect 32510 4498 32562 4510
rect 17390 4450 17442 4462
rect 17390 4386 17442 4398
rect 18174 4450 18226 4462
rect 31950 4450 32002 4462
rect 21746 4398 21758 4450
rect 21810 4398 21822 4450
rect 26226 4398 26238 4450
rect 26290 4398 26302 4450
rect 18174 4386 18226 4398
rect 31950 4386 32002 4398
rect 32174 4450 32226 4462
rect 33506 4398 33518 4450
rect 33570 4398 33582 4450
rect 35186 4398 35198 4450
rect 35250 4398 35262 4450
rect 32174 4386 32226 4398
rect 28814 4338 28866 4350
rect 4722 4286 4734 4338
rect 4786 4286 4798 4338
rect 8978 4286 8990 4338
rect 9042 4286 9054 4338
rect 12002 4286 12014 4338
rect 12066 4286 12078 4338
rect 14914 4286 14926 4338
rect 14978 4286 14990 4338
rect 22530 4286 22542 4338
rect 22594 4286 22606 4338
rect 25442 4286 25454 4338
rect 25506 4286 25518 4338
rect 28814 4274 28866 4286
rect 29038 4338 29090 4350
rect 29038 4274 29090 4286
rect 29262 4338 29314 4350
rect 36642 4286 36654 4338
rect 36706 4286 36718 4338
rect 29262 4274 29314 4286
rect 3838 4226 3890 4238
rect 31502 4226 31554 4238
rect 7186 4174 7198 4226
rect 7250 4174 7262 4226
rect 19618 4174 19630 4226
rect 19682 4174 19694 4226
rect 28354 4174 28366 4226
rect 28418 4174 28430 4226
rect 34514 4174 34526 4226
rect 34578 4174 34590 4226
rect 36306 4174 36318 4226
rect 36370 4174 36382 4226
rect 37426 4174 37438 4226
rect 37490 4174 37502 4226
rect 39554 4174 39566 4226
rect 39618 4174 39630 4226
rect 3838 4162 3890 4174
rect 31502 4162 31554 4174
rect 6078 4114 6130 4126
rect 6078 4050 6130 4062
rect 10110 4114 10162 4126
rect 10110 4050 10162 4062
rect 13022 4114 13074 4126
rect 13022 4050 13074 4062
rect 1344 3946 39984 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 39984 3946
rect 1344 3860 39984 3894
rect 35534 3778 35586 3790
rect 35534 3714 35586 3726
rect 35870 3778 35922 3790
rect 35870 3714 35922 3726
rect 38782 3778 38834 3790
rect 38782 3714 38834 3726
rect 7758 3666 7810 3678
rect 7758 3602 7810 3614
rect 9550 3666 9602 3678
rect 28702 3666 28754 3678
rect 11218 3614 11230 3666
rect 11282 3614 11294 3666
rect 9550 3602 9602 3614
rect 28702 3602 28754 3614
rect 38894 3666 38946 3678
rect 38894 3602 38946 3614
rect 5070 3554 5122 3566
rect 13246 3554 13298 3566
rect 31278 3554 31330 3566
rect 5730 3502 5742 3554
rect 5794 3502 5806 3554
rect 8642 3502 8654 3554
rect 8706 3502 8718 3554
rect 12114 3502 12126 3554
rect 12178 3502 12190 3554
rect 14018 3502 14030 3554
rect 14082 3502 14094 3554
rect 16930 3502 16942 3554
rect 16994 3502 17006 3554
rect 5070 3490 5122 3502
rect 13246 3490 13298 3502
rect 31278 3490 31330 3502
rect 32622 3554 32674 3566
rect 32622 3490 32674 3502
rect 3166 3442 3218 3454
rect 3166 3378 3218 3390
rect 3390 3442 3442 3454
rect 3390 3378 3442 3390
rect 3726 3442 3778 3454
rect 3726 3378 3778 3390
rect 5518 3442 5570 3454
rect 31054 3442 31106 3454
rect 18498 3390 18510 3442
rect 18562 3390 18574 3442
rect 5518 3378 5570 3390
rect 31054 3378 31106 3390
rect 31614 3442 31666 3454
rect 31614 3378 31666 3390
rect 32286 3442 32338 3454
rect 39006 3442 39058 3454
rect 33394 3390 33406 3442
rect 33458 3390 33470 3442
rect 37986 3390 37998 3442
rect 38050 3390 38062 3442
rect 32286 3378 32338 3390
rect 39006 3378 39058 3390
rect 14814 3330 14866 3342
rect 14814 3266 14866 3278
rect 19854 3330 19906 3342
rect 19854 3266 19906 3278
rect 20862 3330 20914 3342
rect 20862 3266 20914 3278
rect 22206 3330 22258 3342
rect 22206 3266 22258 3278
rect 1344 3162 39984 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 39984 3162
rect 1344 3076 39984 3110
<< via1 >>
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 9998 39678 10050 39730
rect 18622 39678 18674 39730
rect 21310 39678 21362 39730
rect 12910 39566 12962 39618
rect 15710 39566 15762 39618
rect 24222 39566 24274 39618
rect 24670 39566 24722 39618
rect 12126 39454 12178 39506
rect 16494 39454 16546 39506
rect 23438 39454 23490 39506
rect 13582 39342 13634 39394
rect 15374 39342 15426 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 12126 39006 12178 39058
rect 16494 39006 16546 39058
rect 12014 38894 12066 38946
rect 15038 38894 15090 38946
rect 16606 38894 16658 38946
rect 17726 38894 17778 38946
rect 18286 38894 18338 38946
rect 22878 38894 22930 38946
rect 12686 38782 12738 38834
rect 13134 38782 13186 38834
rect 17390 38782 17442 38834
rect 18062 38782 18114 38834
rect 18174 38782 18226 38834
rect 18734 38782 18786 38834
rect 20190 38782 20242 38834
rect 20414 38782 20466 38834
rect 20974 38782 21026 38834
rect 21646 38782 21698 38834
rect 11678 38670 11730 38722
rect 13582 38670 13634 38722
rect 14702 38670 14754 38722
rect 17614 38670 17666 38722
rect 20638 38670 20690 38722
rect 21310 38670 21362 38722
rect 22430 38670 22482 38722
rect 12238 38558 12290 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18174 38222 18226 38274
rect 22654 38222 22706 38274
rect 9998 38110 10050 38162
rect 10558 38110 10610 38162
rect 13806 38110 13858 38162
rect 17166 38110 17218 38162
rect 20638 38110 20690 38162
rect 21870 38110 21922 38162
rect 22318 38110 22370 38162
rect 9662 37998 9714 38050
rect 11342 37998 11394 38050
rect 13918 37998 13970 38050
rect 14142 37998 14194 38050
rect 15934 37998 15986 38050
rect 16158 37998 16210 38050
rect 16382 37998 16434 38050
rect 17614 37998 17666 38050
rect 18398 37998 18450 38050
rect 18734 37998 18786 38050
rect 19854 37998 19906 38050
rect 21534 37998 21586 38050
rect 22654 37998 22706 38050
rect 11566 37886 11618 37938
rect 12238 37886 12290 37938
rect 12350 37886 12402 37938
rect 12686 37886 12738 37938
rect 13470 37886 13522 37938
rect 16606 37886 16658 37938
rect 18622 37886 18674 37938
rect 18958 37886 19010 37938
rect 19294 37886 19346 37938
rect 20078 37886 20130 37938
rect 20190 37886 20242 37938
rect 21310 37886 21362 37938
rect 21870 37886 21922 37938
rect 12798 37774 12850 37826
rect 13022 37774 13074 37826
rect 13694 37774 13746 37826
rect 16270 37774 16322 37826
rect 19630 37774 19682 37826
rect 20526 37774 20578 37826
rect 21758 37774 21810 37826
rect 23102 37774 23154 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 13470 37438 13522 37490
rect 13582 37438 13634 37490
rect 16830 37438 16882 37490
rect 17502 37438 17554 37490
rect 18062 37438 18114 37490
rect 18174 37438 18226 37490
rect 17390 37326 17442 37378
rect 17614 37326 17666 37378
rect 24446 37326 24498 37378
rect 28814 37326 28866 37378
rect 13358 37214 13410 37266
rect 13918 37214 13970 37266
rect 14366 37214 14418 37266
rect 16494 37214 16546 37266
rect 18286 37214 18338 37266
rect 18734 37214 18786 37266
rect 28254 37214 28306 37266
rect 19070 37102 19122 37154
rect 20414 37102 20466 37154
rect 22206 37102 22258 37154
rect 23550 37102 23602 37154
rect 24558 37102 24610 37154
rect 25342 37102 25394 37154
rect 27582 37102 27634 37154
rect 24670 36990 24722 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 17726 36542 17778 36594
rect 21422 36542 21474 36594
rect 25230 36542 25282 36594
rect 26238 36542 26290 36594
rect 13694 36430 13746 36482
rect 21646 36430 21698 36482
rect 21982 36430 22034 36482
rect 22318 36430 22370 36482
rect 23438 36430 23490 36482
rect 23886 36430 23938 36482
rect 24110 36430 24162 36482
rect 25342 36430 25394 36482
rect 13470 36318 13522 36370
rect 14030 36318 14082 36370
rect 23326 36318 23378 36370
rect 24782 36318 24834 36370
rect 25566 36318 25618 36370
rect 25790 36318 25842 36370
rect 12574 36206 12626 36258
rect 13806 36206 13858 36258
rect 22430 36206 22482 36258
rect 25230 36206 25282 36258
rect 33070 36206 33122 36258
rect 33406 36206 33458 36258
rect 33742 36206 33794 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 24110 35870 24162 35922
rect 12126 35758 12178 35810
rect 14478 35758 14530 35810
rect 14702 35758 14754 35810
rect 19854 35758 19906 35810
rect 22766 35758 22818 35810
rect 6190 35646 6242 35698
rect 13246 35646 13298 35698
rect 13694 35646 13746 35698
rect 14142 35646 14194 35698
rect 14254 35646 14306 35698
rect 19518 35646 19570 35698
rect 22206 35646 22258 35698
rect 24334 35646 24386 35698
rect 28254 35646 28306 35698
rect 6862 35534 6914 35586
rect 8990 35534 9042 35586
rect 9662 35534 9714 35586
rect 12350 35534 12402 35586
rect 13358 35534 13410 35586
rect 14366 35534 14418 35586
rect 21870 35534 21922 35586
rect 23214 35534 23266 35586
rect 28926 35534 28978 35586
rect 31054 35534 31106 35586
rect 31502 35534 31554 35586
rect 12014 35422 12066 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 11566 35086 11618 35138
rect 6414 34974 6466 35026
rect 8542 34974 8594 35026
rect 9662 34974 9714 35026
rect 12126 34974 12178 35026
rect 14254 34974 14306 35026
rect 17502 34974 17554 35026
rect 22878 34974 22930 35026
rect 28366 34974 28418 35026
rect 34414 34974 34466 35026
rect 35758 34974 35810 35026
rect 5630 34862 5682 34914
rect 8878 34862 8930 34914
rect 11566 34862 11618 34914
rect 12462 34862 12514 34914
rect 14142 34862 14194 34914
rect 14926 34862 14978 34914
rect 17278 34862 17330 34914
rect 17950 34862 18002 34914
rect 34750 34862 34802 34914
rect 11230 34750 11282 34802
rect 12910 34750 12962 34802
rect 13470 34750 13522 34802
rect 14814 34750 14866 34802
rect 17838 34750 17890 34802
rect 18398 34750 18450 34802
rect 34078 34750 34130 34802
rect 35422 34750 35474 34802
rect 9214 34638 9266 34690
rect 16942 34638 16994 34690
rect 23326 34638 23378 34690
rect 29374 34638 29426 34690
rect 35646 34638 35698 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 12462 34302 12514 34354
rect 12798 34302 12850 34354
rect 17614 34302 17666 34354
rect 18286 34302 18338 34354
rect 18622 34302 18674 34354
rect 19742 34302 19794 34354
rect 28926 34302 28978 34354
rect 29150 34302 29202 34354
rect 14702 34190 14754 34242
rect 16158 34190 16210 34242
rect 17838 34190 17890 34242
rect 29598 34190 29650 34242
rect 30830 34190 30882 34242
rect 32174 34190 32226 34242
rect 36542 34190 36594 34242
rect 13470 34078 13522 34130
rect 13918 34078 13970 34130
rect 14142 34078 14194 34130
rect 14590 34078 14642 34130
rect 15598 34078 15650 34130
rect 17278 34078 17330 34130
rect 18846 34078 18898 34130
rect 19182 34078 19234 34130
rect 19630 34078 19682 34130
rect 19854 34078 19906 34130
rect 25342 34078 25394 34130
rect 29262 34078 29314 34130
rect 29934 34078 29986 34130
rect 30270 34078 30322 34130
rect 30606 34078 30658 34130
rect 31726 34078 31778 34130
rect 34078 34078 34130 34130
rect 37214 34078 37266 34130
rect 10446 33966 10498 34018
rect 15934 33966 15986 34018
rect 20974 33966 21026 34018
rect 26014 33966 26066 34018
rect 28142 33966 28194 34018
rect 28814 33966 28866 34018
rect 30382 33966 30434 34018
rect 31278 33966 31330 34018
rect 34414 33966 34466 34018
rect 10558 33854 10610 33906
rect 17502 33854 17554 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 14030 33518 14082 33570
rect 7982 33406 8034 33458
rect 9214 33406 9266 33458
rect 15038 33406 15090 33458
rect 17390 33406 17442 33458
rect 19630 33406 19682 33458
rect 25566 33406 25618 33458
rect 25678 33406 25730 33458
rect 26126 33406 26178 33458
rect 31166 33406 31218 33458
rect 7310 33294 7362 33346
rect 9326 33294 9378 33346
rect 9998 33294 10050 33346
rect 10446 33294 10498 33346
rect 10894 33294 10946 33346
rect 14254 33294 14306 33346
rect 14926 33294 14978 33346
rect 15710 33294 15762 33346
rect 16270 33294 16322 33346
rect 16942 33294 16994 33346
rect 17278 33294 17330 33346
rect 17502 33294 17554 33346
rect 18622 33294 18674 33346
rect 19070 33294 19122 33346
rect 20078 33294 20130 33346
rect 20302 33294 20354 33346
rect 20526 33294 20578 33346
rect 21534 33294 21586 33346
rect 26686 33294 26738 33346
rect 29150 33294 29202 33346
rect 34862 33294 34914 33346
rect 35310 33294 35362 33346
rect 8206 33182 8258 33234
rect 9102 33182 9154 33234
rect 9550 33182 9602 33234
rect 11342 33182 11394 33234
rect 11454 33182 11506 33234
rect 12574 33182 12626 33234
rect 12798 33182 12850 33234
rect 20638 33182 20690 33234
rect 28590 33182 28642 33234
rect 35758 33182 35810 33234
rect 11118 33070 11170 33122
rect 12686 33070 12738 33122
rect 15598 33070 15650 33122
rect 15822 33070 15874 33122
rect 16718 33070 16770 33122
rect 21310 33070 21362 33122
rect 21422 33070 21474 33122
rect 21758 33070 21810 33122
rect 25454 33070 25506 33122
rect 26126 33070 26178 33122
rect 26238 33070 26290 33122
rect 26462 33070 26514 33122
rect 28142 33070 28194 33122
rect 28254 33070 28306 33122
rect 28478 33070 28530 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 17502 32734 17554 32786
rect 17726 32734 17778 32786
rect 18062 32734 18114 32786
rect 18286 32734 18338 32786
rect 19630 32734 19682 32786
rect 23550 32734 23602 32786
rect 25230 32734 25282 32786
rect 30382 32734 30434 32786
rect 32958 32734 33010 32786
rect 33182 32734 33234 32786
rect 35310 32734 35362 32786
rect 36318 32734 36370 32786
rect 11790 32622 11842 32674
rect 22318 32622 22370 32674
rect 25566 32622 25618 32674
rect 26126 32622 26178 32674
rect 26798 32622 26850 32674
rect 28702 32622 28754 32674
rect 35086 32622 35138 32674
rect 15486 32510 15538 32562
rect 17390 32510 17442 32562
rect 17950 32510 18002 32562
rect 19854 32510 19906 32562
rect 23102 32510 23154 32562
rect 26462 32510 26514 32562
rect 27470 32510 27522 32562
rect 28142 32510 28194 32562
rect 29486 32510 29538 32562
rect 29822 32510 29874 32562
rect 30158 32510 30210 32562
rect 30270 32510 30322 32562
rect 30494 32510 30546 32562
rect 31278 32510 31330 32562
rect 31838 32510 31890 32562
rect 32062 32510 32114 32562
rect 33294 32510 33346 32562
rect 34526 32510 34578 32562
rect 35422 32510 35474 32562
rect 35534 32510 35586 32562
rect 35758 32510 35810 32562
rect 36654 32510 36706 32562
rect 15934 32398 15986 32450
rect 19294 32398 19346 32450
rect 20190 32398 20242 32450
rect 31502 32398 31554 32450
rect 34750 32398 34802 32450
rect 37438 32398 37490 32450
rect 39566 32398 39618 32450
rect 19518 32286 19570 32338
rect 30942 32286 30994 32338
rect 32398 32286 32450 32338
rect 34190 32286 34242 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 30830 31950 30882 32002
rect 37326 31950 37378 32002
rect 8430 31838 8482 31890
rect 10446 31838 10498 31890
rect 12574 31838 12626 31890
rect 17166 31838 17218 31890
rect 35534 31838 35586 31890
rect 36990 31838 37042 31890
rect 8878 31726 8930 31778
rect 10110 31726 10162 31778
rect 11566 31726 11618 31778
rect 12126 31726 12178 31778
rect 14254 31726 14306 31778
rect 14926 31726 14978 31778
rect 16382 31726 16434 31778
rect 16942 31726 16994 31778
rect 17726 31726 17778 31778
rect 20526 31726 20578 31778
rect 31166 31726 31218 31778
rect 31502 31726 31554 31778
rect 31950 31726 32002 31778
rect 34414 31726 34466 31778
rect 35086 31726 35138 31778
rect 9326 31614 9378 31666
rect 9662 31614 9714 31666
rect 12014 31614 12066 31666
rect 14814 31614 14866 31666
rect 16158 31614 16210 31666
rect 17950 31614 18002 31666
rect 18062 31614 18114 31666
rect 20302 31614 20354 31666
rect 21758 31614 21810 31666
rect 34750 31614 34802 31666
rect 35534 31614 35586 31666
rect 11230 31502 11282 31554
rect 11790 31502 11842 31554
rect 14702 31502 14754 31554
rect 16270 31502 16322 31554
rect 16606 31502 16658 31554
rect 17278 31502 17330 31554
rect 17502 31502 17554 31554
rect 18622 31502 18674 31554
rect 18958 31502 19010 31554
rect 22094 31502 22146 31554
rect 30942 31502 30994 31554
rect 31614 31502 31666 31554
rect 31838 31502 31890 31554
rect 35310 31502 35362 31554
rect 35646 31502 35698 31554
rect 37214 31502 37266 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 14030 31166 14082 31218
rect 16942 31166 16994 31218
rect 29710 31166 29762 31218
rect 32286 31166 32338 31218
rect 33182 31166 33234 31218
rect 35870 31166 35922 31218
rect 7198 31054 7250 31106
rect 9662 31054 9714 31106
rect 17390 31054 17442 31106
rect 18846 31054 18898 31106
rect 23214 31054 23266 31106
rect 29934 31054 29986 31106
rect 30270 31054 30322 31106
rect 34302 31054 34354 31106
rect 37774 31054 37826 31106
rect 2830 30942 2882 30994
rect 6638 30942 6690 30994
rect 8542 30942 8594 30994
rect 8766 30942 8818 30994
rect 8990 30942 9042 30994
rect 9550 30942 9602 30994
rect 9886 30942 9938 30994
rect 10110 30942 10162 30994
rect 13806 30942 13858 30994
rect 16046 30942 16098 30994
rect 16270 30942 16322 30994
rect 16494 30942 16546 30994
rect 17614 30942 17666 30994
rect 17838 30942 17890 30994
rect 22654 30942 22706 30994
rect 23662 30942 23714 30994
rect 29598 30942 29650 30994
rect 30382 30942 30434 30994
rect 31838 30942 31890 30994
rect 32062 30942 32114 30994
rect 32398 30942 32450 30994
rect 33406 30942 33458 30994
rect 35758 30942 35810 30994
rect 36542 30942 36594 30994
rect 36990 30942 37042 30994
rect 37550 30942 37602 30994
rect 3614 30830 3666 30882
rect 5742 30830 5794 30882
rect 6414 30830 6466 30882
rect 24110 30830 24162 30882
rect 32174 30830 32226 30882
rect 34078 30830 34130 30882
rect 10558 30718 10610 30770
rect 18734 30718 18786 30770
rect 30270 30718 30322 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 13918 30382 13970 30434
rect 27806 30382 27858 30434
rect 32174 30382 32226 30434
rect 11790 30270 11842 30322
rect 23662 30270 23714 30322
rect 23998 30270 24050 30322
rect 26462 30270 26514 30322
rect 27694 30270 27746 30322
rect 36318 30270 36370 30322
rect 37326 30270 37378 30322
rect 5966 30158 6018 30210
rect 6414 30158 6466 30210
rect 8094 30158 8146 30210
rect 8654 30158 8706 30210
rect 8766 30158 8818 30210
rect 10222 30158 10274 30210
rect 10558 30158 10610 30210
rect 11678 30158 11730 30210
rect 14366 30158 14418 30210
rect 14926 30158 14978 30210
rect 17054 30158 17106 30210
rect 17502 30158 17554 30210
rect 18398 30158 18450 30210
rect 24222 30158 24274 30210
rect 26126 30158 26178 30210
rect 27470 30158 27522 30210
rect 29934 30158 29986 30210
rect 30942 30158 30994 30210
rect 31166 30158 31218 30210
rect 31390 30158 31442 30210
rect 31502 30158 31554 30210
rect 35870 30158 35922 30210
rect 36878 30158 36930 30210
rect 37550 30158 37602 30210
rect 37662 30158 37714 30210
rect 10782 30046 10834 30098
rect 11230 30046 11282 30098
rect 13694 30046 13746 30098
rect 14478 30046 14530 30098
rect 17390 30046 17442 30098
rect 18174 30046 18226 30098
rect 18734 30046 18786 30098
rect 27022 30046 27074 30098
rect 27358 30046 27410 30098
rect 30158 30046 30210 30098
rect 31950 30046 32002 30098
rect 38670 30046 38722 30098
rect 39230 30046 39282 30098
rect 39342 30046 39394 30098
rect 6750 29934 6802 29986
rect 10894 29934 10946 29986
rect 13806 29934 13858 29986
rect 14254 29934 14306 29986
rect 16718 29934 16770 29986
rect 17166 29934 17218 29986
rect 18398 29934 18450 29986
rect 24894 29934 24946 29986
rect 31278 29934 31330 29986
rect 32510 29934 32562 29986
rect 36206 29934 36258 29986
rect 36430 29934 36482 29986
rect 39006 29934 39058 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 5182 29598 5234 29650
rect 10446 29598 10498 29650
rect 10558 29598 10610 29650
rect 11342 29598 11394 29650
rect 13918 29598 13970 29650
rect 14478 29598 14530 29650
rect 17390 29598 17442 29650
rect 26798 29598 26850 29650
rect 28254 29598 28306 29650
rect 31390 29598 31442 29650
rect 36878 29598 36930 29650
rect 36990 29598 37042 29650
rect 11566 29486 11618 29538
rect 17614 29486 17666 29538
rect 17726 29486 17778 29538
rect 18174 29486 18226 29538
rect 19070 29486 19122 29538
rect 19182 29486 19234 29538
rect 26350 29486 26402 29538
rect 26462 29486 26514 29538
rect 26574 29486 26626 29538
rect 26686 29486 26738 29538
rect 28366 29486 28418 29538
rect 31166 29486 31218 29538
rect 37774 29486 37826 29538
rect 37998 29486 38050 29538
rect 1934 29374 1986 29426
rect 10110 29374 10162 29426
rect 10334 29374 10386 29426
rect 10670 29374 10722 29426
rect 11006 29374 11058 29426
rect 14030 29374 14082 29426
rect 14254 29374 14306 29426
rect 14590 29374 14642 29426
rect 19406 29374 19458 29426
rect 20638 29374 20690 29426
rect 23998 29374 24050 29426
rect 27134 29374 27186 29426
rect 27358 29374 27410 29426
rect 27918 29374 27970 29426
rect 28478 29374 28530 29426
rect 30942 29374 30994 29426
rect 31614 29374 31666 29426
rect 36766 29374 36818 29426
rect 37438 29374 37490 29426
rect 2606 29262 2658 29314
rect 4734 29262 4786 29314
rect 21310 29262 21362 29314
rect 23438 29262 23490 29314
rect 30606 29262 30658 29314
rect 37662 29262 37714 29314
rect 11678 29150 11730 29202
rect 13918 29150 13970 29202
rect 27694 29150 27746 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 10446 28814 10498 28866
rect 11006 28814 11058 28866
rect 11790 28814 11842 28866
rect 29822 28814 29874 28866
rect 32510 28814 32562 28866
rect 8542 28702 8594 28754
rect 9438 28702 9490 28754
rect 10670 28702 10722 28754
rect 11566 28702 11618 28754
rect 13694 28702 13746 28754
rect 22766 28702 22818 28754
rect 31166 28702 31218 28754
rect 33406 28702 33458 28754
rect 7982 28590 8034 28642
rect 8430 28590 8482 28642
rect 8654 28590 8706 28642
rect 9214 28590 9266 28642
rect 9550 28590 9602 28642
rect 10222 28590 10274 28642
rect 10894 28590 10946 28642
rect 12014 28590 12066 28642
rect 12126 28590 12178 28642
rect 13470 28590 13522 28642
rect 13918 28590 13970 28642
rect 14030 28590 14082 28642
rect 14366 28590 14418 28642
rect 14814 28590 14866 28642
rect 20190 28590 20242 28642
rect 20750 28590 20802 28642
rect 27470 28590 27522 28642
rect 28142 28590 28194 28642
rect 28366 28590 28418 28642
rect 31390 28590 31442 28642
rect 31614 28590 31666 28642
rect 32846 28590 32898 28642
rect 8990 28478 9042 28530
rect 12350 28478 12402 28530
rect 20414 28478 20466 28530
rect 23774 28478 23826 28530
rect 27134 28478 27186 28530
rect 28702 28478 28754 28530
rect 29710 28478 29762 28530
rect 30830 28478 30882 28530
rect 9774 28366 9826 28418
rect 14030 28366 14082 28418
rect 26798 28366 26850 28418
rect 26910 28366 26962 28418
rect 28590 28366 28642 28418
rect 29822 28366 29874 28418
rect 30494 28366 30546 28418
rect 32622 28366 32674 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 8990 28030 9042 28082
rect 11230 28030 11282 28082
rect 15374 28030 15426 28082
rect 21758 28030 21810 28082
rect 22654 28030 22706 28082
rect 8542 27918 8594 27970
rect 10334 27918 10386 27970
rect 21646 27918 21698 27970
rect 21982 27918 22034 27970
rect 23102 27918 23154 27970
rect 33630 27918 33682 27970
rect 37214 27918 37266 27970
rect 3838 27806 3890 27858
rect 7870 27806 7922 27858
rect 8430 27806 8482 27858
rect 10446 27806 10498 27858
rect 10894 27806 10946 27858
rect 22206 27806 22258 27858
rect 26910 27806 26962 27858
rect 28254 27806 28306 27858
rect 33406 27806 33458 27858
rect 37662 27806 37714 27858
rect 4622 27694 4674 27746
rect 6750 27694 6802 27746
rect 26238 27694 26290 27746
rect 31838 27694 31890 27746
rect 35534 27694 35586 27746
rect 38110 27694 38162 27746
rect 11118 27582 11170 27634
rect 15038 27582 15090 27634
rect 15374 27582 15426 27634
rect 22318 27582 22370 27634
rect 22878 27582 22930 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 4622 27134 4674 27186
rect 8878 27134 8930 27186
rect 9774 27134 9826 27186
rect 10446 27134 10498 27186
rect 11118 27134 11170 27186
rect 11902 27134 11954 27186
rect 18846 27134 18898 27186
rect 25902 27134 25954 27186
rect 26686 27134 26738 27186
rect 29374 27134 29426 27186
rect 30158 27134 30210 27186
rect 31838 27134 31890 27186
rect 33966 27134 34018 27186
rect 35198 27134 35250 27186
rect 37326 27134 37378 27186
rect 1822 27022 1874 27074
rect 9326 27022 9378 27074
rect 11566 27022 11618 27074
rect 13470 27022 13522 27074
rect 15038 27022 15090 27074
rect 16046 27022 16098 27074
rect 25230 27022 25282 27074
rect 26798 27022 26850 27074
rect 29486 27022 29538 27074
rect 34750 27022 34802 27074
rect 35870 27022 35922 27074
rect 35982 27022 36034 27074
rect 36094 27022 36146 27074
rect 37438 27022 37490 27074
rect 38334 27022 38386 27074
rect 39230 27022 39282 27074
rect 2494 26910 2546 26962
rect 5070 26910 5122 26962
rect 7198 26910 7250 26962
rect 13806 26910 13858 26962
rect 14814 26910 14866 26962
rect 16718 26910 16770 26962
rect 26126 26910 26178 26962
rect 27470 26910 27522 26962
rect 31502 26910 31554 26962
rect 36206 26910 36258 26962
rect 36430 26910 36482 26962
rect 36990 26910 37042 26962
rect 38558 26910 38610 26962
rect 39006 26910 39058 26962
rect 15598 26798 15650 26850
rect 38446 26798 38498 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 27246 26462 27298 26514
rect 27470 26462 27522 26514
rect 27918 26462 27970 26514
rect 34638 26462 34690 26514
rect 34974 26462 35026 26514
rect 35310 26462 35362 26514
rect 35870 26462 35922 26514
rect 6638 26350 6690 26402
rect 27806 26350 27858 26402
rect 37438 26350 37490 26402
rect 6414 26238 6466 26290
rect 13022 26238 13074 26290
rect 20078 26238 20130 26290
rect 25454 26238 25506 26290
rect 26798 26238 26850 26290
rect 27022 26238 27074 26290
rect 28142 26238 28194 26290
rect 28926 26238 28978 26290
rect 30718 26238 30770 26290
rect 31166 26238 31218 26290
rect 36206 26238 36258 26290
rect 36318 26238 36370 26290
rect 36766 26238 36818 26290
rect 16270 26126 16322 26178
rect 17502 26126 17554 26178
rect 20750 26126 20802 26178
rect 22878 26126 22930 26178
rect 23326 26126 23378 26178
rect 25790 26126 25842 26178
rect 27246 26126 27298 26178
rect 29150 26126 29202 26178
rect 29710 26126 29762 26178
rect 31390 26126 31442 26178
rect 39566 26126 39618 26178
rect 26126 26014 26178 26066
rect 28254 26014 28306 26066
rect 28702 26014 28754 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 3166 25678 3218 25730
rect 13470 25566 13522 25618
rect 15598 25566 15650 25618
rect 20750 25566 20802 25618
rect 26238 25566 26290 25618
rect 30158 25566 30210 25618
rect 7310 25454 7362 25506
rect 16270 25454 16322 25506
rect 17950 25454 18002 25506
rect 25790 25454 25842 25506
rect 26126 25454 26178 25506
rect 27246 25454 27298 25506
rect 27694 25454 27746 25506
rect 30046 25454 30098 25506
rect 3502 25342 3554 25394
rect 7534 25342 7586 25394
rect 7982 25342 8034 25394
rect 18622 25342 18674 25394
rect 26686 25342 26738 25394
rect 28366 25342 28418 25394
rect 29374 25342 29426 25394
rect 3278 25230 3330 25282
rect 8206 25230 8258 25282
rect 16830 25230 16882 25282
rect 17502 25230 17554 25282
rect 22766 25230 22818 25282
rect 27246 25230 27298 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 2382 24894 2434 24946
rect 22094 24894 22146 24946
rect 2270 24782 2322 24834
rect 4286 24782 4338 24834
rect 5966 24782 6018 24834
rect 6526 24782 6578 24834
rect 6862 24782 6914 24834
rect 27806 24782 27858 24834
rect 27918 24782 27970 24834
rect 28142 24782 28194 24834
rect 28366 24782 28418 24834
rect 28926 24782 28978 24834
rect 29374 24782 29426 24834
rect 2494 24670 2546 24722
rect 2830 24670 2882 24722
rect 3502 24670 3554 24722
rect 4398 24670 4450 24722
rect 4958 24670 5010 24722
rect 5742 24670 5794 24722
rect 18286 24670 18338 24722
rect 18846 24670 18898 24722
rect 19294 24670 19346 24722
rect 22430 24670 22482 24722
rect 22878 24670 22930 24722
rect 24670 24670 24722 24722
rect 25566 24670 25618 24722
rect 26238 24670 26290 24722
rect 27358 24670 27410 24722
rect 27582 24670 27634 24722
rect 28590 24670 28642 24722
rect 29150 24670 29202 24722
rect 29710 24670 29762 24722
rect 30046 24670 30098 24722
rect 36094 24670 36146 24722
rect 37102 24670 37154 24722
rect 3614 24558 3666 24610
rect 23326 24558 23378 24610
rect 25790 24558 25842 24610
rect 29038 24558 29090 24610
rect 29822 24558 29874 24610
rect 35870 24558 35922 24610
rect 36766 24558 36818 24610
rect 37662 24558 37714 24610
rect 27022 24446 27074 24498
rect 27134 24446 27186 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 15262 24110 15314 24162
rect 15710 24110 15762 24162
rect 5630 23998 5682 24050
rect 11342 23998 11394 24050
rect 12798 23998 12850 24050
rect 15262 23998 15314 24050
rect 15710 23998 15762 24050
rect 18958 23998 19010 24050
rect 24558 23998 24610 24050
rect 35198 23998 35250 24050
rect 35982 23998 36034 24050
rect 36430 23998 36482 24050
rect 37550 23998 37602 24050
rect 3726 23886 3778 23938
rect 4062 23886 4114 23938
rect 4398 23886 4450 23938
rect 4622 23886 4674 23938
rect 4846 23886 4898 23938
rect 8430 23886 8482 23938
rect 11902 23886 11954 23938
rect 16046 23886 16098 23938
rect 21758 23886 21810 23938
rect 25006 23886 25058 23938
rect 26574 23886 26626 23938
rect 31950 23886 32002 23938
rect 32286 23886 32338 23938
rect 37102 23886 37154 23938
rect 37438 23886 37490 23938
rect 5966 23774 6018 23826
rect 7646 23774 7698 23826
rect 7870 23774 7922 23826
rect 9102 23774 9154 23826
rect 13694 23774 13746 23826
rect 16830 23774 16882 23826
rect 22430 23774 22482 23826
rect 26686 23774 26738 23826
rect 26910 23774 26962 23826
rect 33070 23774 33122 23826
rect 37550 23774 37602 23826
rect 3838 23662 3890 23714
rect 4734 23662 4786 23714
rect 5742 23662 5794 23714
rect 7758 23662 7810 23714
rect 12910 23662 12962 23714
rect 13918 23662 13970 23714
rect 14030 23662 14082 23714
rect 14142 23662 14194 23714
rect 19518 23662 19570 23714
rect 31390 23662 31442 23714
rect 37214 23662 37266 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 4734 23326 4786 23378
rect 16270 23326 16322 23378
rect 17502 23326 17554 23378
rect 18622 23326 18674 23378
rect 19518 23326 19570 23378
rect 22878 23326 22930 23378
rect 27582 23326 27634 23378
rect 31502 23326 31554 23378
rect 3166 23214 3218 23266
rect 6862 23214 6914 23266
rect 8430 23214 8482 23266
rect 16158 23214 16210 23266
rect 19070 23214 19122 23266
rect 22542 23214 22594 23266
rect 26910 23214 26962 23266
rect 31278 23214 31330 23266
rect 35422 23214 35474 23266
rect 37102 23214 37154 23266
rect 3502 23102 3554 23154
rect 5294 23102 5346 23154
rect 7198 23102 7250 23154
rect 7982 23102 8034 23154
rect 15262 23102 15314 23154
rect 15598 23102 15650 23154
rect 15934 23102 15986 23154
rect 17390 23102 17442 23154
rect 17726 23102 17778 23154
rect 18174 23102 18226 23154
rect 18510 23102 18562 23154
rect 18846 23102 18898 23154
rect 19406 23102 19458 23154
rect 19630 23102 19682 23154
rect 19966 23102 20018 23154
rect 22766 23102 22818 23154
rect 22990 23102 23042 23154
rect 27246 23102 27298 23154
rect 27694 23102 27746 23154
rect 28590 23102 28642 23154
rect 31166 23102 31218 23154
rect 31614 23102 31666 23154
rect 32062 23102 32114 23154
rect 32286 23102 32338 23154
rect 37326 23102 37378 23154
rect 38222 23102 38274 23154
rect 38558 23102 38610 23154
rect 38894 23102 38946 23154
rect 12462 22990 12514 23042
rect 14590 22990 14642 23042
rect 16830 22990 16882 23042
rect 20414 22990 20466 23042
rect 22094 22990 22146 23042
rect 23438 22990 23490 23042
rect 23886 22990 23938 23042
rect 28478 22990 28530 23042
rect 30382 22990 30434 23042
rect 30830 22990 30882 23042
rect 31838 22990 31890 23042
rect 34078 22990 34130 23042
rect 37438 22990 37490 23042
rect 39118 22990 39170 23042
rect 5070 22878 5122 22930
rect 8094 22878 8146 22930
rect 8318 22878 8370 22930
rect 17950 22878 18002 22930
rect 27470 22878 27522 22930
rect 28254 22878 28306 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 7646 22542 7698 22594
rect 14030 22542 14082 22594
rect 30494 22542 30546 22594
rect 8206 22430 8258 22482
rect 14478 22430 14530 22482
rect 16942 22430 16994 22482
rect 27694 22430 27746 22482
rect 30270 22430 30322 22482
rect 35758 22430 35810 22482
rect 36990 22430 37042 22482
rect 37326 22430 37378 22482
rect 5854 22318 5906 22370
rect 6302 22318 6354 22370
rect 6750 22318 6802 22370
rect 6974 22318 7026 22370
rect 7422 22318 7474 22370
rect 7982 22318 8034 22370
rect 9886 22318 9938 22370
rect 10334 22318 10386 22370
rect 13470 22318 13522 22370
rect 13694 22318 13746 22370
rect 14254 22318 14306 22370
rect 15150 22318 15202 22370
rect 15710 22318 15762 22370
rect 16046 22318 16098 22370
rect 17950 22318 18002 22370
rect 18286 22318 18338 22370
rect 18958 22318 19010 22370
rect 20078 22318 20130 22370
rect 29262 22318 29314 22370
rect 29934 22318 29986 22370
rect 30046 22318 30098 22370
rect 32174 22318 32226 22370
rect 32846 22318 32898 22370
rect 36430 22318 36482 22370
rect 37438 22318 37490 22370
rect 5966 22206 6018 22258
rect 8878 22206 8930 22258
rect 9998 22206 10050 22258
rect 10110 22206 10162 22258
rect 10782 22206 10834 22258
rect 14590 22206 14642 22258
rect 15486 22206 15538 22258
rect 15598 22206 15650 22258
rect 19070 22206 19122 22258
rect 19854 22206 19906 22258
rect 20414 22206 20466 22258
rect 29374 22206 29426 22258
rect 31950 22206 32002 22258
rect 32510 22206 32562 22258
rect 33630 22206 33682 22258
rect 36094 22206 36146 22258
rect 6190 22094 6242 22146
rect 6862 22094 6914 22146
rect 7310 22094 7362 22146
rect 8542 22094 8594 22146
rect 13918 22094 13970 22146
rect 16606 22094 16658 22146
rect 17838 22094 17890 22146
rect 18174 22094 18226 22146
rect 18958 22094 19010 22146
rect 20750 22094 20802 22146
rect 28254 22094 28306 22146
rect 29822 22094 29874 22146
rect 30942 22094 30994 22146
rect 31502 22094 31554 22146
rect 31726 22094 31778 22146
rect 31838 22094 31890 22146
rect 32398 22094 32450 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 8430 21758 8482 21810
rect 14702 21758 14754 21810
rect 18734 21758 18786 21810
rect 25342 21758 25394 21810
rect 32622 21758 32674 21810
rect 7758 21646 7810 21698
rect 8654 21646 8706 21698
rect 9550 21646 9602 21698
rect 9774 21646 9826 21698
rect 14366 21646 14418 21698
rect 26686 21646 26738 21698
rect 27806 21646 27858 21698
rect 31838 21646 31890 21698
rect 33182 21646 33234 21698
rect 3726 21534 3778 21586
rect 5070 21534 5122 21586
rect 6414 21534 6466 21586
rect 6974 21534 7026 21586
rect 7534 21534 7586 21586
rect 8206 21534 8258 21586
rect 8878 21534 8930 21586
rect 13470 21534 13522 21586
rect 13806 21534 13858 21586
rect 14590 21534 14642 21586
rect 14926 21534 14978 21586
rect 15150 21534 15202 21586
rect 18510 21534 18562 21586
rect 18846 21534 18898 21586
rect 19070 21534 19122 21586
rect 19406 21534 19458 21586
rect 25902 21534 25954 21586
rect 26350 21534 26402 21586
rect 27022 21534 27074 21586
rect 31166 21534 31218 21586
rect 36654 21534 36706 21586
rect 3054 21422 3106 21474
rect 3950 21422 4002 21474
rect 5406 21422 5458 21474
rect 7870 21422 7922 21474
rect 9886 21422 9938 21474
rect 13918 21422 13970 21474
rect 15598 21422 15650 21474
rect 22990 21422 23042 21474
rect 29934 21422 29986 21474
rect 30494 21422 30546 21474
rect 31390 21422 31442 21474
rect 34302 21422 34354 21474
rect 36430 21422 36482 21474
rect 37438 21422 37490 21474
rect 39566 21422 39618 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 9550 20974 9602 21026
rect 11566 20974 11618 21026
rect 18846 20974 18898 21026
rect 19406 20974 19458 21026
rect 19630 20974 19682 21026
rect 19966 20974 20018 21026
rect 37438 20974 37490 21026
rect 4622 20862 4674 20914
rect 7422 20862 7474 20914
rect 7646 20862 7698 20914
rect 18846 20862 18898 20914
rect 25678 20862 25730 20914
rect 31838 20862 31890 20914
rect 32286 20862 32338 20914
rect 33070 20862 33122 20914
rect 37550 20862 37602 20914
rect 1822 20750 1874 20802
rect 7870 20750 7922 20802
rect 8654 20750 8706 20802
rect 10446 20750 10498 20802
rect 19742 20750 19794 20802
rect 20078 20750 20130 20802
rect 22878 20750 22930 20802
rect 26350 20750 26402 20802
rect 26798 20750 26850 20802
rect 27246 20750 27298 20802
rect 27694 20750 27746 20802
rect 31614 20750 31666 20802
rect 33406 20750 33458 20802
rect 37774 20750 37826 20802
rect 2494 20638 2546 20690
rect 8318 20638 8370 20690
rect 9662 20638 9714 20690
rect 10110 20638 10162 20690
rect 11678 20638 11730 20690
rect 15038 20638 15090 20690
rect 21646 20638 21698 20690
rect 23550 20638 23602 20690
rect 26014 20638 26066 20690
rect 27582 20638 27634 20690
rect 28254 20638 28306 20690
rect 5070 20526 5122 20578
rect 7086 20526 7138 20578
rect 11230 20526 11282 20578
rect 11566 20526 11618 20578
rect 14702 20526 14754 20578
rect 19294 20526 19346 20578
rect 21310 20526 21362 20578
rect 27470 20526 27522 20578
rect 30494 20526 30546 20578
rect 33742 20526 33794 20578
rect 37102 20526 37154 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 5854 20190 5906 20242
rect 8654 20190 8706 20242
rect 14142 20190 14194 20242
rect 2942 20078 2994 20130
rect 3166 20078 3218 20130
rect 6414 20078 6466 20130
rect 9550 20078 9602 20130
rect 10782 20078 10834 20130
rect 12686 20078 12738 20130
rect 15150 20078 15202 20130
rect 15486 20078 15538 20130
rect 16382 20078 16434 20130
rect 16718 20078 16770 20130
rect 17390 20078 17442 20130
rect 20526 20078 20578 20130
rect 21534 20078 21586 20130
rect 26910 20078 26962 20130
rect 27022 20078 27074 20130
rect 28030 20078 28082 20130
rect 35982 20078 36034 20130
rect 6302 19966 6354 20018
rect 6526 19966 6578 20018
rect 8430 19966 8482 20018
rect 9774 19966 9826 20018
rect 12238 19966 12290 20018
rect 12798 19966 12850 20018
rect 13358 19966 13410 20018
rect 14478 19966 14530 20018
rect 14814 19966 14866 20018
rect 15934 19966 15986 20018
rect 18958 19966 19010 20018
rect 19406 19966 19458 20018
rect 19742 19966 19794 20018
rect 19966 19966 20018 20018
rect 20078 19966 20130 20018
rect 22094 19966 22146 20018
rect 23102 19966 23154 20018
rect 23774 19966 23826 20018
rect 24222 19966 24274 20018
rect 24446 19966 24498 20018
rect 25902 19966 25954 20018
rect 26126 19966 26178 20018
rect 26350 19966 26402 20018
rect 26686 19966 26738 20018
rect 28590 19966 28642 20018
rect 35758 19966 35810 20018
rect 2830 19854 2882 19906
rect 4286 19854 4338 19906
rect 12462 19854 12514 19906
rect 13806 19854 13858 19906
rect 17838 19854 17890 19906
rect 21198 19854 21250 19906
rect 21646 19854 21698 19906
rect 21870 19854 21922 19906
rect 22654 19854 22706 19906
rect 23998 19854 24050 19906
rect 28142 19854 28194 19906
rect 9998 19742 10050 19794
rect 10222 19742 10274 19794
rect 23214 19742 23266 19794
rect 25454 19742 25506 19794
rect 27470 19742 27522 19794
rect 27806 19742 27858 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 3838 19406 3890 19458
rect 5630 19406 5682 19458
rect 13694 19406 13746 19458
rect 22094 19406 22146 19458
rect 23214 19406 23266 19458
rect 26350 19406 26402 19458
rect 31166 19406 31218 19458
rect 31502 19406 31554 19458
rect 33406 19406 33458 19458
rect 14590 19294 14642 19346
rect 15934 19294 15986 19346
rect 20638 19294 20690 19346
rect 23438 19294 23490 19346
rect 26798 19294 26850 19346
rect 37550 19294 37602 19346
rect 3614 19182 3666 19234
rect 4062 19182 4114 19234
rect 5070 19182 5122 19234
rect 5966 19182 6018 19234
rect 6190 19182 6242 19234
rect 9102 19182 9154 19234
rect 11118 19182 11170 19234
rect 13470 19182 13522 19234
rect 14254 19182 14306 19234
rect 17054 19182 17106 19234
rect 21310 19182 21362 19234
rect 23550 19182 23602 19234
rect 27022 19182 27074 19234
rect 27246 19182 27298 19234
rect 31726 19182 31778 19234
rect 32062 19182 32114 19234
rect 32174 19182 32226 19234
rect 32510 19182 32562 19234
rect 33406 19182 33458 19234
rect 37326 19182 37378 19234
rect 3502 19070 3554 19122
rect 4734 19070 4786 19122
rect 9214 19070 9266 19122
rect 12910 19070 12962 19122
rect 14814 19070 14866 19122
rect 19630 19070 19682 19122
rect 21534 19070 21586 19122
rect 21646 19070 21698 19122
rect 22766 19070 22818 19122
rect 23102 19070 23154 19122
rect 33742 19070 33794 19122
rect 36206 19070 36258 19122
rect 36318 19070 36370 19122
rect 12798 18958 12850 19010
rect 14030 18958 14082 19010
rect 14590 18958 14642 19010
rect 15150 18958 15202 19010
rect 15486 18958 15538 19010
rect 17390 18958 17442 19010
rect 19294 18958 19346 19010
rect 20190 18958 20242 19010
rect 27694 18958 27746 19010
rect 36542 18958 36594 19010
rect 36990 18958 37042 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 4286 18622 4338 18674
rect 14590 18622 14642 18674
rect 18286 18622 18338 18674
rect 19742 18622 19794 18674
rect 31950 18622 32002 18674
rect 33070 18622 33122 18674
rect 38334 18622 38386 18674
rect 19854 18510 19906 18562
rect 26462 18510 26514 18562
rect 31726 18510 31778 18562
rect 35758 18510 35810 18562
rect 36094 18510 36146 18562
rect 38110 18510 38162 18562
rect 4510 18398 4562 18450
rect 13694 18398 13746 18450
rect 18398 18398 18450 18450
rect 18846 18398 18898 18450
rect 26126 18398 26178 18450
rect 32286 18398 32338 18450
rect 33742 18398 33794 18450
rect 35870 18398 35922 18450
rect 36318 18398 36370 18450
rect 37102 18398 37154 18450
rect 38222 18398 38274 18450
rect 13918 18286 13970 18338
rect 14702 18286 14754 18338
rect 33966 18286 34018 18338
rect 34414 18286 34466 18338
rect 35982 18286 36034 18338
rect 37550 18286 37602 18338
rect 4174 18174 4226 18226
rect 14142 18174 14194 18226
rect 18286 18174 18338 18226
rect 19742 18174 19794 18226
rect 31614 18174 31666 18226
rect 33182 18174 33234 18226
rect 33406 18174 33458 18226
rect 37214 18174 37266 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 20190 17838 20242 17890
rect 23438 17838 23490 17890
rect 31278 17838 31330 17890
rect 31614 17838 31666 17890
rect 2494 17726 2546 17778
rect 4622 17726 4674 17778
rect 5070 17726 5122 17778
rect 19070 17726 19122 17778
rect 25118 17726 25170 17778
rect 34750 17726 34802 17778
rect 37102 17726 37154 17778
rect 1822 17614 1874 17666
rect 5742 17614 5794 17666
rect 8766 17614 8818 17666
rect 15822 17614 15874 17666
rect 16158 17614 16210 17666
rect 19630 17614 19682 17666
rect 19742 17614 19794 17666
rect 22542 17614 22594 17666
rect 23214 17614 23266 17666
rect 23774 17614 23826 17666
rect 36990 17614 37042 17666
rect 37214 17614 37266 17666
rect 5966 17502 6018 17554
rect 8430 17502 8482 17554
rect 8542 17502 8594 17554
rect 16942 17502 16994 17554
rect 19518 17502 19570 17554
rect 22878 17502 22930 17554
rect 23998 17502 24050 17554
rect 24334 17502 24386 17554
rect 24558 17502 24610 17554
rect 32622 17502 32674 17554
rect 37438 17502 37490 17554
rect 37886 17502 37938 17554
rect 37998 17502 38050 17554
rect 23662 17390 23714 17442
rect 24446 17390 24498 17442
rect 31614 17390 31666 17442
rect 37662 17390 37714 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 11678 17054 11730 17106
rect 17614 17054 17666 17106
rect 18846 17054 18898 17106
rect 22878 17054 22930 17106
rect 23438 17054 23490 17106
rect 29934 17054 29986 17106
rect 30494 17054 30546 17106
rect 32062 17054 32114 17106
rect 36654 17054 36706 17106
rect 7310 16942 7362 16994
rect 7646 16942 7698 16994
rect 10558 16942 10610 16994
rect 11118 16942 11170 16994
rect 18398 16942 18450 16994
rect 23214 16942 23266 16994
rect 23550 16942 23602 16994
rect 24558 16942 24610 16994
rect 25230 16942 25282 16994
rect 27470 16942 27522 16994
rect 30046 16942 30098 16994
rect 30942 16942 30994 16994
rect 31614 16942 31666 16994
rect 35310 16942 35362 16994
rect 10110 16830 10162 16882
rect 10446 16830 10498 16882
rect 17838 16830 17890 16882
rect 17950 16830 18002 16882
rect 18174 16830 18226 16882
rect 23662 16830 23714 16882
rect 24110 16830 24162 16882
rect 24334 16830 24386 16882
rect 25566 16830 25618 16882
rect 26798 16830 26850 16882
rect 31390 16830 31442 16882
rect 32174 16830 32226 16882
rect 32958 16830 33010 16882
rect 11230 16718 11282 16770
rect 19294 16718 19346 16770
rect 29598 16718 29650 16770
rect 37214 16718 37266 16770
rect 10894 16606 10946 16658
rect 24222 16606 24274 16658
rect 32062 16606 32114 16658
rect 36990 16606 37042 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 6078 16270 6130 16322
rect 6302 16270 6354 16322
rect 7758 16270 7810 16322
rect 22654 16270 22706 16322
rect 30046 16270 30098 16322
rect 3502 16158 3554 16210
rect 9886 16158 9938 16210
rect 10446 16158 10498 16210
rect 12574 16158 12626 16210
rect 15710 16158 15762 16210
rect 18174 16158 18226 16210
rect 18734 16158 18786 16210
rect 19854 16158 19906 16210
rect 31614 16158 31666 16210
rect 33742 16158 33794 16210
rect 36990 16158 37042 16210
rect 4286 16046 4338 16098
rect 5854 16046 5906 16098
rect 6750 16046 6802 16098
rect 7086 16046 7138 16098
rect 9214 16046 9266 16098
rect 9774 16046 9826 16098
rect 23214 16046 23266 16098
rect 24446 16046 24498 16098
rect 25566 16046 25618 16098
rect 26686 16046 26738 16098
rect 27022 16046 27074 16098
rect 28590 16046 28642 16098
rect 30494 16046 30546 16098
rect 34414 16046 34466 16098
rect 35534 16046 35586 16098
rect 37438 16046 37490 16098
rect 37886 16046 37938 16098
rect 38558 16046 38610 16098
rect 3950 15934 4002 15986
rect 5630 15934 5682 15986
rect 7646 15934 7698 15986
rect 13918 15934 13970 15986
rect 14142 15934 14194 15986
rect 14366 15934 14418 15986
rect 14590 15934 14642 15986
rect 18622 15934 18674 15986
rect 18846 15934 18898 15986
rect 19294 15934 19346 15986
rect 19406 15934 19458 15986
rect 22430 15934 22482 15986
rect 23102 15934 23154 15986
rect 23326 15934 23378 15986
rect 23886 15934 23938 15986
rect 25454 15934 25506 15986
rect 27246 15934 27298 15986
rect 27806 15934 27858 15986
rect 29934 15934 29986 15986
rect 34862 15934 34914 15986
rect 35198 15934 35250 15986
rect 35870 15934 35922 15986
rect 38334 15934 38386 15986
rect 4062 15822 4114 15874
rect 7422 15822 7474 15874
rect 14478 15822 14530 15874
rect 14926 15822 14978 15874
rect 15262 15822 15314 15874
rect 19070 15822 19122 15874
rect 23998 15822 24050 15874
rect 27358 15822 27410 15874
rect 28030 15822 28082 15874
rect 30046 15822 30098 15874
rect 31054 15822 31106 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 3614 15486 3666 15538
rect 6078 15486 6130 15538
rect 7758 15486 7810 15538
rect 16046 15486 16098 15538
rect 17726 15486 17778 15538
rect 17838 15486 17890 15538
rect 19742 15486 19794 15538
rect 20078 15486 20130 15538
rect 20750 15486 20802 15538
rect 23102 15486 23154 15538
rect 23438 15486 23490 15538
rect 24334 15486 24386 15538
rect 30606 15486 30658 15538
rect 31278 15486 31330 15538
rect 32062 15486 32114 15538
rect 36318 15486 36370 15538
rect 4846 15374 4898 15426
rect 5070 15374 5122 15426
rect 5630 15374 5682 15426
rect 6302 15374 6354 15426
rect 7198 15374 7250 15426
rect 8990 15374 9042 15426
rect 10334 15374 10386 15426
rect 12014 15374 12066 15426
rect 14814 15374 14866 15426
rect 19854 15374 19906 15426
rect 29598 15374 29650 15426
rect 35310 15374 35362 15426
rect 2830 15262 2882 15314
rect 3054 15262 3106 15314
rect 3278 15262 3330 15314
rect 4062 15262 4114 15314
rect 4174 15262 4226 15314
rect 4398 15262 4450 15314
rect 4622 15262 4674 15314
rect 5294 15262 5346 15314
rect 5854 15262 5906 15314
rect 6862 15262 6914 15314
rect 6974 15262 7026 15314
rect 7310 15262 7362 15314
rect 8542 15262 8594 15314
rect 11566 15262 11618 15314
rect 15598 15262 15650 15314
rect 17614 15262 17666 15314
rect 17950 15262 18002 15314
rect 18174 15262 18226 15314
rect 19070 15262 19122 15314
rect 19294 15262 19346 15314
rect 20302 15262 20354 15314
rect 29822 15262 29874 15314
rect 31950 15262 32002 15314
rect 32174 15262 32226 15314
rect 32622 15262 32674 15314
rect 32958 15262 33010 15314
rect 36654 15262 36706 15314
rect 8094 15150 8146 15202
rect 10110 15150 10162 15202
rect 12686 15150 12738 15202
rect 18398 15150 18450 15202
rect 19518 15150 19570 15202
rect 23774 15150 23826 15202
rect 37438 15150 37490 15202
rect 39566 15150 39618 15202
rect 2718 15038 2770 15090
rect 6190 15038 6242 15090
rect 18846 15038 18898 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 3502 14702 3554 14754
rect 3726 14702 3778 14754
rect 18622 14702 18674 14754
rect 23886 14702 23938 14754
rect 4510 14590 4562 14642
rect 11566 14590 11618 14642
rect 19854 14590 19906 14642
rect 29598 14590 29650 14642
rect 30494 14590 30546 14642
rect 30942 14590 30994 14642
rect 31726 14590 31778 14642
rect 3950 14478 4002 14530
rect 4958 14478 5010 14530
rect 6750 14478 6802 14530
rect 12126 14478 12178 14530
rect 12462 14478 12514 14530
rect 12574 14478 12626 14530
rect 15150 14478 15202 14530
rect 18734 14478 18786 14530
rect 18958 14478 19010 14530
rect 19182 14478 19234 14530
rect 19518 14478 19570 14530
rect 19966 14478 20018 14530
rect 20190 14478 20242 14530
rect 22542 14478 22594 14530
rect 29934 14478 29986 14530
rect 3390 14366 3442 14418
rect 4734 14366 4786 14418
rect 5854 14366 5906 14418
rect 6190 14366 6242 14418
rect 6526 14366 6578 14418
rect 13582 14366 13634 14418
rect 23774 14366 23826 14418
rect 29486 14366 29538 14418
rect 29710 14366 29762 14418
rect 30606 14366 30658 14418
rect 31166 14366 31218 14418
rect 37326 14366 37378 14418
rect 11454 14254 11506 14306
rect 11678 14254 11730 14306
rect 12350 14254 12402 14306
rect 12798 14254 12850 14306
rect 13470 14254 13522 14306
rect 14590 14254 14642 14306
rect 17614 14254 17666 14306
rect 17950 14254 18002 14306
rect 18286 14254 18338 14306
rect 19742 14254 19794 14306
rect 22878 14254 22930 14306
rect 26014 14254 26066 14306
rect 28590 14254 28642 14306
rect 30382 14254 30434 14306
rect 31054 14254 31106 14306
rect 39678 14254 39730 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 9662 13918 9714 13970
rect 16270 13918 16322 13970
rect 17614 13918 17666 13970
rect 18174 13918 18226 13970
rect 18398 13918 18450 13970
rect 19966 13918 20018 13970
rect 26126 13918 26178 13970
rect 33182 13918 33234 13970
rect 37102 13918 37154 13970
rect 37214 13918 37266 13970
rect 37326 13918 37378 13970
rect 2606 13806 2658 13858
rect 19182 13806 19234 13858
rect 19406 13806 19458 13858
rect 25342 13806 25394 13858
rect 25902 13806 25954 13858
rect 31278 13806 31330 13858
rect 35870 13806 35922 13858
rect 37438 13806 37490 13858
rect 37662 13806 37714 13858
rect 38110 13806 38162 13858
rect 38334 13806 38386 13858
rect 38558 13806 38610 13858
rect 38782 13806 38834 13858
rect 1934 13694 1986 13746
rect 12014 13694 12066 13746
rect 17950 13694 18002 13746
rect 18510 13694 18562 13746
rect 25790 13694 25842 13746
rect 26350 13694 26402 13746
rect 38894 13694 38946 13746
rect 4734 13582 4786 13634
rect 5182 13582 5234 13634
rect 9550 13582 9602 13634
rect 15038 13582 15090 13634
rect 22654 13582 22706 13634
rect 37998 13582 38050 13634
rect 39342 13582 39394 13634
rect 19070 13470 19122 13522
rect 22766 13470 22818 13522
rect 25454 13470 25506 13522
rect 33742 13470 33794 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19742 13134 19794 13186
rect 38446 13134 38498 13186
rect 7198 13022 7250 13074
rect 10670 13022 10722 13074
rect 18734 13022 18786 13074
rect 23438 13022 23490 13074
rect 24894 13022 24946 13074
rect 29262 13022 29314 13074
rect 33182 13022 33234 13074
rect 34414 13022 34466 13074
rect 36430 13022 36482 13074
rect 37662 13022 37714 13074
rect 8094 12910 8146 12962
rect 19070 12910 19122 12962
rect 22318 12910 22370 12962
rect 22766 12910 22818 12962
rect 23886 12910 23938 12962
rect 25230 12910 25282 12962
rect 26014 12910 26066 12962
rect 26238 12910 26290 12962
rect 27134 12910 27186 12962
rect 27694 12910 27746 12962
rect 28142 12910 28194 12962
rect 29486 12910 29538 12962
rect 29934 12910 29986 12962
rect 30942 12910 30994 12962
rect 31390 12910 31442 12962
rect 32398 12910 32450 12962
rect 32622 12910 32674 12962
rect 33294 12910 33346 12962
rect 33630 12910 33682 12962
rect 34190 12910 34242 12962
rect 34862 12910 34914 12962
rect 37214 12910 37266 12962
rect 8206 12798 8258 12850
rect 11118 12798 11170 12850
rect 12574 12798 12626 12850
rect 19294 12798 19346 12850
rect 19630 12798 19682 12850
rect 22990 12798 23042 12850
rect 25678 12798 25730 12850
rect 27470 12798 27522 12850
rect 28478 12798 28530 12850
rect 30046 12798 30098 12850
rect 30718 12798 30770 12850
rect 31614 12798 31666 12850
rect 31950 12798 32002 12850
rect 32174 12798 32226 12850
rect 33966 12798 34018 12850
rect 34526 12798 34578 12850
rect 37774 12798 37826 12850
rect 37998 12798 38050 12850
rect 38334 12798 38386 12850
rect 38446 12798 38498 12850
rect 7310 12686 7362 12738
rect 8430 12686 8482 12738
rect 12462 12686 12514 12738
rect 18734 12686 18786 12738
rect 18846 12686 18898 12738
rect 19742 12686 19794 12738
rect 30158 12686 30210 12738
rect 31166 12686 31218 12738
rect 31726 12686 31778 12738
rect 32398 12686 32450 12738
rect 33070 12686 33122 12738
rect 34974 12686 35026 12738
rect 35198 12686 35250 12738
rect 36990 12686 37042 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 5630 12350 5682 12402
rect 6638 12350 6690 12402
rect 8094 12350 8146 12402
rect 8766 12350 8818 12402
rect 18286 12350 18338 12402
rect 19294 12350 19346 12402
rect 19406 12350 19458 12402
rect 21422 12350 21474 12402
rect 25790 12350 25842 12402
rect 30270 12350 30322 12402
rect 33406 12350 33458 12402
rect 33630 12350 33682 12402
rect 33742 12350 33794 12402
rect 34862 12350 34914 12402
rect 37102 12350 37154 12402
rect 3054 12238 3106 12290
rect 12462 12238 12514 12290
rect 17950 12238 18002 12290
rect 25342 12238 25394 12290
rect 25566 12238 25618 12290
rect 26238 12238 26290 12290
rect 26574 12238 26626 12290
rect 29150 12238 29202 12290
rect 34078 12238 34130 12290
rect 35870 12238 35922 12290
rect 37214 12238 37266 12290
rect 37550 12238 37602 12290
rect 2270 12126 2322 12178
rect 6302 12126 6354 12178
rect 7758 12126 7810 12178
rect 8094 12126 8146 12178
rect 8318 12126 8370 12178
rect 8542 12126 8594 12178
rect 8878 12126 8930 12178
rect 9998 12126 10050 12178
rect 10446 12126 10498 12178
rect 17614 12126 17666 12178
rect 18286 12126 18338 12178
rect 18622 12126 18674 12178
rect 18846 12126 18898 12178
rect 19070 12126 19122 12178
rect 19630 12126 19682 12178
rect 19966 12126 20018 12178
rect 21758 12126 21810 12178
rect 22206 12126 22258 12178
rect 25790 12126 25842 12178
rect 26014 12126 26066 12178
rect 28142 12126 28194 12178
rect 28590 12126 28642 12178
rect 33182 12126 33234 12178
rect 35086 12126 35138 12178
rect 36206 12126 36258 12178
rect 36990 12126 37042 12178
rect 37438 12126 37490 12178
rect 5182 12014 5234 12066
rect 5406 12014 5458 12066
rect 9550 12014 9602 12066
rect 12574 12014 12626 12066
rect 17838 12014 17890 12066
rect 24782 12014 24834 12066
rect 33966 12014 34018 12066
rect 5854 11902 5906 11954
rect 6078 11902 6130 11954
rect 7310 11902 7362 11954
rect 7646 11902 7698 11954
rect 12238 11902 12290 11954
rect 34302 11902 34354 11954
rect 36206 11902 36258 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 6414 11566 6466 11618
rect 7422 11566 7474 11618
rect 18846 11566 18898 11618
rect 22206 11566 22258 11618
rect 28254 11566 28306 11618
rect 37886 11566 37938 11618
rect 7310 11454 7362 11506
rect 13694 11454 13746 11506
rect 15822 11454 15874 11506
rect 22430 11454 22482 11506
rect 29262 11454 29314 11506
rect 32622 11454 32674 11506
rect 36430 11454 36482 11506
rect 37102 11454 37154 11506
rect 5854 11342 5906 11394
rect 6750 11342 6802 11394
rect 8654 11342 8706 11394
rect 9550 11342 9602 11394
rect 11454 11342 11506 11394
rect 11790 11342 11842 11394
rect 12014 11342 12066 11394
rect 12574 11342 12626 11394
rect 16606 11342 16658 11394
rect 17726 11342 17778 11394
rect 18622 11342 18674 11394
rect 19070 11342 19122 11394
rect 19406 11342 19458 11394
rect 19630 11342 19682 11394
rect 19966 11342 20018 11394
rect 20750 11342 20802 11394
rect 21870 11342 21922 11394
rect 23214 11342 23266 11394
rect 25790 11342 25842 11394
rect 26686 11342 26738 11394
rect 27470 11342 27522 11394
rect 5966 11230 6018 11282
rect 8094 11230 8146 11282
rect 11566 11230 11618 11282
rect 17950 11230 18002 11282
rect 21646 11230 21698 11282
rect 22766 11230 22818 11282
rect 22878 11230 22930 11282
rect 22990 11230 23042 11282
rect 23662 11230 23714 11282
rect 26574 11230 26626 11282
rect 27358 11230 27410 11282
rect 28366 11230 28418 11282
rect 31726 11230 31778 11282
rect 32286 11230 32338 11282
rect 35534 11230 35586 11282
rect 38110 11230 38162 11282
rect 38558 11230 38610 11282
rect 38670 11230 38722 11282
rect 6190 11118 6242 11170
rect 6526 11118 6578 11170
rect 7198 11118 7250 11170
rect 9662 11118 9714 11170
rect 12350 11118 12402 11170
rect 12462 11118 12514 11170
rect 17054 11118 17106 11170
rect 17838 11118 17890 11170
rect 18174 11118 18226 11170
rect 18958 11118 19010 11170
rect 19854 11118 19906 11170
rect 22094 11118 22146 11170
rect 25230 11118 25282 11170
rect 31838 11118 31890 11170
rect 32062 11118 32114 11170
rect 32510 11118 32562 11170
rect 35870 11118 35922 11170
rect 36990 11118 37042 11170
rect 37214 11118 37266 11170
rect 37438 11118 37490 11170
rect 37998 11118 38050 11170
rect 38894 11118 38946 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 7086 10782 7138 10834
rect 7310 10782 7362 10834
rect 8206 10782 8258 10834
rect 18846 10782 18898 10834
rect 19070 10782 19122 10834
rect 19742 10782 19794 10834
rect 20190 10782 20242 10834
rect 29262 10782 29314 10834
rect 35422 10782 35474 10834
rect 37438 10782 37490 10834
rect 37662 10782 37714 10834
rect 38670 10782 38722 10834
rect 7870 10670 7922 10722
rect 7982 10670 8034 10722
rect 16606 10670 16658 10722
rect 17950 10670 18002 10722
rect 18622 10670 18674 10722
rect 28030 10670 28082 10722
rect 30158 10670 30210 10722
rect 33518 10670 33570 10722
rect 38782 10670 38834 10722
rect 7534 10558 7586 10610
rect 13022 10558 13074 10610
rect 17726 10558 17778 10610
rect 18398 10558 18450 10610
rect 21198 10558 21250 10610
rect 24558 10558 24610 10610
rect 26574 10558 26626 10610
rect 27022 10558 27074 10610
rect 27694 10558 27746 10610
rect 28590 10558 28642 10610
rect 29038 10558 29090 10610
rect 29598 10558 29650 10610
rect 29822 10558 29874 10610
rect 31950 10558 32002 10610
rect 32510 10558 32562 10610
rect 33070 10558 33122 10610
rect 33294 10558 33346 10610
rect 33742 10558 33794 10610
rect 34862 10558 34914 10610
rect 35310 10558 35362 10610
rect 35534 10558 35586 10610
rect 36318 10558 36370 10610
rect 36542 10558 36594 10610
rect 37886 10558 37938 10610
rect 38110 10558 38162 10610
rect 38558 10558 38610 10610
rect 39118 10558 39170 10610
rect 7422 10446 7474 10498
rect 18174 10446 18226 10498
rect 21870 10446 21922 10498
rect 23998 10446 24050 10498
rect 28142 10446 28194 10498
rect 29150 10446 29202 10498
rect 30046 10446 30098 10498
rect 33630 10446 33682 10498
rect 35982 10446 36034 10498
rect 38222 10446 38274 10498
rect 18734 10334 18786 10386
rect 32174 10334 32226 10386
rect 36990 10334 37042 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 2830 9998 2882 10050
rect 22318 9998 22370 10050
rect 30494 9998 30546 10050
rect 31726 9998 31778 10050
rect 33518 9998 33570 10050
rect 22430 9886 22482 9938
rect 23102 9886 23154 9938
rect 23998 9886 24050 9938
rect 26350 9886 26402 9938
rect 29486 9886 29538 9938
rect 32734 9886 32786 9938
rect 3166 9774 3218 9826
rect 8542 9774 8594 9826
rect 9550 9774 9602 9826
rect 13582 9774 13634 9826
rect 14142 9774 14194 9826
rect 14254 9774 14306 9826
rect 14702 9774 14754 9826
rect 23550 9774 23602 9826
rect 26574 9774 26626 9826
rect 27022 9774 27074 9826
rect 27582 9774 27634 9826
rect 28254 9774 28306 9826
rect 29150 9774 29202 9826
rect 29598 9774 29650 9826
rect 29822 9774 29874 9826
rect 30718 9774 30770 9826
rect 31278 9774 31330 9826
rect 31838 9774 31890 9826
rect 32398 9774 32450 9826
rect 36990 9774 37042 9826
rect 37550 9774 37602 9826
rect 39230 9774 39282 9826
rect 4062 9662 4114 9714
rect 8318 9662 8370 9714
rect 9998 9662 10050 9714
rect 13918 9662 13970 9714
rect 15038 9662 15090 9714
rect 18062 9662 18114 9714
rect 18398 9662 18450 9714
rect 19070 9662 19122 9714
rect 27246 9662 27298 9714
rect 27918 9662 27970 9714
rect 28590 9662 28642 9714
rect 32174 9662 32226 9714
rect 32622 9662 32674 9714
rect 35646 9662 35698 9714
rect 37998 9662 38050 9714
rect 39118 9662 39170 9714
rect 2942 9550 2994 9602
rect 4398 9550 4450 9602
rect 13358 9550 13410 9602
rect 16942 9550 16994 9602
rect 17390 9550 17442 9602
rect 18734 9550 18786 9602
rect 26798 9550 26850 9602
rect 29374 9550 29426 9602
rect 30158 9550 30210 9602
rect 31726 9550 31778 9602
rect 32734 9550 32786 9602
rect 33294 9550 33346 9602
rect 37214 9550 37266 9602
rect 37326 9550 37378 9602
rect 37438 9550 37490 9602
rect 38334 9550 38386 9602
rect 38894 9550 38946 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 9662 9214 9714 9266
rect 33630 9214 33682 9266
rect 34302 9214 34354 9266
rect 34526 9214 34578 9266
rect 35758 9214 35810 9266
rect 36318 9214 36370 9266
rect 39006 9214 39058 9266
rect 2494 9102 2546 9154
rect 12238 9102 12290 9154
rect 13918 9102 13970 9154
rect 28702 9102 28754 9154
rect 31166 9102 31218 9154
rect 34078 9102 34130 9154
rect 36990 9102 37042 9154
rect 37326 9102 37378 9154
rect 37662 9102 37714 9154
rect 37998 9102 38050 9154
rect 38334 9102 38386 9154
rect 1822 8990 1874 9042
rect 9438 8990 9490 9042
rect 9886 8990 9938 9042
rect 10110 8990 10162 9042
rect 13246 8990 13298 9042
rect 24670 8990 24722 9042
rect 25342 8990 25394 9042
rect 31278 8990 31330 9042
rect 33070 8990 33122 9042
rect 33518 8990 33570 9042
rect 33742 8990 33794 9042
rect 34638 8990 34690 9042
rect 35870 8990 35922 9042
rect 36206 8990 36258 9042
rect 38558 8990 38610 9042
rect 39230 8990 39282 9042
rect 4622 8878 4674 8930
rect 5070 8878 5122 8930
rect 11790 8878 11842 8930
rect 31726 8878 31778 8930
rect 31166 8766 31218 8818
rect 31614 8766 31666 8818
rect 36318 8766 36370 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 13582 8430 13634 8482
rect 34078 8430 34130 8482
rect 3950 8318 4002 8370
rect 12462 8318 12514 8370
rect 16046 8318 16098 8370
rect 16494 8318 16546 8370
rect 18622 8318 18674 8370
rect 19854 8318 19906 8370
rect 29598 8318 29650 8370
rect 30158 8318 30210 8370
rect 31838 8318 31890 8370
rect 37998 8318 38050 8370
rect 2382 8206 2434 8258
rect 3726 8206 3778 8258
rect 12238 8206 12290 8258
rect 12686 8206 12738 8258
rect 13918 8206 13970 8258
rect 15262 8206 15314 8258
rect 15934 8206 15986 8258
rect 19406 8206 19458 8258
rect 26238 8206 26290 8258
rect 29486 8206 29538 8258
rect 29934 8206 29986 8258
rect 30494 8206 30546 8258
rect 31614 8206 31666 8258
rect 32622 8206 32674 8258
rect 33182 8206 33234 8258
rect 33406 8206 33458 8258
rect 33630 8206 33682 8258
rect 34526 8206 34578 8258
rect 36542 8206 36594 8258
rect 37326 8206 37378 8258
rect 37774 8206 37826 8258
rect 38110 8206 38162 8258
rect 38894 8206 38946 8258
rect 2718 8094 2770 8146
rect 3054 8094 3106 8146
rect 5070 8094 5122 8146
rect 5630 8094 5682 8146
rect 5966 8094 6018 8146
rect 8878 8094 8930 8146
rect 12910 8094 12962 8146
rect 14142 8094 14194 8146
rect 14702 8094 14754 8146
rect 15150 8094 15202 8146
rect 15374 8094 15426 8146
rect 29710 8094 29762 8146
rect 31950 8094 32002 8146
rect 32286 8094 32338 8146
rect 32398 8094 32450 8146
rect 34302 8094 34354 8146
rect 36206 8094 36258 8146
rect 36318 8094 36370 8146
rect 36990 8094 37042 8146
rect 37550 8094 37602 8146
rect 39006 8094 39058 8146
rect 2606 7982 2658 8034
rect 4958 7982 5010 8034
rect 8990 7982 9042 8034
rect 26574 7982 26626 8034
rect 30718 7982 30770 8034
rect 30830 7982 30882 8034
rect 30942 7982 30994 8034
rect 31054 7982 31106 8034
rect 37102 7982 37154 8034
rect 38558 7982 38610 8034
rect 39230 7982 39282 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 6638 7646 6690 7698
rect 9662 7646 9714 7698
rect 9886 7646 9938 7698
rect 10558 7646 10610 7698
rect 15822 7646 15874 7698
rect 17726 7646 17778 7698
rect 20750 7646 20802 7698
rect 21422 7646 21474 7698
rect 28590 7646 28642 7698
rect 29598 7646 29650 7698
rect 32174 7646 32226 7698
rect 32398 7646 32450 7698
rect 2718 7534 2770 7586
rect 8094 7534 8146 7586
rect 9774 7534 9826 7586
rect 10670 7534 10722 7586
rect 14478 7534 14530 7586
rect 21758 7534 21810 7586
rect 24222 7534 24274 7586
rect 24446 7534 24498 7586
rect 25678 7534 25730 7586
rect 29038 7534 29090 7586
rect 30158 7534 30210 7586
rect 30830 7534 30882 7586
rect 35646 7534 35698 7586
rect 35982 7534 36034 7586
rect 37662 7534 37714 7586
rect 39230 7534 39282 7586
rect 1934 7422 1986 7474
rect 6750 7422 6802 7474
rect 7310 7422 7362 7474
rect 7982 7422 8034 7474
rect 9998 7422 10050 7474
rect 10222 7422 10274 7474
rect 13582 7422 13634 7474
rect 13806 7422 13858 7474
rect 20974 7422 21026 7474
rect 21086 7422 21138 7474
rect 22094 7422 22146 7474
rect 23774 7422 23826 7474
rect 26126 7422 26178 7474
rect 26350 7422 26402 7474
rect 26574 7422 26626 7474
rect 27022 7422 27074 7474
rect 27470 7422 27522 7474
rect 27918 7422 27970 7474
rect 28478 7422 28530 7474
rect 28814 7422 28866 7474
rect 29374 7422 29426 7474
rect 31502 7422 31554 7474
rect 32510 7422 32562 7474
rect 4846 7310 4898 7362
rect 5294 7310 5346 7362
rect 8654 7310 8706 7362
rect 22542 7310 22594 7362
rect 28590 7310 28642 7362
rect 29598 7310 29650 7362
rect 31166 7310 31218 7362
rect 33854 7310 33906 7362
rect 35310 7310 35362 7362
rect 36542 7310 36594 7362
rect 38110 7310 38162 7362
rect 7310 7198 7362 7250
rect 7646 7198 7698 7250
rect 8094 7198 8146 7250
rect 24110 7198 24162 7250
rect 26014 7198 26066 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 8990 6862 9042 6914
rect 9774 6862 9826 6914
rect 29710 6862 29762 6914
rect 33294 6862 33346 6914
rect 6862 6750 6914 6802
rect 10558 6750 10610 6802
rect 13694 6750 13746 6802
rect 20750 6750 20802 6802
rect 23550 6750 23602 6802
rect 25678 6750 25730 6802
rect 36990 6750 37042 6802
rect 37102 6750 37154 6802
rect 38222 6750 38274 6802
rect 7198 6638 7250 6690
rect 9326 6638 9378 6690
rect 10334 6638 10386 6690
rect 11230 6638 11282 6690
rect 11678 6638 11730 6690
rect 14142 6638 14194 6690
rect 14590 6638 14642 6690
rect 15374 6638 15426 6690
rect 15598 6638 15650 6690
rect 16382 6638 16434 6690
rect 16718 6638 16770 6690
rect 17054 6638 17106 6690
rect 17838 6638 17890 6690
rect 18622 6638 18674 6690
rect 22878 6638 22930 6690
rect 28142 6638 28194 6690
rect 29374 6638 29426 6690
rect 34414 6638 34466 6690
rect 34750 6638 34802 6690
rect 35758 6638 35810 6690
rect 7758 6526 7810 6578
rect 8430 6526 8482 6578
rect 15150 6526 15202 6578
rect 16942 6526 16994 6578
rect 28366 6526 28418 6578
rect 29150 6526 29202 6578
rect 34302 6526 34354 6578
rect 34862 6526 34914 6578
rect 36318 6526 36370 6578
rect 37214 6526 37266 6578
rect 39118 6526 39170 6578
rect 8094 6414 8146 6466
rect 8878 6414 8930 6466
rect 9998 6414 10050 6466
rect 10894 6414 10946 6466
rect 12686 6414 12738 6466
rect 15038 6414 15090 6466
rect 15262 6414 15314 6466
rect 17502 6414 17554 6466
rect 26126 6414 26178 6466
rect 29598 6414 29650 6466
rect 33406 6414 33458 6466
rect 33518 6414 33570 6466
rect 35870 6414 35922 6466
rect 37774 6414 37826 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4958 6078 5010 6130
rect 5406 6078 5458 6130
rect 10558 6078 10610 6130
rect 11454 6078 11506 6130
rect 12686 6078 12738 6130
rect 13470 6078 13522 6130
rect 13918 6078 13970 6130
rect 16942 6078 16994 6130
rect 18398 6078 18450 6130
rect 22878 6078 22930 6130
rect 24670 6078 24722 6130
rect 28254 6078 28306 6130
rect 29262 6078 29314 6130
rect 34190 6078 34242 6130
rect 39118 6078 39170 6130
rect 5630 5966 5682 6018
rect 5742 5966 5794 6018
rect 11790 5966 11842 6018
rect 14254 5966 14306 6018
rect 15150 5966 15202 6018
rect 15822 5966 15874 6018
rect 25342 5966 25394 6018
rect 25566 5966 25618 6018
rect 35758 5966 35810 6018
rect 38334 5966 38386 6018
rect 6078 5854 6130 5906
rect 9662 5854 9714 5906
rect 10334 5854 10386 5906
rect 11006 5854 11058 5906
rect 13134 5854 13186 5906
rect 15374 5854 15426 5906
rect 16158 5854 16210 5906
rect 16494 5854 16546 5906
rect 17390 5854 17442 5906
rect 17838 5854 17890 5906
rect 21870 5854 21922 5906
rect 22318 5854 22370 5906
rect 28590 5854 28642 5906
rect 29038 5854 29090 5906
rect 39342 5854 39394 5906
rect 9886 5742 9938 5794
rect 10446 5742 10498 5794
rect 12910 5742 12962 5794
rect 16270 5742 16322 5794
rect 17614 5742 17666 5794
rect 21422 5742 21474 5794
rect 32286 5742 32338 5794
rect 33406 5742 33458 5794
rect 33630 5742 33682 5794
rect 34526 5742 34578 5794
rect 7086 5630 7138 5682
rect 9998 5630 10050 5682
rect 14366 5630 14418 5682
rect 17950 5630 18002 5682
rect 25230 5630 25282 5682
rect 33854 5630 33906 5682
rect 36206 5630 36258 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 8878 5294 8930 5346
rect 12798 5294 12850 5346
rect 21646 5294 21698 5346
rect 35870 5294 35922 5346
rect 4734 5182 4786 5234
rect 5630 5182 5682 5234
rect 7758 5182 7810 5234
rect 8990 5182 9042 5234
rect 10334 5182 10386 5234
rect 12462 5182 12514 5234
rect 14142 5182 14194 5234
rect 16270 5182 16322 5234
rect 17614 5182 17666 5234
rect 22094 5182 22146 5234
rect 24670 5182 24722 5234
rect 26798 5182 26850 5234
rect 27246 5182 27298 5234
rect 28590 5182 28642 5234
rect 29262 5182 29314 5234
rect 31390 5182 31442 5234
rect 33406 5182 33458 5234
rect 35534 5182 35586 5234
rect 39230 5182 39282 5234
rect 1934 5070 1986 5122
rect 8542 5070 8594 5122
rect 9214 5070 9266 5122
rect 9550 5070 9602 5122
rect 13582 5070 13634 5122
rect 16942 5070 16994 5122
rect 21310 5070 21362 5122
rect 23886 5070 23938 5122
rect 32062 5070 32114 5122
rect 32622 5070 32674 5122
rect 2606 4958 2658 5010
rect 12910 4958 12962 5010
rect 36094 4958 36146 5010
rect 37102 4958 37154 5010
rect 13806 4846 13858 4898
rect 21534 4846 21586 4898
rect 35982 4846 36034 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 3950 4510 4002 4562
rect 4958 4510 5010 4562
rect 5854 4510 5906 4562
rect 5966 4510 6018 4562
rect 22990 4510 23042 4562
rect 29710 4510 29762 4562
rect 32510 4510 32562 4562
rect 17390 4398 17442 4450
rect 18174 4398 18226 4450
rect 21758 4398 21810 4450
rect 26238 4398 26290 4450
rect 31950 4398 32002 4450
rect 32174 4398 32226 4450
rect 33518 4398 33570 4450
rect 35198 4398 35250 4450
rect 4734 4286 4786 4338
rect 8990 4286 9042 4338
rect 12014 4286 12066 4338
rect 14926 4286 14978 4338
rect 22542 4286 22594 4338
rect 25454 4286 25506 4338
rect 28814 4286 28866 4338
rect 29038 4286 29090 4338
rect 29262 4286 29314 4338
rect 36654 4286 36706 4338
rect 3838 4174 3890 4226
rect 7198 4174 7250 4226
rect 19630 4174 19682 4226
rect 28366 4174 28418 4226
rect 31502 4174 31554 4226
rect 34526 4174 34578 4226
rect 36318 4174 36370 4226
rect 37438 4174 37490 4226
rect 39566 4174 39618 4226
rect 6078 4062 6130 4114
rect 10110 4062 10162 4114
rect 13022 4062 13074 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 35534 3726 35586 3778
rect 35870 3726 35922 3778
rect 38782 3726 38834 3778
rect 7758 3614 7810 3666
rect 9550 3614 9602 3666
rect 11230 3614 11282 3666
rect 28702 3614 28754 3666
rect 38894 3614 38946 3666
rect 5070 3502 5122 3554
rect 5742 3502 5794 3554
rect 8654 3502 8706 3554
rect 12126 3502 12178 3554
rect 13246 3502 13298 3554
rect 14030 3502 14082 3554
rect 16942 3502 16994 3554
rect 31278 3502 31330 3554
rect 32622 3502 32674 3554
rect 3166 3390 3218 3442
rect 3390 3390 3442 3442
rect 3726 3390 3778 3442
rect 5518 3390 5570 3442
rect 18510 3390 18562 3442
rect 31054 3390 31106 3442
rect 31614 3390 31666 3442
rect 32286 3390 32338 3442
rect 33406 3390 33458 3442
rect 37998 3390 38050 3442
rect 39006 3390 39058 3442
rect 14814 3278 14866 3330
rect 19854 3278 19906 3330
rect 20862 3278 20914 3330
rect 22206 3278 22258 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 9996 39730 10052 39742
rect 9996 39678 9998 39730
rect 10050 39678 10052 39730
rect 9996 38836 10052 39678
rect 17724 39732 17780 39742
rect 12908 39618 12964 39630
rect 12908 39566 12910 39618
rect 12962 39566 12964 39618
rect 12124 39506 12180 39518
rect 12124 39454 12126 39506
rect 12178 39454 12180 39506
rect 11788 39060 11844 39070
rect 9996 38770 10052 38780
rect 11340 38836 11396 38846
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 9660 38276 9716 38286
rect 9660 38050 9716 38220
rect 10556 38276 10612 38286
rect 9996 38164 10052 38174
rect 9660 37998 9662 38050
rect 9714 37998 9716 38050
rect 9660 37986 9716 37998
rect 9884 38108 9996 38164
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 6188 35698 6244 35710
rect 6188 35646 6190 35698
rect 6242 35646 6244 35698
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 5628 35252 5684 35262
rect 5628 34914 5684 35196
rect 6188 35252 6244 35646
rect 6188 35186 6244 35196
rect 6860 35586 6916 35598
rect 6860 35534 6862 35586
rect 6914 35534 6916 35586
rect 6412 35028 6468 35038
rect 6412 34934 6468 34972
rect 5628 34862 5630 34914
rect 5682 34862 5684 34914
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 2828 30994 2884 31006
rect 2828 30942 2830 30994
rect 2882 30942 2884 30994
rect 1932 29428 1988 29438
rect 1932 29334 1988 29372
rect 2828 29428 2884 30942
rect 3612 30882 3668 30894
rect 3612 30830 3614 30882
rect 3666 30830 3668 30882
rect 3612 30436 3668 30830
rect 5628 30660 5684 34862
rect 6860 33460 6916 35534
rect 8988 35586 9044 35598
rect 8988 35534 8990 35586
rect 9042 35534 9044 35586
rect 8988 35140 9044 35534
rect 8988 35074 9044 35084
rect 9660 35586 9716 35598
rect 9660 35534 9662 35586
rect 9714 35534 9716 35586
rect 9660 35252 9716 35534
rect 8540 35028 8596 35038
rect 8316 35026 8932 35028
rect 8316 34974 8542 35026
rect 8594 34974 8932 35026
rect 8316 34972 8932 34974
rect 6860 33394 6916 33404
rect 7980 33460 8036 33470
rect 8316 33460 8372 34972
rect 8540 34962 8596 34972
rect 8876 34914 8932 34972
rect 9660 35026 9716 35196
rect 9660 34974 9662 35026
rect 9714 34974 9716 35026
rect 9660 34962 9716 34974
rect 8876 34862 8878 34914
rect 8930 34862 8932 34914
rect 8876 34850 8932 34862
rect 9212 34692 9268 34702
rect 9212 34690 9380 34692
rect 9212 34638 9214 34690
rect 9266 34638 9380 34690
rect 9212 34636 9380 34638
rect 9212 34626 9268 34636
rect 9212 33460 9268 33470
rect 7980 33458 8372 33460
rect 7980 33406 7982 33458
rect 8034 33406 8372 33458
rect 7980 33404 8372 33406
rect 8876 33458 9268 33460
rect 8876 33406 9214 33458
rect 9266 33406 9268 33458
rect 8876 33404 9268 33406
rect 7980 33394 8036 33404
rect 7308 33348 7364 33358
rect 6972 33346 7364 33348
rect 6972 33294 7310 33346
rect 7362 33294 7364 33346
rect 6972 33292 7364 33294
rect 6636 30994 6692 31006
rect 6636 30942 6638 30994
rect 6690 30942 6692 30994
rect 5740 30882 5796 30894
rect 5740 30830 5742 30882
rect 5794 30830 5796 30882
rect 5740 30772 5796 30830
rect 6412 30882 6468 30894
rect 6412 30830 6414 30882
rect 6466 30830 6468 30882
rect 6412 30772 6468 30830
rect 5740 30716 6468 30772
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5180 30604 6020 30660
rect 3612 30370 3668 30380
rect 2828 29362 2884 29372
rect 5180 29650 5236 30604
rect 5964 30210 6020 30604
rect 5964 30158 5966 30210
rect 6018 30158 6020 30210
rect 5964 30146 6020 30158
rect 6412 30210 6468 30716
rect 6412 30158 6414 30210
rect 6466 30158 6468 30210
rect 6412 30146 6468 30158
rect 5180 29598 5182 29650
rect 5234 29598 5236 29650
rect 5180 29428 5236 29598
rect 5180 29362 5236 29372
rect 2604 29316 2660 29326
rect 4732 29316 4788 29326
rect 2604 29314 2772 29316
rect 2604 29262 2606 29314
rect 2658 29262 2772 29314
rect 2604 29260 2772 29262
rect 2604 29250 2660 29260
rect 2716 27300 2772 29260
rect 4732 29222 4788 29260
rect 6636 29316 6692 30942
rect 6748 29986 6804 29998
rect 6748 29934 6750 29986
rect 6802 29934 6804 29986
rect 6748 29540 6804 29934
rect 6748 29474 6804 29484
rect 6636 29092 6692 29260
rect 4476 29036 4740 29046
rect 6636 29036 6916 29092
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 3836 27858 3892 27870
rect 3836 27806 3838 27858
rect 3890 27806 3892 27858
rect 2716 27244 3220 27300
rect 1820 27074 1876 27086
rect 1820 27022 1822 27074
rect 1874 27022 1876 27074
rect 1820 26964 1876 27022
rect 1820 26898 1876 26908
rect 2492 26962 2548 26974
rect 2492 26910 2494 26962
rect 2546 26910 2548 26962
rect 2380 24948 2436 24958
rect 2492 24948 2548 26910
rect 3164 25730 3220 27244
rect 3836 26964 3892 27806
rect 4620 27748 4676 27758
rect 6748 27748 6804 27758
rect 4620 27746 4900 27748
rect 4620 27694 4622 27746
rect 4674 27694 4900 27746
rect 4620 27692 4900 27694
rect 4620 27682 4676 27692
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 3836 26898 3892 26908
rect 4620 27186 4676 27198
rect 4620 27134 4622 27186
rect 4674 27134 4676 27186
rect 4620 26292 4676 27134
rect 4620 26226 4676 26236
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3164 25678 3166 25730
rect 3218 25678 3220 25730
rect 3164 25666 3220 25678
rect 3500 25396 3556 25406
rect 3500 25394 4340 25396
rect 3500 25342 3502 25394
rect 3554 25342 4340 25394
rect 3500 25340 4340 25342
rect 3500 25330 3556 25340
rect 2380 24946 2548 24948
rect 2380 24894 2382 24946
rect 2434 24894 2548 24946
rect 2380 24892 2548 24894
rect 3276 25282 3332 25294
rect 3276 25230 3278 25282
rect 3330 25230 3332 25282
rect 2380 24882 2436 24892
rect 2268 24834 2324 24846
rect 2268 24782 2270 24834
rect 2322 24782 2324 24834
rect 2268 22708 2324 24782
rect 2492 24724 2548 24734
rect 2828 24724 2884 24734
rect 2492 24722 2884 24724
rect 2492 24670 2494 24722
rect 2546 24670 2830 24722
rect 2882 24670 2884 24722
rect 2492 24668 2884 24670
rect 2492 24658 2548 24668
rect 2828 24658 2884 24668
rect 3276 23940 3332 25230
rect 4284 24834 4340 25340
rect 4284 24782 4286 24834
rect 4338 24782 4340 24834
rect 4284 24770 4340 24782
rect 3276 23604 3332 23884
rect 3500 24724 3556 24734
rect 3500 23716 3556 24668
rect 4396 24722 4452 24734
rect 4396 24670 4398 24722
rect 4450 24670 4452 24722
rect 3612 24610 3668 24622
rect 3612 24558 3614 24610
rect 3666 24558 3668 24610
rect 3612 23940 3668 24558
rect 4396 24500 4452 24670
rect 4060 24444 4452 24500
rect 3724 23940 3780 23950
rect 3612 23938 4004 23940
rect 3612 23886 3726 23938
rect 3778 23886 4004 23938
rect 3612 23884 4004 23886
rect 3724 23874 3780 23884
rect 3836 23716 3892 23726
rect 3500 23714 3892 23716
rect 3500 23662 3838 23714
rect 3890 23662 3892 23714
rect 3500 23660 3892 23662
rect 3948 23716 4004 23884
rect 4060 23938 4116 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4844 24164 4900 27692
rect 6748 27654 6804 27692
rect 5068 26964 5124 27002
rect 5068 26898 5124 26908
rect 6860 26628 6916 29036
rect 6860 26562 6916 26572
rect 6636 26402 6692 26414
rect 6636 26350 6638 26402
rect 6690 26350 6692 26402
rect 6412 26292 6468 26302
rect 6412 25508 6468 26236
rect 6412 25442 6468 25452
rect 6636 26292 6692 26350
rect 6972 26292 7028 33292
rect 7308 33282 7364 33292
rect 8204 33236 8260 33246
rect 8204 33142 8260 33180
rect 8428 31890 8484 31902
rect 8428 31838 8430 31890
rect 8482 31838 8484 31890
rect 7196 31108 7252 31118
rect 7196 31014 7252 31052
rect 8428 31108 8484 31838
rect 8876 31778 8932 33404
rect 9212 33394 9268 33404
rect 9324 33348 9380 34636
rect 9324 33254 9380 33292
rect 9548 34020 9604 34030
rect 8876 31726 8878 31778
rect 8930 31726 8932 31778
rect 8876 31714 8932 31726
rect 9100 33234 9156 33246
rect 9100 33182 9102 33234
rect 9154 33182 9156 33234
rect 8428 31042 8484 31052
rect 8764 31220 8820 31230
rect 8540 30996 8596 31006
rect 8764 30996 8820 31164
rect 8540 30902 8596 30940
rect 8652 30994 8820 30996
rect 8652 30942 8766 30994
rect 8818 30942 8820 30994
rect 8652 30940 8820 30942
rect 8092 30210 8148 30222
rect 8092 30158 8094 30210
rect 8146 30158 8148 30210
rect 7980 28868 8036 28878
rect 7980 28642 8036 28812
rect 7980 28590 7982 28642
rect 8034 28590 8036 28642
rect 7980 28578 8036 28590
rect 7868 27860 7924 27870
rect 7756 27858 7924 27860
rect 7756 27806 7870 27858
rect 7922 27806 7924 27858
rect 7756 27804 7924 27806
rect 7756 27412 7812 27804
rect 7868 27794 7924 27804
rect 6636 26236 7028 26292
rect 7084 27356 7812 27412
rect 6636 25284 6692 26236
rect 6636 25228 6804 25284
rect 5740 24948 5796 24958
rect 4956 24836 5012 24846
rect 4956 24722 5012 24780
rect 4956 24670 4958 24722
rect 5010 24670 5012 24722
rect 4956 24658 5012 24670
rect 5740 24722 5796 24892
rect 5964 24836 6020 24846
rect 6020 24780 6356 24836
rect 5964 24742 6020 24780
rect 5740 24670 5742 24722
rect 5794 24670 5796 24722
rect 5740 24658 5796 24670
rect 4732 24108 4900 24164
rect 4060 23886 4062 23938
rect 4114 23886 4116 23938
rect 4060 23874 4116 23886
rect 4396 23940 4452 23950
rect 4396 23846 4452 23884
rect 4620 23938 4676 23950
rect 4620 23886 4622 23938
rect 4674 23886 4676 23938
rect 4620 23716 4676 23886
rect 3948 23660 4676 23716
rect 3836 23650 3892 23660
rect 3276 23548 3556 23604
rect 3164 23266 3220 23278
rect 3164 23214 3166 23266
rect 3218 23214 3220 23266
rect 3164 22708 3220 23214
rect 3500 23154 3556 23548
rect 4620 23380 4676 23660
rect 4732 23714 4788 24108
rect 5628 24050 5684 24062
rect 5628 23998 5630 24050
rect 5682 23998 5684 24050
rect 4844 23940 4900 23950
rect 4844 23846 4900 23884
rect 5628 23940 5684 23998
rect 5628 23874 5684 23884
rect 5964 23828 6020 23838
rect 5964 23826 6132 23828
rect 5964 23774 5966 23826
rect 6018 23774 6132 23826
rect 5964 23772 6132 23774
rect 5964 23762 6020 23772
rect 5740 23716 5796 23726
rect 4732 23662 4734 23714
rect 4786 23662 4788 23714
rect 4732 23650 4788 23662
rect 5292 23714 5908 23716
rect 5292 23662 5742 23714
rect 5794 23662 5908 23714
rect 5292 23660 5908 23662
rect 4732 23380 4788 23390
rect 4620 23378 4788 23380
rect 4620 23326 4734 23378
rect 4786 23326 4788 23378
rect 4620 23324 4788 23326
rect 4732 23314 4788 23324
rect 3500 23102 3502 23154
rect 3554 23102 3556 23154
rect 3500 22932 3556 23102
rect 5292 23154 5348 23660
rect 5740 23650 5796 23660
rect 5292 23102 5294 23154
rect 5346 23102 5348 23154
rect 5292 23090 5348 23102
rect 3500 22866 3556 22876
rect 5068 22930 5124 22942
rect 5068 22878 5070 22930
rect 5122 22878 5124 22930
rect 2268 22652 3220 22708
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 1820 20802 1876 20814
rect 1820 20750 1822 20802
rect 1874 20750 1876 20802
rect 1820 17668 1876 20750
rect 2492 20690 2548 20702
rect 2492 20638 2494 20690
rect 2546 20638 2548 20690
rect 2492 20188 2548 20638
rect 2492 20132 2884 20188
rect 2828 19906 2884 20132
rect 2828 19854 2830 19906
rect 2882 19854 2884 19906
rect 2828 19842 2884 19854
rect 2940 20130 2996 22652
rect 5068 22148 5124 22878
rect 5852 22820 5908 23660
rect 6076 23156 6132 23772
rect 5852 22764 6020 22820
rect 5852 22484 5908 22494
rect 5852 22370 5908 22428
rect 5852 22318 5854 22370
rect 5906 22318 5908 22370
rect 5852 22306 5908 22318
rect 5964 22372 6020 22764
rect 5964 22258 6020 22316
rect 5964 22206 5966 22258
rect 6018 22206 6020 22258
rect 5964 22194 6020 22206
rect 5068 22082 5124 22092
rect 5852 22148 5908 22158
rect 5852 22036 5908 22092
rect 6076 22036 6132 23100
rect 6300 22484 6356 24780
rect 6524 24834 6580 24846
rect 6524 24782 6526 24834
rect 6578 24782 6580 24834
rect 6524 24724 6580 24782
rect 6748 24836 6804 25228
rect 6860 24836 6916 24846
rect 6748 24834 6916 24836
rect 6748 24782 6862 24834
rect 6914 24782 6916 24834
rect 6748 24780 6916 24782
rect 6860 24724 6916 24780
rect 6972 24724 7028 24734
rect 6580 24668 6692 24724
rect 6860 24668 6972 24724
rect 6524 24658 6580 24668
rect 6636 23604 6692 24668
rect 6972 24658 7028 24668
rect 7084 23716 7140 27356
rect 7196 26964 7252 27002
rect 8092 26908 8148 30158
rect 8652 30210 8708 30940
rect 8764 30930 8820 30940
rect 8988 30994 9044 31006
rect 8988 30942 8990 30994
rect 9042 30942 9044 30994
rect 8652 30158 8654 30210
rect 8706 30158 8708 30210
rect 8652 30146 8708 30158
rect 8764 30324 8820 30334
rect 8764 30210 8820 30268
rect 8764 30158 8766 30210
rect 8818 30158 8820 30210
rect 8764 30146 8820 30158
rect 8652 29428 8708 29438
rect 8428 29316 8484 29326
rect 8428 28642 8484 29260
rect 8540 28756 8596 28766
rect 8540 28662 8596 28700
rect 8428 28590 8430 28642
rect 8482 28590 8484 28642
rect 8428 28578 8484 28590
rect 8652 28642 8708 29372
rect 8876 28868 8932 28878
rect 8652 28590 8654 28642
rect 8706 28590 8708 28642
rect 8652 28578 8708 28590
rect 8764 28644 8820 28654
rect 8428 28084 8484 28094
rect 8428 27858 8484 28028
rect 8540 27972 8596 27982
rect 8764 27972 8820 28588
rect 8540 27970 8820 27972
rect 8540 27918 8542 27970
rect 8594 27918 8820 27970
rect 8540 27916 8820 27918
rect 8540 27906 8596 27916
rect 8428 27806 8430 27858
rect 8482 27806 8484 27858
rect 8428 27794 8484 27806
rect 8876 27186 8932 28812
rect 8988 28530 9044 30942
rect 9100 29316 9156 33182
rect 9548 33234 9604 33964
rect 9548 33182 9550 33234
rect 9602 33182 9604 33234
rect 9548 33170 9604 33182
rect 9660 33236 9716 33246
rect 9660 32452 9716 33180
rect 9884 33012 9940 38108
rect 9996 38070 10052 38108
rect 10556 38162 10612 38220
rect 10556 38110 10558 38162
rect 10610 38110 10612 38162
rect 10556 38098 10612 38110
rect 11340 38050 11396 38780
rect 11676 38724 11732 38734
rect 11676 38630 11732 38668
rect 11340 37998 11342 38050
rect 11394 37998 11396 38050
rect 11228 34802 11284 34814
rect 11228 34750 11230 34802
rect 11282 34750 11284 34802
rect 10444 34020 10500 34030
rect 10444 33926 10500 33964
rect 10556 33908 10612 33918
rect 11228 33908 11284 34750
rect 11340 34020 11396 37998
rect 11564 38052 11620 38062
rect 11564 37938 11620 37996
rect 11564 37886 11566 37938
rect 11618 37886 11620 37938
rect 11564 37874 11620 37886
rect 11564 36372 11620 36382
rect 11564 35138 11620 36316
rect 11564 35086 11566 35138
rect 11618 35086 11620 35138
rect 11564 35074 11620 35086
rect 11788 35252 11844 39004
rect 12124 39058 12180 39454
rect 12124 39006 12126 39058
rect 12178 39006 12180 39058
rect 12124 38994 12180 39006
rect 12908 39060 12964 39566
rect 15708 39618 15764 39630
rect 15708 39566 15710 39618
rect 15762 39566 15764 39618
rect 12908 38994 12964 39004
rect 13580 39394 13636 39406
rect 13580 39342 13582 39394
rect 13634 39342 13636 39394
rect 13580 39060 13636 39342
rect 13580 38994 13636 39004
rect 15372 39396 15428 39406
rect 15708 39396 15764 39566
rect 16492 39508 16548 39518
rect 16492 39506 16772 39508
rect 16492 39454 16494 39506
rect 16546 39454 16772 39506
rect 16492 39452 16772 39454
rect 16492 39442 16548 39452
rect 15372 39394 15764 39396
rect 15372 39342 15374 39394
rect 15426 39342 15764 39394
rect 15372 39340 15764 39342
rect 15372 39060 15428 39340
rect 16492 39060 16548 39070
rect 15372 38994 15428 39004
rect 16380 39058 16548 39060
rect 16380 39006 16494 39058
rect 16546 39006 16548 39058
rect 16380 39004 16548 39006
rect 12012 38946 12068 38958
rect 12012 38894 12014 38946
rect 12066 38894 12068 38946
rect 12012 38724 12068 38894
rect 15036 38946 15092 38958
rect 15036 38894 15038 38946
rect 15090 38894 15092 38946
rect 12684 38836 12740 38846
rect 12684 38742 12740 38780
rect 13132 38834 13188 38846
rect 13132 38782 13134 38834
rect 13186 38782 13188 38834
rect 12012 38612 12180 38668
rect 12012 38276 12068 38286
rect 11564 34914 11620 34926
rect 11564 34862 11566 34914
rect 11618 34862 11620 34914
rect 11564 34356 11620 34862
rect 11564 34290 11620 34300
rect 11340 33954 11396 33964
rect 10556 33906 11284 33908
rect 10556 33854 10558 33906
rect 10610 33854 11284 33906
rect 10556 33852 11284 33854
rect 10556 33572 10612 33852
rect 10332 33516 10612 33572
rect 11340 33572 11396 33582
rect 9996 33346 10052 33358
rect 9996 33294 9998 33346
rect 10050 33294 10052 33346
rect 9996 33236 10052 33294
rect 9996 33170 10052 33180
rect 9884 32956 10052 33012
rect 9548 32396 9716 32452
rect 9324 31666 9380 31678
rect 9324 31614 9326 31666
rect 9378 31614 9380 31666
rect 9324 30212 9380 31614
rect 9548 30994 9604 32396
rect 9660 31668 9716 31678
rect 9660 31666 9828 31668
rect 9660 31614 9662 31666
rect 9714 31614 9828 31666
rect 9660 31612 9828 31614
rect 9660 31602 9716 31612
rect 9660 31108 9716 31118
rect 9660 31014 9716 31052
rect 9548 30942 9550 30994
rect 9602 30942 9604 30994
rect 9548 30930 9604 30942
rect 9772 30996 9828 31612
rect 9884 30996 9940 31006
rect 9772 30994 9940 30996
rect 9772 30942 9886 30994
rect 9938 30942 9940 30994
rect 9772 30940 9940 30942
rect 9324 30146 9380 30156
rect 9884 29428 9940 30940
rect 9996 30996 10052 32956
rect 10332 31892 10388 33516
rect 10444 33346 10500 33358
rect 10444 33294 10446 33346
rect 10498 33294 10500 33346
rect 10444 33012 10500 33294
rect 10892 33348 10948 33358
rect 10892 33346 11284 33348
rect 10892 33294 10894 33346
rect 10946 33294 11284 33346
rect 10892 33292 11284 33294
rect 10892 33282 10948 33292
rect 11116 33122 11172 33134
rect 11116 33070 11118 33122
rect 11170 33070 11172 33122
rect 11116 33012 11172 33070
rect 10444 32956 11172 33012
rect 10444 31892 10500 31902
rect 10332 31890 10500 31892
rect 10332 31838 10446 31890
rect 10498 31838 10500 31890
rect 10332 31836 10500 31838
rect 10444 31826 10500 31836
rect 11228 31892 11284 33292
rect 11340 33234 11396 33516
rect 11340 33182 11342 33234
rect 11394 33182 11396 33234
rect 11340 33170 11396 33182
rect 11452 33234 11508 33246
rect 11452 33182 11454 33234
rect 11506 33182 11508 33234
rect 11228 31826 11284 31836
rect 10108 31780 10164 31790
rect 10108 31778 10388 31780
rect 10108 31726 10110 31778
rect 10162 31726 10388 31778
rect 10108 31724 10388 31726
rect 10108 31714 10164 31724
rect 9996 30930 10052 30940
rect 10108 30994 10164 31006
rect 10108 30942 10110 30994
rect 10162 30942 10164 30994
rect 10108 30324 10164 30942
rect 10108 30258 10164 30268
rect 10220 30212 10276 30222
rect 10220 30118 10276 30156
rect 9884 29362 9940 29372
rect 10108 29988 10164 29998
rect 10108 29426 10164 29932
rect 10332 29652 10388 31724
rect 11228 31554 11284 31566
rect 11228 31502 11230 31554
rect 11282 31502 11284 31554
rect 11228 31220 11284 31502
rect 11228 31154 11284 31164
rect 10556 30772 10612 30782
rect 10556 30770 10724 30772
rect 10556 30718 10558 30770
rect 10610 30718 10724 30770
rect 10556 30716 10724 30718
rect 10556 30706 10612 30716
rect 10556 30212 10612 30222
rect 10108 29374 10110 29426
rect 10162 29374 10164 29426
rect 9100 29250 9156 29260
rect 10108 29316 10164 29374
rect 10108 29250 10164 29260
rect 10220 29596 10388 29652
rect 10444 30210 10612 30212
rect 10444 30158 10558 30210
rect 10610 30158 10612 30210
rect 10444 30156 10612 30158
rect 10444 29650 10500 30156
rect 10556 30146 10612 30156
rect 10444 29598 10446 29650
rect 10498 29598 10500 29650
rect 10220 28868 10276 29596
rect 10444 29586 10500 29598
rect 10556 29764 10612 29774
rect 10556 29650 10612 29708
rect 10556 29598 10558 29650
rect 10610 29598 10612 29650
rect 10556 29586 10612 29598
rect 10668 29652 10724 30716
rect 10780 30156 11060 30212
rect 10780 30098 10836 30156
rect 10780 30046 10782 30098
rect 10834 30046 10836 30098
rect 10780 30034 10836 30046
rect 10668 29586 10724 29596
rect 10892 29986 10948 29998
rect 10892 29934 10894 29986
rect 10946 29934 10948 29986
rect 10332 29428 10388 29438
rect 10668 29428 10724 29438
rect 10332 29334 10388 29372
rect 10444 29426 10836 29428
rect 10444 29374 10670 29426
rect 10722 29374 10836 29426
rect 10444 29372 10836 29374
rect 10220 28812 10388 28868
rect 9436 28756 9492 28766
rect 9436 28662 9492 28700
rect 8988 28478 8990 28530
rect 9042 28478 9044 28530
rect 8988 28466 9044 28478
rect 9212 28642 9268 28654
rect 9212 28590 9214 28642
rect 9266 28590 9268 28642
rect 8988 28084 9044 28094
rect 8988 27990 9044 28028
rect 8876 27134 8878 27186
rect 8930 27134 8932 27186
rect 8876 27122 8932 27134
rect 9212 27860 9268 28590
rect 9548 28644 9604 28654
rect 9548 28550 9604 28588
rect 10220 28644 10276 28654
rect 10220 28550 10276 28588
rect 7196 24612 7252 26908
rect 7980 26852 8148 26908
rect 7532 26628 7588 26638
rect 7308 25508 7364 25518
rect 7308 25414 7364 25452
rect 7532 25396 7588 26572
rect 7532 25394 7924 25396
rect 7532 25342 7534 25394
rect 7586 25342 7924 25394
rect 7532 25340 7924 25342
rect 7532 25330 7588 25340
rect 7868 24948 7924 25340
rect 7196 24546 7252 24556
rect 7644 24724 7700 24734
rect 7644 23826 7700 24668
rect 7644 23774 7646 23826
rect 7698 23774 7700 23826
rect 7084 23660 7364 23716
rect 6636 23548 7028 23604
rect 6300 22370 6356 22428
rect 6860 23266 6916 23278
rect 6860 23214 6862 23266
rect 6914 23214 6916 23266
rect 6300 22318 6302 22370
rect 6354 22318 6356 22370
rect 6300 22306 6356 22318
rect 6748 22372 6804 22382
rect 6860 22372 6916 23214
rect 6804 22316 6916 22372
rect 6972 22370 7028 23548
rect 6972 22318 6974 22370
rect 7026 22318 7028 22370
rect 6748 22278 6804 22316
rect 6188 22148 6244 22158
rect 6188 22146 6468 22148
rect 6188 22094 6190 22146
rect 6242 22094 6468 22146
rect 6188 22092 6468 22094
rect 6188 22082 6244 22092
rect 5852 21980 6132 22036
rect 3724 21588 3780 21598
rect 3724 21494 3780 21532
rect 5068 21588 5124 21598
rect 5068 21494 5124 21532
rect 3052 21474 3108 21486
rect 3052 21422 3054 21474
rect 3106 21422 3108 21474
rect 3052 20188 3108 21422
rect 3948 21474 4004 21486
rect 3948 21422 3950 21474
rect 4002 21422 4004 21474
rect 3052 20132 3220 20188
rect 3948 20132 4004 21422
rect 5404 21474 5460 21486
rect 5404 21422 5406 21474
rect 5458 21422 5460 21474
rect 4956 21364 5012 21374
rect 4844 21308 4956 21364
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4844 21028 4900 21308
rect 4956 21298 5012 21308
rect 5404 21364 5460 21422
rect 5404 21298 5460 21308
rect 4620 20972 4900 21028
rect 4620 20914 4676 20972
rect 4620 20862 4622 20914
rect 4674 20862 4676 20914
rect 4620 20850 4676 20862
rect 5516 20692 5572 20702
rect 5068 20580 5124 20590
rect 5068 20578 5236 20580
rect 5068 20526 5070 20578
rect 5122 20526 5236 20578
rect 5068 20524 5236 20526
rect 5068 20514 5124 20524
rect 2940 20078 2942 20130
rect 2994 20078 2996 20130
rect 2492 19124 2548 19134
rect 2492 17778 2548 19068
rect 2492 17726 2494 17778
rect 2546 17726 2548 17778
rect 2492 17714 2548 17726
rect 1820 13748 1876 17612
rect 1932 16884 1988 16894
rect 1932 15148 1988 16828
rect 2828 15316 2884 15326
rect 2828 15222 2884 15260
rect 1932 15092 2100 15148
rect 1932 13748 1988 13758
rect 1820 13746 1988 13748
rect 1820 13694 1934 13746
rect 1986 13694 1988 13746
rect 1820 13692 1988 13694
rect 1932 13636 1988 13692
rect 1932 13570 1988 13580
rect 1820 9042 1876 9054
rect 1820 8990 1822 9042
rect 1874 8990 1876 9042
rect 1820 7476 1876 8990
rect 1932 7476 1988 7486
rect 1820 7474 1988 7476
rect 1820 7422 1934 7474
rect 1986 7422 1988 7474
rect 1820 7420 1988 7422
rect 1932 6468 1988 7420
rect 1932 5122 1988 6412
rect 1932 5070 1934 5122
rect 1986 5070 1988 5122
rect 1932 5058 1988 5070
rect 2044 3388 2100 15092
rect 2716 15090 2772 15102
rect 2716 15038 2718 15090
rect 2770 15038 2772 15090
rect 2604 13860 2660 13870
rect 2716 13860 2772 15038
rect 2604 13858 2772 13860
rect 2604 13806 2606 13858
rect 2658 13806 2772 13858
rect 2604 13804 2772 13806
rect 2604 13794 2660 13804
rect 2268 13636 2324 13646
rect 2268 12178 2324 13580
rect 2268 12126 2270 12178
rect 2322 12126 2324 12178
rect 2268 12114 2324 12126
rect 2828 10052 2884 10062
rect 2940 10052 2996 20078
rect 3164 20130 3220 20132
rect 3164 20078 3166 20130
rect 3218 20078 3220 20130
rect 3164 20066 3220 20078
rect 3836 20076 3948 20132
rect 3836 19458 3892 20076
rect 3948 20066 4004 20076
rect 5068 20020 5124 20030
rect 3836 19406 3838 19458
rect 3890 19406 3892 19458
rect 3836 19394 3892 19406
rect 4284 19906 4340 19918
rect 4284 19854 4286 19906
rect 4338 19854 4340 19906
rect 4284 19348 4340 19854
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4284 19292 4452 19348
rect 3612 19234 3668 19246
rect 3612 19182 3614 19234
rect 3666 19182 3668 19234
rect 3500 19124 3556 19134
rect 3500 19030 3556 19068
rect 3612 18900 3668 19182
rect 4060 19236 4116 19246
rect 4060 19234 4340 19236
rect 4060 19182 4062 19234
rect 4114 19182 4340 19234
rect 4060 19180 4340 19182
rect 4060 19170 4116 19180
rect 3500 18844 3612 18900
rect 3052 16772 3108 16782
rect 3052 15314 3108 16716
rect 3500 16210 3556 18844
rect 3612 18834 3668 18844
rect 4284 18674 4340 19180
rect 4396 18900 4452 19292
rect 4732 19236 4788 19246
rect 4732 19124 4788 19180
rect 4396 18834 4452 18844
rect 4508 19122 4788 19124
rect 4508 19070 4734 19122
rect 4786 19070 4788 19122
rect 4508 19068 4788 19070
rect 4284 18622 4286 18674
rect 4338 18622 4340 18674
rect 4284 18610 4340 18622
rect 4508 18450 4564 19068
rect 4732 19058 4788 19068
rect 5068 19234 5124 19964
rect 5068 19182 5070 19234
rect 5122 19182 5124 19234
rect 5068 18564 5124 19182
rect 5068 18498 5124 18508
rect 4508 18398 4510 18450
rect 4562 18398 4564 18450
rect 4508 18386 4564 18398
rect 4172 18226 4228 18238
rect 4172 18174 4174 18226
rect 4226 18174 4228 18226
rect 4172 16772 4228 18174
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4620 17780 4676 17790
rect 4620 17686 4676 17724
rect 5068 17780 5124 17790
rect 5180 17780 5236 20524
rect 5068 17778 5236 17780
rect 5068 17726 5070 17778
rect 5122 17726 5236 17778
rect 5068 17724 5236 17726
rect 5068 17668 5124 17724
rect 5068 17602 5124 17612
rect 4172 16706 4228 16716
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 3500 16158 3502 16210
rect 3554 16158 3556 16210
rect 3052 15262 3054 15314
rect 3106 15262 3108 15314
rect 3052 15250 3108 15262
rect 3276 15876 3332 15886
rect 3276 15314 3332 15820
rect 3276 15262 3278 15314
rect 3330 15262 3332 15314
rect 3276 15250 3332 15262
rect 3500 15316 3556 16158
rect 4284 16098 4340 16110
rect 4284 16046 4286 16098
rect 4338 16046 4340 16098
rect 3948 15988 4004 15998
rect 3500 14756 3556 15260
rect 3612 15986 4004 15988
rect 3612 15934 3950 15986
rect 4002 15934 4004 15986
rect 3612 15932 4004 15934
rect 3612 15538 3668 15932
rect 3948 15922 4004 15932
rect 4060 15876 4116 15886
rect 4060 15782 4116 15820
rect 4284 15876 4340 16046
rect 4284 15810 4340 15820
rect 4956 15876 5012 15886
rect 4956 15540 5012 15820
rect 3612 15486 3614 15538
rect 3666 15486 3668 15538
rect 3612 14756 3668 15486
rect 3948 15484 4900 15540
rect 3724 14756 3780 14766
rect 3612 14754 3780 14756
rect 3612 14702 3726 14754
rect 3778 14702 3780 14754
rect 3612 14700 3780 14702
rect 3500 14662 3556 14700
rect 3724 14690 3780 14700
rect 3948 14530 4004 15484
rect 4844 15426 4900 15484
rect 4844 15374 4846 15426
rect 4898 15374 4900 15426
rect 4844 15362 4900 15374
rect 4060 15314 4116 15326
rect 4060 15262 4062 15314
rect 4114 15262 4116 15314
rect 4060 15204 4116 15262
rect 4060 15138 4116 15148
rect 4172 15314 4228 15326
rect 4172 15262 4174 15314
rect 4226 15262 4228 15314
rect 4172 15148 4228 15262
rect 4396 15316 4452 15354
rect 4396 15250 4452 15260
rect 4620 15314 4676 15326
rect 4620 15262 4622 15314
rect 4674 15262 4676 15314
rect 4620 15148 4676 15262
rect 4956 15148 5012 15484
rect 5068 15428 5124 15438
rect 5068 15334 5124 15372
rect 3948 14478 3950 14530
rect 4002 14478 4004 14530
rect 3948 14466 4004 14478
rect 4172 15092 4676 15148
rect 4844 15092 5012 15148
rect 3388 14420 3444 14430
rect 3052 14418 3444 14420
rect 3052 14366 3390 14418
rect 3442 14366 3444 14418
rect 3052 14364 3444 14366
rect 3052 12290 3108 14364
rect 3388 14354 3444 14364
rect 3052 12238 3054 12290
rect 3106 12238 3108 12290
rect 3052 12226 3108 12238
rect 2380 10050 2996 10052
rect 2380 9998 2830 10050
rect 2882 9998 2996 10050
rect 2380 9996 2996 9998
rect 2380 8258 2436 9996
rect 2828 9986 2884 9996
rect 3164 9826 3220 9838
rect 3164 9774 3166 9826
rect 3218 9774 3220 9826
rect 3164 9716 3220 9774
rect 3164 9650 3220 9660
rect 4060 9716 4116 9726
rect 4172 9716 4228 15092
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4508 14756 4564 14766
rect 4508 14642 4564 14700
rect 4508 14590 4510 14642
rect 4562 14590 4564 14642
rect 4508 14578 4564 14590
rect 4732 14420 4788 14430
rect 4844 14420 4900 15092
rect 4732 14418 4900 14420
rect 4732 14366 4734 14418
rect 4786 14366 4900 14418
rect 4732 14364 4900 14366
rect 4956 14532 5012 14542
rect 4732 14354 4788 14364
rect 4956 13748 5012 14476
rect 4732 13692 5012 13748
rect 4732 13634 4788 13692
rect 4732 13582 4734 13634
rect 4786 13582 4788 13634
rect 4732 13570 4788 13582
rect 5180 13636 5236 17724
rect 5292 15314 5348 15326
rect 5292 15262 5294 15314
rect 5346 15262 5348 15314
rect 5292 15204 5348 15262
rect 5292 15138 5348 15148
rect 5180 13542 5236 13580
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 5180 12068 5236 12078
rect 5404 12068 5460 12078
rect 5180 12066 5460 12068
rect 5180 12014 5182 12066
rect 5234 12014 5406 12066
rect 5458 12014 5460 12066
rect 5180 12012 5460 12014
rect 5180 12002 5236 12012
rect 5404 12002 5460 12012
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4116 9660 4228 9716
rect 2940 9602 2996 9614
rect 2940 9550 2942 9602
rect 2994 9550 2996 9602
rect 2940 9268 2996 9550
rect 2492 9212 2996 9268
rect 2492 9154 2548 9212
rect 2492 9102 2494 9154
rect 2546 9102 2548 9154
rect 2492 9090 2548 9102
rect 3948 8372 4004 8382
rect 4060 8372 4116 9660
rect 4396 9602 4452 9614
rect 4396 9550 4398 9602
rect 4450 9550 4452 9602
rect 4396 8932 4452 9550
rect 4620 8932 4676 8942
rect 4396 8930 4676 8932
rect 4396 8878 4622 8930
rect 4674 8878 4676 8930
rect 4396 8876 4676 8878
rect 4620 8820 4676 8876
rect 5068 8932 5124 8942
rect 5068 8930 5236 8932
rect 5068 8878 5070 8930
rect 5122 8878 5236 8930
rect 5068 8876 5236 8878
rect 5068 8866 5124 8876
rect 4620 8754 4676 8764
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 3948 8370 4116 8372
rect 3948 8318 3950 8370
rect 4002 8318 4116 8370
rect 3948 8316 4116 8318
rect 3948 8306 4004 8316
rect 2380 8206 2382 8258
rect 2434 8206 2436 8258
rect 2380 8194 2436 8206
rect 3724 8258 3780 8270
rect 3724 8206 3726 8258
rect 3778 8206 3780 8258
rect 2716 8148 2772 8158
rect 3052 8148 3108 8158
rect 2716 8146 3108 8148
rect 2716 8094 2718 8146
rect 2770 8094 3054 8146
rect 3106 8094 3108 8146
rect 2716 8092 3108 8094
rect 2716 8082 2772 8092
rect 3052 8082 3108 8092
rect 2604 8034 2660 8046
rect 2604 7982 2606 8034
rect 2658 7982 2660 8034
rect 2604 7588 2660 7982
rect 3724 7700 3780 8206
rect 5068 8148 5124 8158
rect 3724 7634 3780 7644
rect 4956 8034 5012 8046
rect 4956 7982 4958 8034
rect 5010 7982 5012 8034
rect 4956 7700 5012 7982
rect 4956 7634 5012 7644
rect 2716 7588 2772 7598
rect 2604 7586 2772 7588
rect 2604 7534 2718 7586
rect 2770 7534 2772 7586
rect 2604 7532 2772 7534
rect 2716 7522 2772 7532
rect 4844 7364 4900 7374
rect 5068 7364 5124 8092
rect 4844 7362 5124 7364
rect 4844 7310 4846 7362
rect 4898 7310 5124 7362
rect 4844 7308 5124 7310
rect 5180 7364 5236 8876
rect 5516 8484 5572 20636
rect 5852 20242 5908 21980
rect 6412 21586 6468 22092
rect 6860 22146 6916 22158
rect 6860 22094 6862 22146
rect 6914 22094 6916 22146
rect 6860 21924 6916 22094
rect 6860 21858 6916 21868
rect 6412 21534 6414 21586
rect 6466 21534 6468 21586
rect 6412 21522 6468 21534
rect 6972 21586 7028 22318
rect 6972 21534 6974 21586
rect 7026 21534 7028 21586
rect 6972 21522 7028 21534
rect 7084 23492 7140 23502
rect 7084 22260 7140 23436
rect 7196 23154 7252 23166
rect 7196 23102 7198 23154
rect 7250 23102 7252 23154
rect 7196 22596 7252 23102
rect 7196 22530 7252 22540
rect 7308 22372 7364 23660
rect 7644 22594 7700 23774
rect 7868 23826 7924 24892
rect 7868 23774 7870 23826
rect 7922 23774 7924 23826
rect 7868 23762 7924 23774
rect 7980 25394 8036 26852
rect 7980 25342 7982 25394
rect 8034 25342 8036 25394
rect 7756 23714 7812 23726
rect 7756 23662 7758 23714
rect 7810 23662 7812 23714
rect 7756 23044 7812 23662
rect 7980 23492 8036 25342
rect 7980 23426 8036 23436
rect 8204 25282 8260 25294
rect 8204 25230 8206 25282
rect 8258 25230 8260 25282
rect 7980 23156 8036 23166
rect 7980 23062 8036 23100
rect 7756 22978 7812 22988
rect 8092 22930 8148 22942
rect 8092 22878 8094 22930
rect 8146 22878 8148 22930
rect 7644 22542 7646 22594
rect 7698 22542 7700 22594
rect 7644 22530 7700 22542
rect 7756 22596 7812 22606
rect 7812 22540 8036 22596
rect 7756 22530 7812 22540
rect 7084 21588 7140 22204
rect 7084 21522 7140 21532
rect 7196 22316 7364 22372
rect 7420 22370 7476 22382
rect 7420 22318 7422 22370
rect 7474 22318 7476 22370
rect 7196 20804 7252 22316
rect 7308 22148 7364 22158
rect 7308 22054 7364 22092
rect 7420 21588 7476 22318
rect 7980 22370 8036 22540
rect 7980 22318 7982 22370
rect 8034 22318 8036 22370
rect 7756 21698 7812 21710
rect 7756 21646 7758 21698
rect 7810 21646 7812 21698
rect 7532 21588 7588 21598
rect 7420 21586 7588 21588
rect 7420 21534 7534 21586
rect 7586 21534 7588 21586
rect 7420 21532 7588 21534
rect 7420 20916 7476 20926
rect 7420 20822 7476 20860
rect 6972 20748 7252 20804
rect 5852 20190 5854 20242
rect 5906 20190 5908 20242
rect 5852 20178 5908 20190
rect 6412 20580 6468 20590
rect 5628 20132 5684 20142
rect 5628 19458 5684 20076
rect 6412 20130 6468 20524
rect 6412 20078 6414 20130
rect 6466 20078 6468 20130
rect 6412 20066 6468 20078
rect 6300 20018 6356 20030
rect 6300 19966 6302 20018
rect 6354 19966 6356 20018
rect 6300 19460 6356 19966
rect 6524 20020 6580 20030
rect 6524 19926 6580 19964
rect 5628 19406 5630 19458
rect 5682 19406 5684 19458
rect 5628 19394 5684 19406
rect 5964 19404 6356 19460
rect 5964 19236 6020 19404
rect 5852 19234 6020 19236
rect 5852 19182 5966 19234
rect 6018 19182 6020 19234
rect 5852 19180 6020 19182
rect 5740 17668 5796 17678
rect 5740 17574 5796 17612
rect 5852 16772 5908 19180
rect 5964 19170 6020 19180
rect 6188 19236 6244 19246
rect 6188 19142 6244 19180
rect 5964 18564 6020 18574
rect 5964 17556 6020 18508
rect 5964 17554 6356 17556
rect 5964 17502 5966 17554
rect 6018 17502 6356 17554
rect 5964 17500 6356 17502
rect 5964 17490 6020 17500
rect 5852 16706 5908 16716
rect 6076 16324 6132 16334
rect 5852 16098 5908 16110
rect 5852 16046 5854 16098
rect 5906 16046 5908 16098
rect 5628 15986 5684 15998
rect 5628 15934 5630 15986
rect 5682 15934 5684 15986
rect 5628 15428 5684 15934
rect 5628 15148 5684 15372
rect 5852 15314 5908 16046
rect 6076 15540 6132 16268
rect 6300 16322 6356 17500
rect 6300 16270 6302 16322
rect 6354 16270 6356 16322
rect 6076 15446 6132 15484
rect 6188 15876 6244 15886
rect 5852 15262 5854 15314
rect 5906 15262 5908 15314
rect 5852 15204 5908 15262
rect 5628 15092 5796 15148
rect 5852 15138 5908 15148
rect 5740 14420 5796 15092
rect 6188 15090 6244 15820
rect 6300 15426 6356 16270
rect 6972 16324 7028 20748
rect 7084 20580 7140 20590
rect 7532 20580 7588 21532
rect 7644 21364 7700 21374
rect 7644 20914 7700 21308
rect 7644 20862 7646 20914
rect 7698 20862 7700 20914
rect 7644 20850 7700 20862
rect 7140 20524 7588 20580
rect 7756 20804 7812 21646
rect 7980 21700 8036 22318
rect 8092 22260 8148 22878
rect 8204 22708 8260 25230
rect 8316 24612 8372 24622
rect 8316 23940 8372 24556
rect 8428 23940 8484 23950
rect 8316 23884 8428 23940
rect 8428 23846 8484 23884
rect 9100 23828 9156 23838
rect 8540 23826 9156 23828
rect 8540 23774 9102 23826
rect 9154 23774 9156 23826
rect 8540 23772 9156 23774
rect 8428 23268 8484 23278
rect 8540 23268 8596 23772
rect 9100 23762 9156 23772
rect 8428 23266 8596 23268
rect 8428 23214 8430 23266
rect 8482 23214 8596 23266
rect 8428 23212 8596 23214
rect 8428 23202 8484 23212
rect 8316 22932 8372 22942
rect 8316 22838 8372 22876
rect 8204 22642 8260 22652
rect 8204 22484 8260 22494
rect 8204 22390 8260 22428
rect 8876 22260 8932 22270
rect 9212 22260 9268 27804
rect 9436 28532 9492 28542
rect 9436 27748 9492 28476
rect 10332 28532 10388 28812
rect 10444 28866 10500 29372
rect 10668 29362 10724 29372
rect 10444 28814 10446 28866
rect 10498 28814 10500 28866
rect 10444 28802 10500 28814
rect 10668 28756 10724 28766
rect 10668 28662 10724 28700
rect 10332 28466 10388 28476
rect 9772 28420 9828 28430
rect 9772 28418 10276 28420
rect 9772 28366 9774 28418
rect 9826 28366 10276 28418
rect 9772 28364 10276 28366
rect 9772 28354 9828 28364
rect 10220 27972 10276 28364
rect 10332 27972 10388 27982
rect 10220 27970 10388 27972
rect 10220 27918 10334 27970
rect 10386 27918 10388 27970
rect 10220 27916 10388 27918
rect 10332 27906 10388 27916
rect 10444 27860 10500 27870
rect 10444 27766 10500 27804
rect 8092 22204 8484 22260
rect 8428 21810 8484 22204
rect 8652 22258 9268 22260
rect 8652 22206 8878 22258
rect 8930 22206 9268 22258
rect 8652 22204 9268 22206
rect 8428 21758 8430 21810
rect 8482 21758 8484 21810
rect 8428 21746 8484 21758
rect 8540 22146 8596 22158
rect 8540 22094 8542 22146
rect 8594 22094 8596 22146
rect 7980 21634 8036 21644
rect 8204 21586 8260 21598
rect 8204 21534 8206 21586
rect 8258 21534 8260 21586
rect 7084 20486 7140 20524
rect 7756 19236 7812 20748
rect 7868 21474 7924 21486
rect 7868 21422 7870 21474
rect 7922 21422 7924 21474
rect 7868 20802 7924 21422
rect 7868 20750 7870 20802
rect 7922 20750 7924 20802
rect 7868 20738 7924 20750
rect 8204 20132 8260 21534
rect 8540 21364 8596 22094
rect 8652 21698 8708 22204
rect 8876 22194 8932 22204
rect 9212 22036 9268 22204
rect 9212 21970 9268 21980
rect 9324 27074 9380 27086
rect 9324 27022 9326 27074
rect 9378 27022 9380 27074
rect 8652 21646 8654 21698
rect 8706 21646 8708 21698
rect 8652 21634 8708 21646
rect 8764 21700 8820 21710
rect 8540 21298 8596 21308
rect 8652 20804 8708 20814
rect 8652 20710 8708 20748
rect 8316 20692 8372 20702
rect 8316 20598 8372 20636
rect 8652 20244 8708 20254
rect 8764 20244 8820 21644
rect 8876 21586 8932 21598
rect 8876 21534 8878 21586
rect 8930 21534 8932 21586
rect 8876 21028 8932 21534
rect 8876 20962 8932 20972
rect 8652 20242 8764 20244
rect 8652 20190 8654 20242
rect 8706 20190 8764 20242
rect 8652 20188 8764 20190
rect 8652 20178 8708 20188
rect 8764 20150 8820 20188
rect 8204 20066 8260 20076
rect 7756 19170 7812 19180
rect 8428 20018 8484 20030
rect 8428 19966 8430 20018
rect 8482 19966 8484 20018
rect 8428 19236 8484 19966
rect 9324 19460 9380 27022
rect 9436 19572 9492 27692
rect 10780 27636 10836 29372
rect 10892 28868 10948 29934
rect 11004 29988 11060 30156
rect 11228 30100 11284 30110
rect 11452 30100 11508 33182
rect 11788 32674 11844 35196
rect 11788 32622 11790 32674
rect 11842 32622 11844 32674
rect 11788 32610 11844 32622
rect 11900 38220 12012 38276
rect 11900 32004 11956 38220
rect 12012 38210 12068 38220
rect 12124 35812 12180 38612
rect 12236 38612 12292 38622
rect 12236 38518 12292 38556
rect 13132 38500 13188 38782
rect 13132 38434 13188 38444
rect 13580 38722 13636 38734
rect 13580 38670 13582 38722
rect 13634 38670 13636 38722
rect 12236 37938 12292 37950
rect 12236 37886 12238 37938
rect 12290 37886 12292 37938
rect 12236 37492 12292 37886
rect 12348 37940 12404 37950
rect 12348 37846 12404 37884
rect 12684 37938 12740 37950
rect 12684 37886 12686 37938
rect 12738 37886 12740 37938
rect 12236 37426 12292 37436
rect 12684 37268 12740 37886
rect 13468 37940 13524 37950
rect 13468 37846 13524 37884
rect 12796 37826 12852 37838
rect 12796 37774 12798 37826
rect 12850 37774 12852 37826
rect 12796 37716 12852 37774
rect 13020 37828 13076 37838
rect 13020 37734 13076 37772
rect 12796 37650 12852 37660
rect 13580 37716 13636 38670
rect 14700 38722 14756 38734
rect 14700 38670 14702 38722
rect 14754 38670 14756 38722
rect 13804 38612 13860 38622
rect 13804 38162 13860 38556
rect 13804 38110 13806 38162
rect 13858 38110 13860 38162
rect 13804 38098 13860 38110
rect 14700 38164 14756 38670
rect 14700 38098 14756 38108
rect 13916 38052 13972 38062
rect 14140 38052 14196 38062
rect 13972 37996 14084 38052
rect 13916 37958 13972 37996
rect 13692 37828 13748 37838
rect 13692 37734 13748 37772
rect 13468 37492 13524 37502
rect 13468 37398 13524 37436
rect 13580 37490 13636 37660
rect 13580 37438 13582 37490
rect 13634 37438 13636 37490
rect 13356 37268 13412 37278
rect 12684 37266 13412 37268
rect 12684 37214 13358 37266
rect 13410 37214 13412 37266
rect 12684 37212 13412 37214
rect 13356 36484 13412 37212
rect 13580 36484 13636 37438
rect 13916 37268 13972 37278
rect 13916 37174 13972 37212
rect 14028 36708 14084 37996
rect 14140 37958 14196 37996
rect 15036 37604 15092 38894
rect 16156 38164 16212 38174
rect 15932 38052 15988 38062
rect 15932 37958 15988 37996
rect 16156 38050 16212 38108
rect 16156 37998 16158 38050
rect 16210 37998 16212 38050
rect 16156 37986 16212 37998
rect 16380 38050 16436 39004
rect 16492 38994 16548 39004
rect 16604 38946 16660 38958
rect 16604 38894 16606 38946
rect 16658 38894 16660 38946
rect 16604 38836 16660 38894
rect 16604 38770 16660 38780
rect 16380 37998 16382 38050
rect 16434 37998 16436 38050
rect 16380 37986 16436 37998
rect 16492 38500 16548 38510
rect 16492 38164 16548 38444
rect 16268 37828 16324 37838
rect 16268 37734 16324 37772
rect 15036 37538 15092 37548
rect 14364 37268 14420 37278
rect 14364 37174 14420 37212
rect 16492 37266 16548 38108
rect 16492 37214 16494 37266
rect 16546 37214 16548 37266
rect 13916 36652 14084 36708
rect 13692 36484 13748 36494
rect 13580 36482 13748 36484
rect 13580 36430 13694 36482
rect 13746 36430 13748 36482
rect 13580 36428 13748 36430
rect 13356 36418 13412 36428
rect 13692 36418 13748 36428
rect 13468 36372 13524 36382
rect 13468 36278 13524 36316
rect 12572 36258 12628 36270
rect 12572 36206 12574 36258
rect 12626 36206 12628 36258
rect 12572 35812 12628 36206
rect 13804 36258 13860 36270
rect 13804 36206 13806 36258
rect 13858 36206 13860 36258
rect 13804 36036 13860 36206
rect 12124 35810 12628 35812
rect 12124 35758 12126 35810
rect 12178 35758 12628 35810
rect 12124 35756 12628 35758
rect 13244 35980 13860 36036
rect 12124 35746 12180 35756
rect 12012 35474 12068 35486
rect 12012 35422 12014 35474
rect 12066 35422 12068 35474
rect 12012 35028 12068 35422
rect 12012 34962 12068 34972
rect 12124 35140 12180 35150
rect 12124 35026 12180 35084
rect 12124 34974 12126 35026
rect 12178 34974 12180 35026
rect 11900 31948 12068 32004
rect 11788 31892 11844 31902
rect 12012 31892 12068 31948
rect 11844 31836 11956 31892
rect 11788 31826 11844 31836
rect 11564 31780 11620 31790
rect 11564 31686 11620 31724
rect 11788 31554 11844 31566
rect 11788 31502 11790 31554
rect 11842 31502 11844 31554
rect 11788 30436 11844 31502
rect 11228 30098 11508 30100
rect 11228 30046 11230 30098
rect 11282 30046 11508 30098
rect 11228 30044 11508 30046
rect 11564 30380 11844 30436
rect 11228 29988 11284 30044
rect 11004 29932 11172 29988
rect 11116 29652 11172 29932
rect 11228 29922 11284 29932
rect 11564 29764 11620 30380
rect 11788 30322 11844 30380
rect 11788 30270 11790 30322
rect 11842 30270 11844 30322
rect 11788 30258 11844 30270
rect 11676 30210 11732 30222
rect 11676 30158 11678 30210
rect 11730 30158 11732 30210
rect 11676 30100 11732 30158
rect 11900 30212 11956 31836
rect 12012 31666 12068 31836
rect 12124 31780 12180 34974
rect 12236 34132 12292 35756
rect 13244 35698 13300 35980
rect 13804 35812 13860 35822
rect 13244 35646 13246 35698
rect 13298 35646 13300 35698
rect 13244 35634 13300 35646
rect 13692 35756 13804 35812
rect 13692 35698 13748 35756
rect 13804 35746 13860 35756
rect 13692 35646 13694 35698
rect 13746 35646 13748 35698
rect 13692 35634 13748 35646
rect 12348 35588 12404 35598
rect 12348 35494 12404 35532
rect 13356 35586 13412 35598
rect 13356 35534 13358 35586
rect 13410 35534 13412 35586
rect 12460 34914 12516 34926
rect 12460 34862 12462 34914
rect 12514 34862 12516 34914
rect 12460 34468 12516 34862
rect 12908 34804 12964 34814
rect 13356 34804 13412 35534
rect 13468 34804 13524 34814
rect 13356 34802 13524 34804
rect 13356 34750 13470 34802
rect 13522 34750 13524 34802
rect 13356 34748 13524 34750
rect 12908 34710 12964 34748
rect 13468 34692 13524 34748
rect 13468 34636 13636 34692
rect 12460 34354 12516 34412
rect 12460 34302 12462 34354
rect 12514 34302 12516 34354
rect 12460 34290 12516 34302
rect 12796 34356 12852 34366
rect 12796 34262 12852 34300
rect 13468 34356 13524 34366
rect 12236 34076 12516 34132
rect 12124 31686 12180 31724
rect 12012 31614 12014 31666
rect 12066 31614 12068 31666
rect 12012 30324 12068 31614
rect 12012 30268 12292 30324
rect 11900 30156 12068 30212
rect 11676 30034 11732 30044
rect 12012 29988 12068 30156
rect 11564 29698 11620 29708
rect 11788 29932 12068 29988
rect 11340 29652 11396 29662
rect 11116 29596 11284 29652
rect 10892 28802 10948 28812
rect 11004 29426 11060 29438
rect 11004 29374 11006 29426
rect 11058 29374 11060 29426
rect 11004 28866 11060 29374
rect 11004 28814 11006 28866
rect 11058 28814 11060 28866
rect 11004 28802 11060 28814
rect 11116 29316 11172 29326
rect 10892 28642 10948 28654
rect 11116 28644 11172 29260
rect 11228 29316 11284 29596
rect 11340 29558 11396 29596
rect 11564 29538 11620 29550
rect 11564 29486 11566 29538
rect 11618 29486 11620 29538
rect 11564 29316 11620 29486
rect 11228 29260 11620 29316
rect 11228 28980 11284 29260
rect 11676 29204 11732 29214
rect 11676 29110 11732 29148
rect 11228 28924 11396 28980
rect 10892 28590 10894 28642
rect 10946 28590 10948 28642
rect 10892 28420 10948 28590
rect 10892 28354 10948 28364
rect 11004 28588 11172 28644
rect 11228 28756 11284 28766
rect 10892 27860 10948 27870
rect 11004 27860 11060 28588
rect 11228 28082 11284 28700
rect 11228 28030 11230 28082
rect 11282 28030 11284 28082
rect 11228 28018 11284 28030
rect 10892 27858 11060 27860
rect 10892 27806 10894 27858
rect 10946 27806 11060 27858
rect 10892 27804 11060 27806
rect 10892 27794 10948 27804
rect 11116 27636 11172 27646
rect 10780 27634 11172 27636
rect 10780 27582 11118 27634
rect 11170 27582 11172 27634
rect 10780 27580 11172 27582
rect 9772 27188 9828 27198
rect 9772 27094 9828 27132
rect 10444 27188 10500 27198
rect 10444 27094 10500 27132
rect 11116 27186 11172 27580
rect 11116 27134 11118 27186
rect 11170 27134 11172 27186
rect 11116 27122 11172 27134
rect 11340 26908 11396 28924
rect 11452 28868 11508 28878
rect 11508 28812 11620 28868
rect 11452 28802 11508 28812
rect 11564 28754 11620 28812
rect 11788 28866 11844 29932
rect 11788 28814 11790 28866
rect 11842 28814 11844 28866
rect 11788 28802 11844 28814
rect 11900 28980 11956 28990
rect 11564 28702 11566 28754
rect 11618 28702 11620 28754
rect 11564 28690 11620 28702
rect 11900 27186 11956 28924
rect 12124 28756 12180 28766
rect 12012 28644 12068 28654
rect 12012 28550 12068 28588
rect 12124 28642 12180 28700
rect 12124 28590 12126 28642
rect 12178 28590 12180 28642
rect 12124 28578 12180 28590
rect 11900 27134 11902 27186
rect 11954 27134 11956 27186
rect 11900 27122 11956 27134
rect 12236 27188 12292 30268
rect 12348 28532 12404 28542
rect 12348 28438 12404 28476
rect 12236 27122 12292 27132
rect 11564 27074 11620 27086
rect 11564 27022 11566 27074
rect 11618 27022 11620 27074
rect 11564 26908 11620 27022
rect 11116 26852 11396 26908
rect 11452 26852 11620 26908
rect 12460 26964 12516 34076
rect 13468 34130 13524 34300
rect 13580 34244 13636 34636
rect 13580 34178 13636 34188
rect 13468 34078 13470 34130
rect 13522 34078 13524 34130
rect 12796 33572 12852 33582
rect 12572 33236 12628 33246
rect 12572 33142 12628 33180
rect 12796 33234 12852 33516
rect 12796 33182 12798 33234
rect 12850 33182 12852 33234
rect 12796 33170 12852 33182
rect 12684 33122 12740 33134
rect 12684 33070 12686 33122
rect 12738 33070 12740 33122
rect 12572 31892 12628 31902
rect 12572 31798 12628 31836
rect 12684 31780 12740 33070
rect 12684 31714 12740 31724
rect 13468 31556 13524 34078
rect 13916 34130 13972 36652
rect 13916 34078 13918 34130
rect 13970 34078 13972 34130
rect 13916 33572 13972 34078
rect 13916 33506 13972 33516
rect 14028 36484 14084 36494
rect 14028 36370 14084 36428
rect 14028 36318 14030 36370
rect 14082 36318 14084 36370
rect 14028 33570 14084 36318
rect 14476 35812 14532 35822
rect 14476 35718 14532 35756
rect 14700 35812 14756 35822
rect 14700 35718 14756 35756
rect 14140 35700 14196 35710
rect 14140 35606 14196 35644
rect 14252 35698 14308 35710
rect 14252 35646 14254 35698
rect 14306 35646 14308 35698
rect 14252 35026 14308 35646
rect 14364 35588 14420 35598
rect 14364 35494 14420 35532
rect 14252 34974 14254 35026
rect 14306 34974 14308 35026
rect 14140 34914 14196 34926
rect 14140 34862 14142 34914
rect 14194 34862 14196 34914
rect 14140 34468 14196 34862
rect 14140 34402 14196 34412
rect 14140 34132 14196 34142
rect 14140 34038 14196 34076
rect 14252 33684 14308 34974
rect 14924 34916 14980 34926
rect 14924 34822 14980 34860
rect 14812 34804 14868 34814
rect 14812 34710 14868 34748
rect 14924 34692 14980 34702
rect 14700 34244 14756 34254
rect 14700 34150 14756 34188
rect 14588 34132 14644 34142
rect 14588 34038 14644 34076
rect 14028 33518 14030 33570
rect 14082 33518 14084 33570
rect 14028 33506 14084 33518
rect 14140 33628 14308 33684
rect 14140 33236 14196 33628
rect 14140 33170 14196 33180
rect 14252 33348 14308 33358
rect 14028 31892 14084 31902
rect 13580 31556 13636 31566
rect 13468 31500 13580 31556
rect 13468 28644 13524 28654
rect 13468 28550 13524 28588
rect 12460 26898 12516 26908
rect 13468 28420 13524 28430
rect 13468 27074 13524 28364
rect 13468 27022 13470 27074
rect 13522 27022 13524 27074
rect 10332 23044 10388 23054
rect 9884 22372 9940 22382
rect 9884 22278 9940 22316
rect 10332 22370 10388 22988
rect 10332 22318 10334 22370
rect 10386 22318 10388 22370
rect 10332 22306 10388 22318
rect 9996 22260 10052 22270
rect 9996 22166 10052 22204
rect 10108 22258 10164 22270
rect 10108 22206 10110 22258
rect 10162 22206 10164 22258
rect 9548 22036 9604 22046
rect 9604 21980 9716 22036
rect 9548 21970 9604 21980
rect 9548 21700 9604 21710
rect 9548 21606 9604 21644
rect 9548 21028 9604 21038
rect 9548 20130 9604 20972
rect 9660 20690 9716 21980
rect 10108 21924 10164 22206
rect 10780 22260 10836 22270
rect 10780 22166 10836 22204
rect 9884 21868 10164 21924
rect 9772 21698 9828 21710
rect 9772 21646 9774 21698
rect 9826 21646 9828 21698
rect 9772 21028 9828 21646
rect 9884 21474 9940 21868
rect 9884 21422 9886 21474
rect 9938 21422 9940 21474
rect 9884 21410 9940 21422
rect 10444 21812 10500 21822
rect 9828 20972 10164 21028
rect 9772 20962 9828 20972
rect 9660 20638 9662 20690
rect 9714 20638 9716 20690
rect 9660 20626 9716 20638
rect 10108 20690 10164 20972
rect 10444 20804 10500 21756
rect 10444 20710 10500 20748
rect 10108 20638 10110 20690
rect 10162 20638 10164 20690
rect 10108 20626 10164 20638
rect 10332 20580 10388 20590
rect 9548 20078 9550 20130
rect 9602 20078 9604 20130
rect 9548 20066 9604 20078
rect 9772 20244 9828 20254
rect 9772 20018 9828 20188
rect 9772 19966 9774 20018
rect 9826 19966 9828 20018
rect 9772 19954 9828 19966
rect 9996 19796 10052 19806
rect 9436 19506 9492 19516
rect 9884 19794 10052 19796
rect 9884 19742 9998 19794
rect 10050 19742 10052 19794
rect 9884 19740 10052 19742
rect 8428 19170 8484 19180
rect 8540 19404 9380 19460
rect 8540 17668 8596 19404
rect 9884 19348 9940 19740
rect 9996 19730 10052 19740
rect 10220 19794 10276 19806
rect 10220 19742 10222 19794
rect 10274 19742 10276 19794
rect 9100 19292 9940 19348
rect 9100 19236 9156 19292
rect 7644 17556 7700 17566
rect 7308 16994 7364 17006
rect 7308 16942 7310 16994
rect 7362 16942 7364 16994
rect 7308 16772 7364 16942
rect 7644 16996 7700 17500
rect 8428 17556 8484 17566
rect 8428 17462 8484 17500
rect 8540 17554 8596 17612
rect 8764 19234 9156 19236
rect 8764 19182 9102 19234
rect 9154 19182 9156 19234
rect 8764 19180 9156 19182
rect 8764 17666 8820 19180
rect 9100 19170 9156 19180
rect 9212 19124 9268 19134
rect 9212 19030 9268 19068
rect 10220 19124 10276 19742
rect 10220 19058 10276 19068
rect 8764 17614 8766 17666
rect 8818 17614 8820 17666
rect 8764 17602 8820 17614
rect 8540 17502 8542 17554
rect 8594 17502 8596 17554
rect 7644 16994 7924 16996
rect 7644 16942 7646 16994
rect 7698 16942 7924 16994
rect 7644 16940 7924 16942
rect 7644 16930 7700 16940
rect 7308 16706 7364 16716
rect 7756 16772 7812 16782
rect 6972 16258 7028 16268
rect 7644 16324 7700 16334
rect 6748 16100 6804 16110
rect 7084 16100 7140 16110
rect 6748 16098 7140 16100
rect 6748 16046 6750 16098
rect 6802 16046 7086 16098
rect 7138 16046 7140 16098
rect 6748 16044 7140 16046
rect 6748 16034 6804 16044
rect 7084 16034 7140 16044
rect 7644 15986 7700 16268
rect 7756 16322 7812 16716
rect 7756 16270 7758 16322
rect 7810 16270 7812 16322
rect 7756 16258 7812 16270
rect 7644 15934 7646 15986
rect 7698 15934 7700 15986
rect 7644 15922 7700 15934
rect 7420 15876 7476 15886
rect 7420 15782 7476 15820
rect 7308 15540 7364 15550
rect 6300 15374 6302 15426
rect 6354 15374 6356 15426
rect 6300 15362 6356 15374
rect 7196 15484 7308 15540
rect 7196 15426 7252 15484
rect 7308 15474 7364 15484
rect 7756 15540 7812 15550
rect 7868 15540 7924 16940
rect 7756 15538 7924 15540
rect 7756 15486 7758 15538
rect 7810 15486 7924 15538
rect 7756 15484 7924 15486
rect 7756 15474 7812 15484
rect 7196 15374 7198 15426
rect 7250 15374 7252 15426
rect 6860 15316 6916 15354
rect 6636 15260 6860 15316
rect 6188 15038 6190 15090
rect 6242 15038 6244 15090
rect 6188 15026 6244 15038
rect 6524 15204 6580 15214
rect 5852 14420 5908 14430
rect 5740 14418 5908 14420
rect 5740 14366 5854 14418
rect 5906 14366 5908 14418
rect 5740 14364 5908 14366
rect 5852 14354 5908 14364
rect 6188 14418 6244 14430
rect 6188 14366 6190 14418
rect 6242 14366 6244 14418
rect 6188 14196 6244 14366
rect 6524 14418 6580 15148
rect 6524 14366 6526 14418
rect 6578 14366 6580 14418
rect 6524 14354 6580 14366
rect 6636 14196 6692 15260
rect 6860 15250 6916 15260
rect 6972 15314 7028 15326
rect 6972 15262 6974 15314
rect 7026 15262 7028 15314
rect 6188 14140 6692 14196
rect 6748 15092 6804 15102
rect 6748 14530 6804 15036
rect 6748 14478 6750 14530
rect 6802 14478 6804 14530
rect 5628 13636 5684 13646
rect 5628 12402 5684 13580
rect 5628 12350 5630 12402
rect 5682 12350 5684 12402
rect 5628 12338 5684 12350
rect 6188 12404 6244 14140
rect 6636 12404 6692 12414
rect 6748 12404 6804 14478
rect 6188 12348 6580 12404
rect 6300 12178 6356 12190
rect 6300 12126 6302 12178
rect 6354 12126 6356 12178
rect 5852 11954 5908 11966
rect 5852 11902 5854 11954
rect 5906 11902 5908 11954
rect 5852 11394 5908 11902
rect 6076 11956 6132 11966
rect 6300 11956 6356 12126
rect 6076 11954 6468 11956
rect 6076 11902 6078 11954
rect 6130 11902 6468 11954
rect 6076 11900 6468 11902
rect 6076 11890 6132 11900
rect 5852 11342 5854 11394
rect 5906 11342 5908 11394
rect 5852 11330 5908 11342
rect 5964 11620 6020 11630
rect 5964 11282 6020 11564
rect 6412 11618 6468 11900
rect 6412 11566 6414 11618
rect 6466 11566 6468 11618
rect 6412 11554 6468 11566
rect 6524 11396 6580 12348
rect 6636 12402 6804 12404
rect 6636 12350 6638 12402
rect 6690 12350 6804 12402
rect 6636 12348 6804 12350
rect 6636 12338 6692 12348
rect 6748 11620 6804 11630
rect 6748 11396 6804 11564
rect 5964 11230 5966 11282
rect 6018 11230 6020 11282
rect 5964 11218 6020 11230
rect 6412 11340 6580 11396
rect 6636 11394 6804 11396
rect 6636 11342 6750 11394
rect 6802 11342 6804 11394
rect 6636 11340 6804 11342
rect 6188 11172 6244 11182
rect 6188 11078 6244 11116
rect 5516 8418 5572 8428
rect 5964 9044 6020 9054
rect 5628 8148 5684 8158
rect 5628 8054 5684 8092
rect 5964 8146 6020 8988
rect 6300 9044 6356 9054
rect 6412 9044 6468 11340
rect 6524 11170 6580 11182
rect 6524 11118 6526 11170
rect 6578 11118 6580 11170
rect 6524 10836 6580 11118
rect 6524 10770 6580 10780
rect 6356 8988 6468 9044
rect 6300 8978 6356 8988
rect 5964 8094 5966 8146
rect 6018 8094 6020 8146
rect 5964 8082 6020 8094
rect 6636 7698 6692 11340
rect 6748 11330 6804 11340
rect 6972 8820 7028 15262
rect 7196 15204 7252 15374
rect 7196 15138 7252 15148
rect 7308 15314 7364 15326
rect 7308 15262 7310 15314
rect 7362 15262 7364 15314
rect 7308 14532 7364 15262
rect 8540 15314 8596 17502
rect 10108 16884 10164 16894
rect 10332 16884 10388 20524
rect 11116 20356 11172 26852
rect 11340 24052 11396 24062
rect 11452 24052 11508 26852
rect 13020 26290 13076 26302
rect 13020 26238 13022 26290
rect 13074 26238 13076 26290
rect 13020 26180 13076 26238
rect 13020 26114 13076 26124
rect 13468 25618 13524 27022
rect 13580 26908 13636 31500
rect 13804 31220 13860 31230
rect 14028 31220 14084 31836
rect 14252 31778 14308 33292
rect 14924 33346 14980 34636
rect 16156 34692 16212 34702
rect 16156 34242 16212 34636
rect 16156 34190 16158 34242
rect 16210 34190 16212 34242
rect 16156 34178 16212 34190
rect 15036 34132 15092 34142
rect 15036 33458 15092 34076
rect 15596 34132 15652 34142
rect 15596 34038 15652 34076
rect 15036 33406 15038 33458
rect 15090 33406 15092 33458
rect 15036 33394 15092 33406
rect 15932 34018 15988 34030
rect 15932 33966 15934 34018
rect 15986 33966 15988 34018
rect 14924 33294 14926 33346
rect 14978 33294 14980 33346
rect 14924 33282 14980 33294
rect 15708 33348 15764 33358
rect 15708 33254 15764 33292
rect 14252 31726 14254 31778
rect 14306 31726 14308 31778
rect 14252 31714 14308 31726
rect 14588 33124 14644 33134
rect 13692 30996 13748 31006
rect 13692 30098 13748 30940
rect 13804 30994 13860 31164
rect 13804 30942 13806 30994
rect 13858 30942 13860 30994
rect 13804 30930 13860 30942
rect 13916 31218 14084 31220
rect 13916 31166 14030 31218
rect 14082 31166 14084 31218
rect 13916 31164 14084 31166
rect 13916 30548 13972 31164
rect 14028 31154 14084 31164
rect 13916 30492 14196 30548
rect 13916 30434 13972 30492
rect 13916 30382 13918 30434
rect 13970 30382 13972 30434
rect 13916 30370 13972 30382
rect 13692 30046 13694 30098
rect 13746 30046 13748 30098
rect 13692 30034 13748 30046
rect 14028 30324 14084 30334
rect 13804 29988 13860 29998
rect 13804 29316 13860 29932
rect 13916 29652 13972 29662
rect 14028 29652 14084 30268
rect 13916 29650 14084 29652
rect 13916 29598 13918 29650
rect 13970 29598 14084 29650
rect 13916 29596 14084 29598
rect 14140 29652 14196 30492
rect 14364 30212 14420 30222
rect 14364 30118 14420 30156
rect 14476 30100 14532 30110
rect 14476 30006 14532 30044
rect 14252 29988 14308 29998
rect 14252 29894 14308 29932
rect 14476 29652 14532 29662
rect 14140 29650 14532 29652
rect 14140 29598 14478 29650
rect 14530 29598 14532 29650
rect 14140 29596 14532 29598
rect 13916 29586 13972 29596
rect 14476 29586 14532 29596
rect 14028 29428 14084 29438
rect 14252 29428 14308 29438
rect 14028 29426 14308 29428
rect 14028 29374 14030 29426
rect 14082 29374 14254 29426
rect 14306 29374 14308 29426
rect 14028 29372 14308 29374
rect 14028 29362 14084 29372
rect 14252 29362 14308 29372
rect 14364 29428 14420 29438
rect 13804 29250 13860 29260
rect 13692 29204 13748 29214
rect 13692 28754 13748 29148
rect 13916 29204 13972 29214
rect 13916 29202 14084 29204
rect 13916 29150 13918 29202
rect 13970 29150 14084 29202
rect 13916 29148 14084 29150
rect 13916 29138 13972 29148
rect 13692 28702 13694 28754
rect 13746 28702 13748 28754
rect 13692 28690 13748 28702
rect 13916 28644 13972 28654
rect 13916 28550 13972 28588
rect 14028 28642 14084 29148
rect 14028 28590 14030 28642
rect 14082 28590 14084 28642
rect 14028 28578 14084 28590
rect 14364 29092 14420 29372
rect 14364 28642 14420 29036
rect 14588 29426 14644 33068
rect 15596 33124 15652 33134
rect 15820 33124 15876 33134
rect 15596 33030 15652 33068
rect 15708 33122 15876 33124
rect 15708 33070 15822 33122
rect 15874 33070 15876 33122
rect 15708 33068 15876 33070
rect 15708 32788 15764 33068
rect 15820 33058 15876 33068
rect 15372 32732 15764 32788
rect 14924 31780 14980 31790
rect 14812 31668 14868 31678
rect 14812 31574 14868 31612
rect 14700 31556 14756 31566
rect 14700 31462 14756 31500
rect 14924 30324 14980 31724
rect 15372 31220 15428 32732
rect 15932 32676 15988 33966
rect 16268 33348 16324 33358
rect 16492 33348 16548 37214
rect 16604 37938 16660 37950
rect 16604 37886 16606 37938
rect 16658 37886 16660 37938
rect 16604 35924 16660 37886
rect 16716 37492 16772 39452
rect 17724 38948 17780 39676
rect 18620 39732 18676 39742
rect 18620 39638 18676 39676
rect 21308 39730 21364 39742
rect 21308 39678 21310 39730
rect 21362 39678 21364 39730
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 17500 38946 17780 38948
rect 17500 38894 17726 38946
rect 17778 38894 17780 38946
rect 17500 38892 17780 38894
rect 17388 38834 17444 38846
rect 17388 38782 17390 38834
rect 17442 38782 17444 38834
rect 16716 37426 16772 37436
rect 16828 38388 16884 38398
rect 16828 37604 16884 38332
rect 17164 38276 17220 38286
rect 17164 38162 17220 38220
rect 17164 38110 17166 38162
rect 17218 38110 17220 38162
rect 17164 38098 17220 38110
rect 17388 38164 17444 38782
rect 17388 38098 17444 38108
rect 17500 38052 17556 38892
rect 17724 38882 17780 38892
rect 18284 38946 18340 38958
rect 18284 38894 18286 38946
rect 18338 38894 18340 38946
rect 18060 38834 18116 38846
rect 18060 38782 18062 38834
rect 18114 38782 18116 38834
rect 17612 38722 17668 38734
rect 17612 38670 17614 38722
rect 17666 38670 17668 38722
rect 17612 38668 17668 38670
rect 18060 38668 18116 38782
rect 18172 38836 18228 38846
rect 18284 38836 18340 38894
rect 21308 38948 21364 39678
rect 24220 39620 24276 39630
rect 24668 39620 24724 39630
rect 24220 39618 24724 39620
rect 24220 39566 24222 39618
rect 24274 39566 24670 39618
rect 24722 39566 24724 39618
rect 24220 39564 24724 39566
rect 24220 39554 24276 39564
rect 23436 39508 23492 39518
rect 18396 38836 18452 38846
rect 18732 38836 18788 38846
rect 20188 38836 20244 38846
rect 20300 38836 20356 38846
rect 18284 38780 18396 38836
rect 18452 38780 18676 38836
rect 18172 38742 18228 38780
rect 18396 38770 18452 38780
rect 18620 38668 18676 38780
rect 18732 38834 19908 38836
rect 18732 38782 18734 38834
rect 18786 38782 19908 38834
rect 18732 38780 19908 38782
rect 18732 38770 18788 38780
rect 17612 38612 18004 38668
rect 18060 38612 18452 38668
rect 18620 38612 18788 38668
rect 17836 38276 17892 38286
rect 17948 38276 18004 38612
rect 18172 38276 18228 38286
rect 17948 38274 18228 38276
rect 17948 38222 18174 38274
rect 18226 38222 18228 38274
rect 17948 38220 18228 38222
rect 17612 38052 17668 38062
rect 17500 38050 17668 38052
rect 17500 37998 17614 38050
rect 17666 37998 17668 38050
rect 17500 37996 17668 37998
rect 17612 37986 17668 37996
rect 16828 37490 16884 37548
rect 16828 37438 16830 37490
rect 16882 37438 16884 37490
rect 16604 33908 16660 35868
rect 16604 33842 16660 33852
rect 16828 33572 16884 37438
rect 17388 37828 17444 37838
rect 17388 37378 17444 37772
rect 17836 37604 17892 38220
rect 18172 38210 18228 38220
rect 18396 38050 18452 38612
rect 18396 37998 18398 38050
rect 18450 37998 18452 38050
rect 18172 37940 18228 37950
rect 17724 37548 18116 37604
rect 17500 37492 17556 37502
rect 17500 37398 17556 37436
rect 17388 37326 17390 37378
rect 17442 37326 17444 37378
rect 17388 37314 17444 37326
rect 17612 37380 17668 37390
rect 17612 37286 17668 37324
rect 17724 36594 17780 37548
rect 18060 37490 18116 37548
rect 18060 37438 18062 37490
rect 18114 37438 18116 37490
rect 18060 37426 18116 37438
rect 18172 37490 18228 37884
rect 18172 37438 18174 37490
rect 18226 37438 18228 37490
rect 18172 37426 18228 37438
rect 18060 37268 18116 37278
rect 18116 37212 18228 37268
rect 18060 37202 18116 37212
rect 17724 36542 17726 36594
rect 17778 36542 17780 36594
rect 17724 36530 17780 36542
rect 17500 35364 17556 35374
rect 17500 35026 17556 35308
rect 17500 34974 17502 35026
rect 17554 34974 17556 35026
rect 17500 34962 17556 34974
rect 17276 34916 17332 34926
rect 17276 34822 17332 34860
rect 17948 34916 18004 34954
rect 17948 34850 18004 34860
rect 17836 34802 17892 34814
rect 17836 34750 17838 34802
rect 17890 34750 17892 34802
rect 16940 34692 16996 34702
rect 17612 34692 17668 34702
rect 17836 34692 17892 34750
rect 16940 34690 17332 34692
rect 16940 34638 16942 34690
rect 16994 34638 17332 34690
rect 16940 34636 17332 34638
rect 16940 34626 16996 34636
rect 17276 34130 17332 34636
rect 17276 34078 17278 34130
rect 17330 34078 17332 34130
rect 17276 34066 17332 34078
rect 17668 34636 17892 34692
rect 17612 34354 17668 34636
rect 17612 34302 17614 34354
rect 17666 34302 17668 34354
rect 17500 33906 17556 33918
rect 17500 33854 17502 33906
rect 17554 33854 17556 33906
rect 16828 33516 17220 33572
rect 16940 33348 16996 33358
rect 16268 33346 16548 33348
rect 16268 33294 16270 33346
rect 16322 33294 16548 33346
rect 16268 33292 16548 33294
rect 16828 33346 16996 33348
rect 16828 33294 16942 33346
rect 16994 33294 16996 33346
rect 16828 33292 16996 33294
rect 16268 33282 16324 33292
rect 16716 33124 16772 33134
rect 16828 33124 16884 33292
rect 16940 33282 16996 33292
rect 16716 33122 16884 33124
rect 16716 33070 16718 33122
rect 16770 33070 16884 33122
rect 16716 33068 16884 33070
rect 15932 32620 16436 32676
rect 15372 31154 15428 31164
rect 15484 32562 15540 32574
rect 15484 32510 15486 32562
rect 15538 32510 15540 32562
rect 15484 32452 15540 32510
rect 15932 32452 15988 32462
rect 15484 32450 15988 32452
rect 15484 32398 15934 32450
rect 15986 32398 15988 32450
rect 15484 32396 15988 32398
rect 14924 30210 14980 30268
rect 14924 30158 14926 30210
rect 14978 30158 14980 30210
rect 14924 30146 14980 30158
rect 14588 29374 14590 29426
rect 14642 29374 14644 29426
rect 14588 28980 14644 29374
rect 14588 28914 14644 28924
rect 14364 28590 14366 28642
rect 14418 28590 14420 28642
rect 14364 28578 14420 28590
rect 14700 28644 14756 28654
rect 14812 28644 14868 28654
rect 14756 28642 14868 28644
rect 14756 28590 14814 28642
rect 14866 28590 14868 28642
rect 14756 28588 14868 28590
rect 13804 28532 13860 28542
rect 13804 26962 13860 28476
rect 13804 26910 13806 26962
rect 13858 26910 13860 26962
rect 13580 26852 13748 26908
rect 13468 25566 13470 25618
rect 13522 25566 13524 25618
rect 13468 25554 13524 25566
rect 11340 24050 11508 24052
rect 11340 23998 11342 24050
rect 11394 23998 11508 24050
rect 11340 23996 11508 23998
rect 12796 24052 12852 24062
rect 11340 21812 11396 23996
rect 12796 23958 12852 23996
rect 11900 23940 11956 23950
rect 11900 23846 11956 23884
rect 13692 23826 13748 26852
rect 13692 23774 13694 23826
rect 13746 23774 13748 23826
rect 13692 23762 13748 23774
rect 13804 24052 13860 26910
rect 14028 28418 14084 28430
rect 14028 28366 14030 28418
rect 14082 28366 14084 28418
rect 14028 25620 14084 28366
rect 14028 25554 14084 25564
rect 14252 26964 14308 26974
rect 12908 23716 12964 23726
rect 12908 23622 12964 23660
rect 12460 23042 12516 23054
rect 12460 22990 12462 23042
rect 12514 22990 12516 23042
rect 11564 22932 11620 22942
rect 11340 21746 11396 21756
rect 11452 22036 11508 22046
rect 11228 20580 11284 20590
rect 11228 20578 11396 20580
rect 11228 20526 11230 20578
rect 11282 20526 11396 20578
rect 11228 20524 11396 20526
rect 11228 20514 11284 20524
rect 11116 20300 11284 20356
rect 10780 20132 10836 20142
rect 10780 20038 10836 20076
rect 11116 19236 11172 19246
rect 11116 19142 11172 19180
rect 10108 16882 10276 16884
rect 10108 16830 10110 16882
rect 10162 16830 10276 16882
rect 10108 16828 10276 16830
rect 10108 16818 10164 16828
rect 9884 16660 9940 16670
rect 9772 16212 9828 16222
rect 9212 16098 9268 16110
rect 9212 16046 9214 16098
rect 9266 16046 9268 16098
rect 8988 15428 9044 15438
rect 8988 15334 9044 15372
rect 8540 15262 8542 15314
rect 8594 15262 8596 15314
rect 8540 15250 8596 15262
rect 9212 15316 9268 16046
rect 9772 16098 9828 16156
rect 9884 16210 9940 16604
rect 9884 16158 9886 16210
rect 9938 16158 9940 16210
rect 9884 16146 9940 16158
rect 9772 16046 9774 16098
rect 9826 16046 9828 16098
rect 9772 16034 9828 16046
rect 9212 15250 9268 15260
rect 10220 15540 10276 16828
rect 10332 16818 10388 16828
rect 10444 17108 10500 17118
rect 10444 16882 10500 17052
rect 10556 16996 10612 17006
rect 11116 16996 11172 17006
rect 10556 16994 11172 16996
rect 10556 16942 10558 16994
rect 10610 16942 11118 16994
rect 11170 16942 11172 16994
rect 10556 16940 11172 16942
rect 10556 16930 10612 16940
rect 11116 16930 11172 16940
rect 10444 16830 10446 16882
rect 10498 16830 10500 16882
rect 10444 16818 10500 16830
rect 11228 16770 11284 20300
rect 11340 20132 11396 20524
rect 11340 20066 11396 20076
rect 11228 16718 11230 16770
rect 11282 16718 11284 16770
rect 11228 16706 11284 16718
rect 10892 16660 10948 16670
rect 10892 16566 10948 16604
rect 10444 16212 10500 16222
rect 10444 16118 10500 16156
rect 8092 15202 8148 15214
rect 8092 15150 8094 15202
rect 8146 15150 8148 15202
rect 8092 15148 8148 15150
rect 7196 13524 7252 13534
rect 7308 13524 7364 14476
rect 7252 13468 7364 13524
rect 7980 15092 8148 15148
rect 10108 15204 10164 15242
rect 10108 15138 10164 15148
rect 7196 13074 7252 13468
rect 7196 13022 7198 13074
rect 7250 13022 7252 13074
rect 7196 13010 7252 13022
rect 7308 12740 7364 12750
rect 7308 12738 7476 12740
rect 7308 12686 7310 12738
rect 7362 12686 7476 12738
rect 7308 12684 7476 12686
rect 7308 12674 7364 12684
rect 7308 11954 7364 11966
rect 7308 11902 7310 11954
rect 7362 11902 7364 11954
rect 7308 11506 7364 11902
rect 7420 11620 7476 12684
rect 7980 12404 8036 15092
rect 8204 13972 8260 13982
rect 8092 13524 8148 13534
rect 8092 12962 8148 13468
rect 8092 12910 8094 12962
rect 8146 12910 8148 12962
rect 8092 12898 8148 12910
rect 8204 12850 8260 13916
rect 9660 13972 9716 13982
rect 9660 13878 9716 13916
rect 8204 12798 8206 12850
rect 8258 12798 8260 12850
rect 8204 12786 8260 12798
rect 9548 13634 9604 13646
rect 9548 13582 9550 13634
rect 9602 13582 9604 13634
rect 9548 13524 9604 13582
rect 8428 12740 8484 12750
rect 8428 12738 8820 12740
rect 8428 12686 8430 12738
rect 8482 12686 8820 12738
rect 8428 12684 8820 12686
rect 8428 12674 8484 12684
rect 8092 12404 8148 12414
rect 7980 12402 8148 12404
rect 7980 12350 8094 12402
rect 8146 12350 8148 12402
rect 7980 12348 8148 12350
rect 8092 12338 8148 12348
rect 8764 12402 8820 12684
rect 8764 12350 8766 12402
rect 8818 12350 8820 12402
rect 8764 12338 8820 12350
rect 9548 12292 9604 13468
rect 9324 12236 9604 12292
rect 7756 12180 7812 12190
rect 7644 12178 7812 12180
rect 7644 12126 7758 12178
rect 7810 12126 7812 12178
rect 7644 12124 7812 12126
rect 7644 11954 7700 12124
rect 7756 12114 7812 12124
rect 8092 12180 8148 12190
rect 8204 12180 8260 12190
rect 8092 12178 8204 12180
rect 8092 12126 8094 12178
rect 8146 12126 8204 12178
rect 8092 12124 8204 12126
rect 8092 12114 8148 12124
rect 7644 11902 7646 11954
rect 7698 11902 7700 11954
rect 7644 11890 7700 11902
rect 7420 11618 7924 11620
rect 7420 11566 7422 11618
rect 7474 11566 7924 11618
rect 7420 11564 7924 11566
rect 7420 11554 7476 11564
rect 7308 11454 7310 11506
rect 7362 11454 7364 11506
rect 7308 11442 7364 11454
rect 7084 11172 7140 11182
rect 7084 10834 7140 11116
rect 7196 11170 7252 11182
rect 7196 11118 7198 11170
rect 7250 11118 7252 11170
rect 7196 11060 7252 11118
rect 7196 11004 7700 11060
rect 7084 10782 7086 10834
rect 7138 10782 7140 10834
rect 7084 10770 7140 10782
rect 7308 10836 7364 10846
rect 7308 10742 7364 10780
rect 7532 10610 7588 10622
rect 7532 10558 7534 10610
rect 7586 10558 7588 10610
rect 7420 10500 7476 10510
rect 7420 10406 7476 10444
rect 7532 10052 7588 10558
rect 7644 10500 7700 11004
rect 7868 10722 7924 11564
rect 8092 11282 8148 11294
rect 8092 11230 8094 11282
rect 8146 11230 8148 11282
rect 8092 11172 8148 11230
rect 8092 11106 8148 11116
rect 8204 10834 8260 12124
rect 8204 10782 8206 10834
rect 8258 10782 8260 10834
rect 8204 10770 8260 10782
rect 8316 12178 8372 12190
rect 8316 12126 8318 12178
rect 8370 12126 8372 12178
rect 7868 10670 7870 10722
rect 7922 10670 7924 10722
rect 7868 10658 7924 10670
rect 7980 10722 8036 10734
rect 7980 10670 7982 10722
rect 8034 10670 8036 10722
rect 7980 10500 8036 10670
rect 7644 10444 8036 10500
rect 7980 10276 8036 10444
rect 7532 9986 7588 9996
rect 7868 10220 8036 10276
rect 8316 10500 8372 12126
rect 6972 8754 7028 8764
rect 6636 7646 6638 7698
rect 6690 7646 6692 7698
rect 6636 7634 6692 7646
rect 6748 7476 6804 7486
rect 7308 7476 7364 7486
rect 6748 7474 7364 7476
rect 6748 7422 6750 7474
rect 6802 7422 7310 7474
rect 7362 7422 7364 7474
rect 6748 7420 7364 7422
rect 5292 7364 5348 7374
rect 5180 7362 5348 7364
rect 5180 7310 5294 7362
rect 5346 7310 5348 7362
rect 5180 7308 5348 7310
rect 4844 7298 4900 7308
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4956 6468 5012 6478
rect 4956 6130 5012 6412
rect 5292 6468 5348 7308
rect 5292 6402 5348 6412
rect 5404 6804 5460 6814
rect 4956 6078 4958 6130
rect 5010 6078 5012 6130
rect 4956 6066 5012 6078
rect 5404 6130 5460 6748
rect 6300 6692 6356 6702
rect 6188 6636 6300 6692
rect 5404 6078 5406 6130
rect 5458 6078 5460 6130
rect 5404 6066 5460 6078
rect 5628 6580 5684 6590
rect 5628 6020 5684 6524
rect 5516 6018 5684 6020
rect 5516 5966 5630 6018
rect 5682 5966 5684 6018
rect 5516 5964 5684 5966
rect 4956 5908 5012 5918
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4732 5236 4788 5246
rect 4732 5142 4788 5180
rect 2604 5012 2660 5022
rect 2604 4918 2660 4956
rect 3948 4564 4004 4574
rect 3948 4470 4004 4508
rect 4956 4562 5012 5852
rect 5516 5236 5572 5964
rect 5628 5954 5684 5964
rect 5740 6020 5796 6030
rect 5740 5926 5796 5964
rect 6076 5908 6132 5918
rect 6076 5814 6132 5852
rect 5852 5796 5908 5806
rect 5516 5170 5572 5180
rect 5628 5572 5684 5582
rect 5628 5234 5684 5516
rect 5628 5182 5630 5234
rect 5682 5182 5684 5234
rect 5628 5170 5684 5182
rect 4956 4510 4958 4562
rect 5010 4510 5012 4562
rect 4956 4498 5012 4510
rect 5852 4562 5908 5740
rect 6076 5684 6132 5694
rect 5852 4510 5854 4562
rect 5906 4510 5908 4562
rect 5852 4498 5908 4510
rect 5964 5012 6020 5022
rect 5964 4562 6020 4956
rect 5964 4510 5966 4562
rect 6018 4510 6020 4562
rect 5964 4498 6020 4510
rect 4732 4340 4788 4350
rect 4732 4246 4788 4284
rect 5516 4340 5572 4350
rect 6076 4340 6132 5628
rect 3836 4226 3892 4238
rect 3836 4174 3838 4226
rect 3890 4174 3892 4226
rect 1820 3332 2100 3388
rect 3164 3444 3220 3454
rect 3388 3444 3444 3454
rect 3164 3442 3444 3444
rect 3164 3390 3166 3442
rect 3218 3390 3390 3442
rect 3442 3390 3444 3442
rect 3164 3388 3444 3390
rect 1820 800 1876 3332
rect 3164 800 3220 3388
rect 3388 3378 3444 3388
rect 3724 3444 3780 3454
rect 3836 3444 3892 4174
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 3724 3442 3892 3444
rect 3724 3390 3726 3442
rect 3778 3390 3892 3442
rect 3724 3388 3892 3390
rect 5068 3556 5124 3566
rect 5068 3388 5124 3500
rect 3724 3378 3780 3388
rect 4956 3332 5124 3388
rect 5516 3442 5572 4284
rect 5852 4284 6132 4340
rect 5740 3556 5796 3566
rect 5740 3462 5796 3500
rect 5516 3390 5518 3442
rect 5570 3390 5572 3442
rect 5516 3378 5572 3390
rect 4956 2212 5012 3332
rect 4508 2156 5012 2212
rect 4508 800 4564 2156
rect 5852 800 5908 4284
rect 6076 4116 6132 4126
rect 6188 4116 6244 6636
rect 6300 6626 6356 6636
rect 6748 6580 6804 7420
rect 7308 7410 7364 7420
rect 7308 7250 7364 7262
rect 7308 7198 7310 7250
rect 7362 7198 7364 7250
rect 7196 6916 7252 6926
rect 6860 6804 6916 6814
rect 6860 6710 6916 6748
rect 7196 6690 7252 6860
rect 7196 6638 7198 6690
rect 7250 6638 7252 6690
rect 7196 6626 7252 6638
rect 6748 6514 6804 6524
rect 7308 5796 7364 7198
rect 7644 7250 7700 7262
rect 7644 7198 7646 7250
rect 7698 7198 7700 7250
rect 7644 6020 7700 7198
rect 7756 6580 7812 6590
rect 7756 6486 7812 6524
rect 7868 6468 7924 10220
rect 8316 9714 8372 10444
rect 8540 12178 8596 12190
rect 8540 12126 8542 12178
rect 8594 12126 8596 12178
rect 8540 9826 8596 12126
rect 8876 12180 8932 12190
rect 8876 12086 8932 12124
rect 8540 9774 8542 9826
rect 8594 9774 8596 9826
rect 8540 9762 8596 9774
rect 8652 11394 8708 11406
rect 8652 11342 8654 11394
rect 8706 11342 8708 11394
rect 8652 10052 8708 11342
rect 8316 9662 8318 9714
rect 8370 9662 8372 9714
rect 8316 9650 8372 9662
rect 8652 9268 8708 9996
rect 8652 9202 8708 9212
rect 9212 9492 9268 9502
rect 8876 8820 8932 8830
rect 8428 8372 8484 8382
rect 8092 7588 8148 7598
rect 8092 7494 8148 7532
rect 7980 7474 8036 7486
rect 7980 7422 7982 7474
rect 8034 7422 8036 7474
rect 7980 6804 8036 7422
rect 7980 6738 8036 6748
rect 8092 7250 8148 7262
rect 8092 7198 8094 7250
rect 8146 7198 8148 7250
rect 8092 6692 8148 7198
rect 8092 6626 8148 6636
rect 8428 6916 8484 8316
rect 8876 8146 8932 8764
rect 8876 8094 8878 8146
rect 8930 8094 8932 8146
rect 8876 8036 8932 8094
rect 8876 7970 8932 7980
rect 8988 8034 9044 8046
rect 8988 7982 8990 8034
rect 9042 7982 9044 8034
rect 8428 6578 8484 6860
rect 8652 7588 8708 7598
rect 8652 7362 8708 7532
rect 8652 7310 8654 7362
rect 8706 7310 8708 7362
rect 8652 6916 8708 7310
rect 8652 6850 8708 6860
rect 8988 6914 9044 7982
rect 8988 6862 8990 6914
rect 9042 6862 9044 6914
rect 8988 6850 9044 6862
rect 9212 6692 9268 9436
rect 9324 8372 9380 12236
rect 9996 12178 10052 12190
rect 9996 12126 9998 12178
rect 10050 12126 10052 12178
rect 9548 12066 9604 12078
rect 9548 12014 9550 12066
rect 9602 12014 9604 12066
rect 9548 11394 9604 12014
rect 9548 11342 9550 11394
rect 9602 11342 9604 11394
rect 9548 11330 9604 11342
rect 9996 11284 10052 12126
rect 10220 12180 10276 15484
rect 10332 15428 10388 15438
rect 10332 15334 10388 15372
rect 11452 15148 11508 21980
rect 11564 21026 11620 22876
rect 12460 22372 12516 22990
rect 13468 22372 13524 22382
rect 12460 22306 12516 22316
rect 13356 22370 13524 22372
rect 13356 22318 13470 22370
rect 13522 22318 13524 22370
rect 13356 22316 13524 22318
rect 12796 22260 12852 22270
rect 11564 20974 11566 21026
rect 11618 20974 11620 21026
rect 11564 20962 11620 20974
rect 12684 21588 12740 21598
rect 11676 20690 11732 20702
rect 11676 20638 11678 20690
rect 11730 20638 11732 20690
rect 11564 20578 11620 20590
rect 11564 20526 11566 20578
rect 11618 20526 11620 20578
rect 11564 20020 11620 20526
rect 11564 19954 11620 19964
rect 11676 20132 11732 20638
rect 11676 19012 11732 20076
rect 12684 20130 12740 21532
rect 12684 20078 12686 20130
rect 12738 20078 12740 20130
rect 12684 20066 12740 20078
rect 12236 20018 12292 20030
rect 12236 19966 12238 20018
rect 12290 19966 12292 20018
rect 11676 18956 11956 19012
rect 11788 18004 11844 18014
rect 11676 17892 11732 17902
rect 11676 17108 11732 17836
rect 11676 17014 11732 17052
rect 11788 16212 11844 17948
rect 11788 16146 11844 16156
rect 11340 15092 11508 15148
rect 11564 15314 11620 15326
rect 11564 15262 11566 15314
rect 11618 15262 11620 15314
rect 10668 13524 10724 13534
rect 10668 13074 10724 13468
rect 10668 13022 10670 13074
rect 10722 13022 10724 13074
rect 10668 13010 10724 13022
rect 11116 12852 11172 12862
rect 11116 12758 11172 12796
rect 10444 12180 10500 12190
rect 10220 12178 10500 12180
rect 10220 12126 10446 12178
rect 10498 12126 10500 12178
rect 10220 12124 10500 12126
rect 10444 12114 10500 12124
rect 9996 11218 10052 11228
rect 9660 11172 9716 11182
rect 9548 11170 9716 11172
rect 9548 11118 9662 11170
rect 9714 11118 9716 11170
rect 9548 11116 9716 11118
rect 9548 9826 9604 11116
rect 9660 11106 9716 11116
rect 9548 9774 9550 9826
rect 9602 9774 9604 9826
rect 9548 9762 9604 9774
rect 9996 9714 10052 9726
rect 9996 9662 9998 9714
rect 10050 9662 10052 9714
rect 9996 9604 10052 9662
rect 9996 9538 10052 9548
rect 9660 9268 9716 9278
rect 9660 9174 9716 9212
rect 9436 9044 9492 9054
rect 9436 8950 9492 8988
rect 9884 9042 9940 9054
rect 10108 9044 10164 9054
rect 9884 8990 9886 9042
rect 9938 8990 9940 9042
rect 9324 8306 9380 8316
rect 9884 8148 9940 8990
rect 9884 8082 9940 8092
rect 9996 9042 10164 9044
rect 9996 8990 10110 9042
rect 10162 8990 10164 9042
rect 9996 8988 10164 8990
rect 9660 7700 9716 7710
rect 9660 7606 9716 7644
rect 9884 7700 9940 7710
rect 9996 7700 10052 8988
rect 10108 8978 10164 8988
rect 11340 8596 11396 15092
rect 11564 14642 11620 15262
rect 11564 14590 11566 14642
rect 11618 14590 11620 14642
rect 11564 14578 11620 14590
rect 11788 15204 11844 15214
rect 11452 14306 11508 14318
rect 11452 14254 11454 14306
rect 11506 14254 11508 14306
rect 11452 13524 11508 14254
rect 11676 14308 11732 14318
rect 11676 14214 11732 14252
rect 11452 13458 11508 13468
rect 11452 11620 11508 11630
rect 11788 11620 11844 15148
rect 11900 14980 11956 18956
rect 12236 16772 12292 19966
rect 12796 20018 12852 22204
rect 13356 22260 13412 22316
rect 13468 22306 13524 22316
rect 13692 22372 13748 22382
rect 13804 22372 13860 23996
rect 13916 23716 13972 23726
rect 13916 23622 13972 23660
rect 14028 23714 14084 23726
rect 14028 23662 14030 23714
rect 14082 23662 14084 23714
rect 14028 23268 14084 23662
rect 14028 23202 14084 23212
rect 14140 23714 14196 23726
rect 14140 23662 14142 23714
rect 14194 23662 14196 23714
rect 14028 22596 14084 22606
rect 14028 22502 14084 22540
rect 13692 22370 13860 22372
rect 13692 22318 13694 22370
rect 13746 22318 13860 22370
rect 13692 22316 13860 22318
rect 13692 22306 13748 22316
rect 13356 22194 13412 22204
rect 13468 21588 13524 21598
rect 13468 21494 13524 21532
rect 13804 21586 13860 22316
rect 13916 22146 13972 22158
rect 13916 22094 13918 22146
rect 13970 22094 13972 22146
rect 13916 21812 13972 22094
rect 14140 22148 14196 23662
rect 14140 22082 14196 22092
rect 14252 22370 14308 26908
rect 14588 23044 14644 23054
rect 14476 23042 14644 23044
rect 14476 22990 14590 23042
rect 14642 22990 14644 23042
rect 14476 22988 14644 22990
rect 14476 22482 14532 22988
rect 14588 22978 14644 22988
rect 14700 22932 14756 28588
rect 14812 28578 14868 28588
rect 15372 28532 15428 28542
rect 15372 28082 15428 28476
rect 15372 28030 15374 28082
rect 15426 28030 15428 28082
rect 15036 27634 15092 27646
rect 15036 27582 15038 27634
rect 15090 27582 15092 27634
rect 15036 27074 15092 27582
rect 15372 27634 15428 28030
rect 15372 27582 15374 27634
rect 15426 27582 15428 27634
rect 15372 27570 15428 27582
rect 15036 27022 15038 27074
rect 15090 27022 15092 27074
rect 14812 26964 14868 27002
rect 14812 26898 14868 26908
rect 14812 22932 14868 22942
rect 14700 22876 14812 22932
rect 14476 22430 14478 22482
rect 14530 22430 14532 22482
rect 14476 22418 14532 22430
rect 14252 22318 14254 22370
rect 14306 22318 14308 22370
rect 14252 22036 14308 22318
rect 14588 22260 14644 22270
rect 14588 22166 14644 22204
rect 14700 22148 14756 22158
rect 14252 21980 14532 22036
rect 14364 21812 14420 21822
rect 13916 21756 14364 21812
rect 14364 21698 14420 21756
rect 14364 21646 14366 21698
rect 14418 21646 14420 21698
rect 14364 21634 14420 21646
rect 14476 21700 14532 21980
rect 14700 21810 14756 22092
rect 14700 21758 14702 21810
rect 14754 21758 14756 21810
rect 14700 21746 14756 21758
rect 14476 21634 14532 21644
rect 13804 21534 13806 21586
rect 13858 21534 13860 21586
rect 13804 21522 13860 21534
rect 14588 21588 14644 21598
rect 14588 21494 14644 21532
rect 13916 21474 13972 21486
rect 13916 21422 13918 21474
rect 13970 21422 13972 21474
rect 12796 19966 12798 20018
rect 12850 19966 12852 20018
rect 12796 19954 12852 19966
rect 12908 20804 12964 20814
rect 12460 19908 12516 19918
rect 12460 19814 12516 19852
rect 12908 19122 12964 20748
rect 13804 20132 13860 20142
rect 13356 20020 13412 20030
rect 13356 19926 13412 19964
rect 13692 19908 13748 19918
rect 13692 19458 13748 19852
rect 13692 19406 13694 19458
rect 13746 19406 13748 19458
rect 13692 19394 13748 19406
rect 13804 19906 13860 20076
rect 13804 19854 13806 19906
rect 13858 19854 13860 19906
rect 13580 19348 13636 19358
rect 13468 19292 13580 19348
rect 13468 19234 13524 19292
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 13468 19170 13524 19182
rect 12908 19070 12910 19122
rect 12962 19070 12964 19122
rect 12908 19058 12964 19070
rect 12796 19010 12852 19022
rect 12796 18958 12798 19010
rect 12850 18958 12852 19010
rect 12796 18452 12852 18958
rect 13580 18452 13636 19292
rect 13692 18452 13748 18462
rect 13580 18450 13748 18452
rect 13580 18398 13694 18450
rect 13746 18398 13748 18450
rect 13580 18396 13748 18398
rect 12796 18386 12852 18396
rect 13692 18386 13748 18396
rect 12236 16706 12292 16716
rect 12572 16660 12628 16670
rect 12572 16212 12628 16604
rect 12012 16210 12628 16212
rect 12012 16158 12574 16210
rect 12626 16158 12628 16210
rect 12012 16156 12628 16158
rect 12012 15426 12068 16156
rect 12572 16146 12628 16156
rect 12012 15374 12014 15426
rect 12066 15374 12068 15426
rect 12012 15362 12068 15374
rect 12684 15876 12740 15886
rect 12684 15202 12740 15820
rect 12684 15150 12686 15202
rect 12738 15150 12740 15202
rect 12684 15148 12740 15150
rect 11900 14914 11956 14924
rect 12572 15092 12740 15148
rect 12124 14532 12180 14542
rect 12460 14532 12516 14542
rect 12124 14530 12516 14532
rect 12124 14478 12126 14530
rect 12178 14478 12462 14530
rect 12514 14478 12516 14530
rect 12124 14476 12516 14478
rect 12124 14466 12180 14476
rect 12460 14466 12516 14476
rect 12572 14530 12628 15092
rect 12572 14478 12574 14530
rect 12626 14478 12628 14530
rect 12572 14466 12628 14478
rect 13580 14868 13636 14878
rect 13580 14418 13636 14812
rect 13580 14366 13582 14418
rect 13634 14366 13636 14418
rect 12348 14306 12404 14318
rect 12796 14308 12852 14318
rect 12348 14254 12350 14306
rect 12402 14254 12404 14306
rect 12348 13972 12404 14254
rect 12348 13906 12404 13916
rect 12572 14306 12852 14308
rect 12572 14254 12798 14306
rect 12850 14254 12852 14306
rect 12572 14252 12852 14254
rect 12012 13748 12068 13758
rect 12012 13654 12068 13692
rect 12572 12852 12628 14252
rect 12796 14242 12852 14252
rect 13468 14308 13524 14318
rect 13468 14214 13524 14252
rect 13580 12852 13636 14366
rect 12572 12850 12964 12852
rect 12572 12798 12574 12850
rect 12626 12798 12964 12850
rect 12572 12796 12964 12798
rect 12572 12786 12628 12796
rect 12460 12740 12516 12750
rect 12348 12738 12516 12740
rect 12348 12686 12462 12738
rect 12514 12686 12516 12738
rect 12348 12684 12516 12686
rect 11452 11394 11508 11564
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 11452 11330 11508 11342
rect 11676 11564 11844 11620
rect 12236 11954 12292 11966
rect 12236 11902 12238 11954
rect 12290 11902 12292 11954
rect 12236 11620 12292 11902
rect 11564 11284 11620 11294
rect 11564 11190 11620 11228
rect 11676 11172 11732 11564
rect 12236 11554 12292 11564
rect 11788 11396 11844 11406
rect 12012 11396 12068 11406
rect 12348 11396 12404 12684
rect 12460 12674 12516 12684
rect 12460 12290 12516 12302
rect 12460 12238 12462 12290
rect 12514 12238 12516 12290
rect 12460 11508 12516 12238
rect 12460 11442 12516 11452
rect 12572 12066 12628 12078
rect 12572 12014 12574 12066
rect 12626 12014 12628 12066
rect 11788 11394 12068 11396
rect 11788 11342 11790 11394
rect 11842 11342 12014 11394
rect 12066 11342 12068 11394
rect 11788 11340 12068 11342
rect 11788 11330 11844 11340
rect 12012 11330 12068 11340
rect 12236 11340 12404 11396
rect 12572 11394 12628 12014
rect 12572 11342 12574 11394
rect 12626 11342 12628 11394
rect 11676 11116 11844 11172
rect 11788 8932 11844 11116
rect 12236 9154 12292 11340
rect 12572 11330 12628 11342
rect 12908 11284 12964 12796
rect 13580 12786 13636 12796
rect 13804 12180 13860 19854
rect 13916 18338 13972 21422
rect 14028 21476 14084 21486
rect 14028 19236 14084 21420
rect 14812 21364 14868 22876
rect 14476 21308 14868 21364
rect 14924 21586 14980 21598
rect 14924 21534 14926 21586
rect 14978 21534 14980 21586
rect 14140 20244 14196 20254
rect 14476 20244 14532 21308
rect 14924 21252 14980 21534
rect 14924 21186 14980 21196
rect 15036 20690 15092 27022
rect 15372 27412 15428 27422
rect 15260 24162 15316 24174
rect 15260 24110 15262 24162
rect 15314 24110 15316 24162
rect 15260 24050 15316 24110
rect 15260 23998 15262 24050
rect 15314 23998 15316 24050
rect 15148 23940 15204 23950
rect 15260 23940 15316 23998
rect 15204 23884 15316 23940
rect 15148 23874 15204 23884
rect 15260 23154 15316 23884
rect 15260 23102 15262 23154
rect 15314 23102 15316 23154
rect 15260 23090 15316 23102
rect 15260 22484 15316 22494
rect 15148 22428 15260 22484
rect 15148 22370 15204 22428
rect 15148 22318 15150 22370
rect 15202 22318 15204 22370
rect 15148 22306 15204 22318
rect 15148 21586 15204 21598
rect 15148 21534 15150 21586
rect 15202 21534 15204 21586
rect 15148 21140 15204 21534
rect 15148 21074 15204 21084
rect 15036 20638 15038 20690
rect 15090 20638 15092 20690
rect 15036 20626 15092 20638
rect 14140 20242 14532 20244
rect 14140 20190 14142 20242
rect 14194 20190 14532 20242
rect 14140 20188 14532 20190
rect 14700 20578 14756 20590
rect 14700 20526 14702 20578
rect 14754 20526 14756 20578
rect 14140 20178 14196 20188
rect 14476 20020 14532 20030
rect 14700 20020 14756 20526
rect 15260 20356 15316 22428
rect 15036 20300 15316 20356
rect 14924 20132 14980 20142
rect 15036 20132 15092 20300
rect 14980 20076 15092 20132
rect 15148 20132 15204 20142
rect 14924 20066 14980 20076
rect 15148 20038 15204 20076
rect 15372 20132 15428 27356
rect 15484 26180 15540 32396
rect 15932 32386 15988 32396
rect 16044 30994 16100 32620
rect 16380 31778 16436 32620
rect 16380 31726 16382 31778
rect 16434 31726 16436 31778
rect 16380 31714 16436 31726
rect 16044 30942 16046 30994
rect 16098 30942 16100 30994
rect 16044 30930 16100 30942
rect 16156 31668 16212 31678
rect 16156 30996 16212 31612
rect 16268 31556 16324 31566
rect 16268 31462 16324 31500
rect 16604 31554 16660 31566
rect 16604 31502 16606 31554
rect 16658 31502 16660 31554
rect 16604 31108 16660 31502
rect 16268 30996 16324 31006
rect 16156 30994 16324 30996
rect 16156 30942 16270 30994
rect 16322 30942 16324 30994
rect 16156 30940 16324 30942
rect 16268 30930 16324 30940
rect 16492 30996 16548 31006
rect 16604 30996 16660 31052
rect 16492 30994 16660 30996
rect 16492 30942 16494 30994
rect 16546 30942 16660 30994
rect 16492 30940 16660 30942
rect 16492 30930 16548 30940
rect 16716 29986 16772 33068
rect 17164 33012 17220 33516
rect 17388 33460 17444 33470
rect 17388 33366 17444 33404
rect 17276 33346 17332 33358
rect 17276 33294 17278 33346
rect 17330 33294 17332 33346
rect 17276 33236 17332 33294
rect 17500 33346 17556 33854
rect 17500 33294 17502 33346
rect 17554 33294 17556 33346
rect 17500 33282 17556 33294
rect 17276 33170 17332 33180
rect 17164 32956 17556 33012
rect 17500 32786 17556 32956
rect 17500 32734 17502 32786
rect 17554 32734 17556 32786
rect 17388 32562 17444 32574
rect 17388 32510 17390 32562
rect 17442 32510 17444 32562
rect 17164 31890 17220 31902
rect 17164 31838 17166 31890
rect 17218 31838 17220 31890
rect 16940 31778 16996 31790
rect 16940 31726 16942 31778
rect 16994 31726 16996 31778
rect 16940 31218 16996 31726
rect 16940 31166 16942 31218
rect 16994 31166 16996 31218
rect 16940 31154 16996 31166
rect 17052 30212 17108 30222
rect 17164 30212 17220 31838
rect 17388 31892 17444 32510
rect 17500 32452 17556 32734
rect 17612 32564 17668 34302
rect 18172 34356 18228 37212
rect 18284 37266 18340 37278
rect 18284 37214 18286 37266
rect 18338 37214 18340 37266
rect 18284 37156 18340 37214
rect 18284 34580 18340 37100
rect 18396 36932 18452 37998
rect 18732 38050 18788 38612
rect 18732 37998 18734 38050
rect 18786 37998 18788 38050
rect 18732 37986 18788 37998
rect 19292 38164 19348 38174
rect 18620 37940 18676 37950
rect 18396 36866 18452 36876
rect 18508 37938 18676 37940
rect 18508 37886 18622 37938
rect 18674 37886 18676 37938
rect 18508 37884 18676 37886
rect 18508 35812 18564 37884
rect 18620 37874 18676 37884
rect 18956 37940 19012 37950
rect 18956 37846 19012 37884
rect 19292 37938 19348 38108
rect 19852 38050 19908 38780
rect 20188 38834 20300 38836
rect 20188 38782 20190 38834
rect 20242 38782 20300 38834
rect 20188 38780 20300 38782
rect 20188 38770 20244 38780
rect 20300 38770 20356 38780
rect 20412 38834 20468 38846
rect 20412 38782 20414 38834
rect 20466 38782 20468 38834
rect 19852 37998 19854 38050
rect 19906 37998 19908 38050
rect 19852 37986 19908 37998
rect 20076 38388 20132 38398
rect 19292 37886 19294 37938
rect 19346 37886 19348 37938
rect 19292 37874 19348 37886
rect 20076 37938 20132 38332
rect 20076 37886 20078 37938
rect 20130 37886 20132 37938
rect 20076 37874 20132 37886
rect 20188 37938 20244 37950
rect 20188 37886 20190 37938
rect 20242 37886 20244 37938
rect 18732 37828 18788 37838
rect 18732 37266 18788 37772
rect 19628 37828 19684 37838
rect 19628 37734 19684 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18732 37214 18734 37266
rect 18786 37214 18788 37266
rect 18732 37202 18788 37214
rect 19068 37156 19124 37166
rect 20188 37156 20244 37886
rect 20412 37604 20468 38782
rect 20972 38836 21028 38846
rect 20972 38742 21028 38780
rect 20636 38724 20692 38734
rect 20636 38722 20916 38724
rect 20636 38670 20638 38722
rect 20690 38670 20916 38722
rect 20636 38668 20916 38670
rect 21308 38722 21364 38892
rect 22652 39506 23492 39508
rect 22652 39454 23438 39506
rect 23490 39454 23492 39506
rect 22652 39452 23492 39454
rect 21308 38670 21310 38722
rect 21362 38670 21364 38722
rect 20636 38658 20692 38668
rect 20860 38612 21252 38668
rect 21308 38658 21364 38670
rect 21644 38834 21700 38846
rect 21644 38782 21646 38834
rect 21698 38782 21700 38834
rect 20860 38500 20916 38510
rect 20636 38444 20860 38500
rect 20636 38162 20692 38444
rect 20860 38434 20916 38444
rect 21196 38276 21252 38612
rect 21644 38500 21700 38782
rect 21196 38220 21588 38276
rect 20636 38110 20638 38162
rect 20690 38110 20692 38162
rect 20636 38098 20692 38110
rect 21532 38050 21588 38220
rect 21532 37998 21534 38050
rect 21586 37998 21588 38050
rect 21532 37986 21588 37998
rect 21308 37938 21364 37950
rect 21308 37886 21310 37938
rect 21362 37886 21364 37938
rect 20524 37828 20580 37838
rect 20524 37734 20580 37772
rect 20412 37548 20580 37604
rect 20412 37156 20468 37166
rect 20188 37100 20412 37156
rect 19068 37062 19124 37100
rect 20412 37062 20468 37100
rect 20524 36932 20580 37548
rect 20524 36866 20580 36876
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 18396 35756 18564 35812
rect 19852 35810 19908 35822
rect 19852 35758 19854 35810
rect 19906 35758 19908 35810
rect 18396 35364 18452 35756
rect 18396 34802 18452 35308
rect 18396 34750 18398 34802
rect 18450 34750 18452 34802
rect 18396 34738 18452 34750
rect 19516 35698 19572 35710
rect 19516 35646 19518 35698
rect 19570 35646 19572 35698
rect 18284 34524 18452 34580
rect 18284 34356 18340 34366
rect 18172 34354 18340 34356
rect 18172 34302 18286 34354
rect 18338 34302 18340 34354
rect 18172 34300 18340 34302
rect 17836 34242 17892 34254
rect 17836 34190 17838 34242
rect 17890 34190 17892 34242
rect 17836 33908 17892 34190
rect 17836 33842 17892 33852
rect 17724 32788 17780 32798
rect 18060 32788 18116 32798
rect 17724 32786 18116 32788
rect 17724 32734 17726 32786
rect 17778 32734 18062 32786
rect 18114 32734 18116 32786
rect 17724 32732 18116 32734
rect 17724 32722 17780 32732
rect 18060 32722 18116 32732
rect 17948 32564 18004 32574
rect 17612 32562 18004 32564
rect 17612 32510 17950 32562
rect 18002 32510 18004 32562
rect 17612 32508 18004 32510
rect 17948 32498 18004 32508
rect 17500 32396 17892 32452
rect 17388 31826 17444 31836
rect 17724 32228 17780 32238
rect 17724 31778 17780 32172
rect 17724 31726 17726 31778
rect 17778 31726 17780 31778
rect 17724 31714 17780 31726
rect 17276 31556 17332 31566
rect 17276 31462 17332 31500
rect 17500 31556 17556 31566
rect 17388 31108 17444 31118
rect 17388 31014 17444 31052
rect 17500 30436 17556 31500
rect 17052 30210 17220 30212
rect 17052 30158 17054 30210
rect 17106 30158 17220 30210
rect 17052 30156 17220 30158
rect 17276 30380 17556 30436
rect 17612 30994 17668 31006
rect 17612 30942 17614 30994
rect 17666 30942 17668 30994
rect 17052 30146 17108 30156
rect 16716 29934 16718 29986
rect 16770 29934 16772 29986
rect 16716 29876 16772 29934
rect 17164 29988 17220 29998
rect 17164 29894 17220 29932
rect 16716 27412 16772 29820
rect 17276 29764 17332 30380
rect 17612 30324 17668 30942
rect 17836 30994 17892 32396
rect 17948 31892 18004 31902
rect 17948 31666 18004 31836
rect 17948 31614 17950 31666
rect 18002 31614 18004 31666
rect 17948 31602 18004 31614
rect 18060 31668 18116 31678
rect 18060 31574 18116 31612
rect 17836 30942 17838 30994
rect 17890 30942 17892 30994
rect 17836 30930 17892 30942
rect 18172 30436 18228 34300
rect 18284 34020 18340 34300
rect 18284 33954 18340 33964
rect 18284 33236 18340 33246
rect 18284 32786 18340 33180
rect 18284 32734 18286 32786
rect 18338 32734 18340 32786
rect 18284 32722 18340 32734
rect 18396 32564 18452 34524
rect 18620 34468 18676 34478
rect 18620 34354 18676 34412
rect 19516 34356 19572 35646
rect 19852 35700 19908 35758
rect 19852 35634 19908 35644
rect 21196 35588 21252 35598
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 18620 34302 18622 34354
rect 18674 34302 18676 34354
rect 18620 33346 18676 34302
rect 19068 34300 19572 34356
rect 19740 34356 19796 34366
rect 19740 34354 20132 34356
rect 19740 34302 19742 34354
rect 19794 34302 20132 34354
rect 19740 34300 20132 34302
rect 18844 34132 18900 34142
rect 19068 34132 19124 34300
rect 19740 34290 19796 34300
rect 18844 34130 19124 34132
rect 18844 34078 18846 34130
rect 18898 34078 19124 34130
rect 18844 34076 19124 34078
rect 19180 34130 19236 34142
rect 19180 34078 19182 34130
rect 19234 34078 19236 34130
rect 18620 33294 18622 33346
rect 18674 33294 18676 33346
rect 18620 33282 18676 33294
rect 18732 33348 18788 33358
rect 17500 30210 17556 30222
rect 17500 30158 17502 30210
rect 17554 30158 17556 30210
rect 16716 27346 16772 27356
rect 17164 29708 17332 29764
rect 17388 30098 17444 30110
rect 17388 30046 17390 30098
rect 17442 30046 17444 30098
rect 16044 27074 16100 27086
rect 16044 27022 16046 27074
rect 16098 27022 16100 27074
rect 15596 26852 15652 26862
rect 16044 26852 16100 27022
rect 16716 26962 16772 26974
rect 16716 26910 16718 26962
rect 16770 26910 16772 26962
rect 16716 26908 16772 26910
rect 15596 26850 16100 26852
rect 15596 26798 15598 26850
rect 15650 26798 16100 26850
rect 15596 26796 16100 26798
rect 15596 26786 15652 26796
rect 16044 26180 16100 26796
rect 16380 26852 16772 26908
rect 16268 26180 16324 26190
rect 16044 26178 16324 26180
rect 16044 26126 16270 26178
rect 16322 26126 16324 26178
rect 16044 26124 16324 26126
rect 15484 26114 15540 26124
rect 15596 25620 15652 25630
rect 15596 25526 15652 25564
rect 16268 25506 16324 26124
rect 16268 25454 16270 25506
rect 16322 25454 16324 25506
rect 16268 25284 16324 25454
rect 15708 24162 15764 24174
rect 15708 24110 15710 24162
rect 15762 24110 15764 24162
rect 15708 24052 15764 24110
rect 16268 24052 16324 25228
rect 15708 24050 16324 24052
rect 15708 23998 15710 24050
rect 15762 23998 16324 24050
rect 15708 23996 16324 23998
rect 15708 23986 15764 23996
rect 16044 23938 16100 23996
rect 16044 23886 16046 23938
rect 16098 23886 16100 23938
rect 16044 23874 16100 23886
rect 16268 23380 16324 23390
rect 16380 23380 16436 26852
rect 16828 25284 16884 25294
rect 16828 25190 16884 25228
rect 16268 23378 16436 23380
rect 16268 23326 16270 23378
rect 16322 23326 16436 23378
rect 16268 23324 16436 23326
rect 16828 23826 16884 23838
rect 16828 23774 16830 23826
rect 16882 23774 16884 23826
rect 16828 23380 16884 23774
rect 17052 23380 17108 23390
rect 16828 23324 17052 23380
rect 16268 23314 16324 23324
rect 17052 23314 17108 23324
rect 15596 23268 15652 23278
rect 15596 23154 15652 23212
rect 16156 23266 16212 23278
rect 16156 23214 16158 23266
rect 16210 23214 16212 23266
rect 15596 23102 15598 23154
rect 15650 23102 15652 23154
rect 15596 23090 15652 23102
rect 15932 23154 15988 23166
rect 15932 23102 15934 23154
rect 15986 23102 15988 23154
rect 15932 22820 15988 23102
rect 15932 22754 15988 22764
rect 16156 22484 16212 23214
rect 16828 23042 16884 23054
rect 16828 22990 16830 23042
rect 16882 22990 16884 23042
rect 16828 22932 16884 22990
rect 16828 22866 16884 22876
rect 16156 22418 16212 22428
rect 16940 22484 16996 22494
rect 16940 22390 16996 22428
rect 15708 22372 15764 22382
rect 15708 22278 15764 22316
rect 16044 22372 16100 22382
rect 16044 22278 16100 22316
rect 15484 22258 15540 22270
rect 15484 22206 15486 22258
rect 15538 22206 15540 22258
rect 15484 22036 15540 22206
rect 15596 22260 15652 22270
rect 15596 22166 15652 22204
rect 16604 22146 16660 22158
rect 16604 22094 16606 22146
rect 16658 22094 16660 22146
rect 16604 22036 16660 22094
rect 15484 21980 16660 22036
rect 15596 21476 15652 21486
rect 15652 21420 15764 21476
rect 15596 21382 15652 21420
rect 15484 20132 15540 20142
rect 15372 20130 15540 20132
rect 15372 20078 15486 20130
rect 15538 20078 15540 20130
rect 15372 20076 15540 20078
rect 14812 20020 14868 20030
rect 14476 20018 14868 20020
rect 14476 19966 14478 20018
rect 14530 19966 14814 20018
rect 14866 19966 14868 20018
rect 14476 19964 14868 19966
rect 14252 19236 14308 19246
rect 14028 19234 14308 19236
rect 14028 19182 14254 19234
rect 14306 19182 14308 19234
rect 14028 19180 14308 19182
rect 14252 19170 14308 19180
rect 14028 19012 14084 19022
rect 14028 19010 14308 19012
rect 14028 18958 14030 19010
rect 14082 18958 14308 19010
rect 14028 18956 14308 18958
rect 14028 18946 14084 18956
rect 13916 18286 13918 18338
rect 13970 18286 13972 18338
rect 13916 15986 13972 18286
rect 14140 18226 14196 18238
rect 14140 18174 14142 18226
rect 14194 18174 14196 18226
rect 14140 17668 14196 18174
rect 13916 15934 13918 15986
rect 13970 15934 13972 15986
rect 13916 15922 13972 15934
rect 14028 17612 14196 17668
rect 13692 11508 13748 11518
rect 13692 11414 13748 11452
rect 12684 11228 12964 11284
rect 12236 9102 12238 9154
rect 12290 9102 12292 9154
rect 12236 9090 12292 9102
rect 12348 11172 12404 11182
rect 11788 8838 11844 8876
rect 11340 8530 11396 8540
rect 12124 8484 12180 8494
rect 11676 8260 11732 8270
rect 9884 7698 10052 7700
rect 9884 7646 9886 7698
rect 9938 7646 10052 7698
rect 9884 7644 10052 7646
rect 10556 8148 10612 8158
rect 10556 7698 10612 8092
rect 10556 7646 10558 7698
rect 10610 7646 10612 7698
rect 9884 7634 9940 7644
rect 10556 7634 10612 7646
rect 11228 7924 11284 7934
rect 9772 7588 9828 7598
rect 9772 7494 9828 7532
rect 10668 7588 10724 7598
rect 9996 7474 10052 7486
rect 9996 7422 9998 7474
rect 10050 7422 10052 7474
rect 9772 6916 9828 6926
rect 9996 6916 10052 7422
rect 10220 7476 10276 7486
rect 10220 7382 10276 7420
rect 9772 6914 10052 6916
rect 9772 6862 9774 6914
rect 9826 6862 10052 6914
rect 9772 6860 10052 6862
rect 9772 6850 9828 6860
rect 10556 6804 10612 6814
rect 10668 6804 10724 7532
rect 10556 6802 10668 6804
rect 10556 6750 10558 6802
rect 10610 6750 10668 6802
rect 10556 6748 10668 6750
rect 9324 6692 9380 6702
rect 9100 6690 9380 6692
rect 9100 6638 9326 6690
rect 9378 6638 9380 6690
rect 9100 6636 9380 6638
rect 8428 6526 8430 6578
rect 8482 6526 8484 6578
rect 8428 6514 8484 6526
rect 8764 6580 8820 6590
rect 8092 6468 8148 6478
rect 7868 6466 8148 6468
rect 7868 6414 8094 6466
rect 8146 6414 8148 6466
rect 7868 6412 8148 6414
rect 7644 5954 7700 5964
rect 7308 5730 7364 5740
rect 7084 5684 7140 5694
rect 7084 5590 7140 5628
rect 8092 5572 8148 6412
rect 8092 5506 8148 5516
rect 8652 5348 8708 5358
rect 8764 5348 8820 6524
rect 8876 6468 8932 6478
rect 8876 6374 8932 6412
rect 8876 5348 8932 5358
rect 8764 5346 8932 5348
rect 8764 5294 8878 5346
rect 8930 5294 8932 5346
rect 8764 5292 8932 5294
rect 7756 5236 7812 5246
rect 7756 5142 7812 5180
rect 8540 5124 8596 5134
rect 8540 5030 8596 5068
rect 6076 4114 6244 4116
rect 6076 4062 6078 4114
rect 6130 4062 6244 4114
rect 6076 4060 6244 4062
rect 7196 4226 7252 4238
rect 7196 4174 7198 4226
rect 7250 4174 7252 4226
rect 6076 4050 6132 4060
rect 7196 800 7252 4174
rect 7756 3668 7812 3678
rect 7756 3574 7812 3612
rect 8540 3668 8596 3678
rect 8540 800 8596 3612
rect 8652 3554 8708 5292
rect 8876 5282 8932 5292
rect 8988 5236 9044 5246
rect 8988 5142 9044 5180
rect 8988 4340 9044 4350
rect 9100 4340 9156 6636
rect 9324 6626 9380 6636
rect 10332 6690 10388 6702
rect 10332 6638 10334 6690
rect 10386 6638 10388 6690
rect 9548 6468 9604 6478
rect 9212 5236 9268 5246
rect 9212 5122 9268 5180
rect 9212 5070 9214 5122
rect 9266 5070 9268 5122
rect 9212 5058 9268 5070
rect 9548 5124 9604 6412
rect 9996 6466 10052 6478
rect 9996 6414 9998 6466
rect 10050 6414 10052 6466
rect 9660 6020 9716 6030
rect 9996 6020 10052 6414
rect 9716 5964 10052 6020
rect 9660 5906 9716 5964
rect 9660 5854 9662 5906
rect 9714 5854 9716 5906
rect 9660 5842 9716 5854
rect 10332 5908 10388 6638
rect 10556 6130 10612 6748
rect 10668 6710 10724 6748
rect 11004 6916 11060 6926
rect 10556 6078 10558 6130
rect 10610 6078 10612 6130
rect 10556 6066 10612 6078
rect 10892 6466 10948 6478
rect 10892 6414 10894 6466
rect 10946 6414 10948 6466
rect 10892 6132 10948 6414
rect 10892 6066 10948 6076
rect 10332 5814 10388 5852
rect 11004 5906 11060 6860
rect 11228 6690 11284 7868
rect 11676 6916 11732 8204
rect 11228 6638 11230 6690
rect 11282 6638 11284 6690
rect 11228 6626 11284 6638
rect 11452 6804 11508 6814
rect 11452 6130 11508 6748
rect 11676 6690 11732 6860
rect 11676 6638 11678 6690
rect 11730 6638 11732 6690
rect 11676 6626 11732 6638
rect 11452 6078 11454 6130
rect 11506 6078 11508 6130
rect 11452 6066 11508 6078
rect 12012 6132 12068 6142
rect 11788 6020 11844 6030
rect 11788 5926 11844 5964
rect 11004 5854 11006 5906
rect 11058 5854 11060 5906
rect 11004 5842 11060 5854
rect 9884 5794 9940 5806
rect 9884 5742 9886 5794
rect 9938 5742 9940 5794
rect 9884 5348 9940 5742
rect 10444 5794 10500 5806
rect 10444 5742 10446 5794
rect 10498 5742 10500 5794
rect 9996 5684 10052 5694
rect 10444 5684 10500 5742
rect 9996 5682 10500 5684
rect 9996 5630 9998 5682
rect 10050 5630 10500 5682
rect 9996 5628 10500 5630
rect 10556 5796 10612 5806
rect 9996 5618 10052 5628
rect 9884 5292 10388 5348
rect 9548 5030 9604 5068
rect 9660 5236 9716 5246
rect 8988 4338 9156 4340
rect 8988 4286 8990 4338
rect 9042 4286 9156 4338
rect 8988 4284 9156 4286
rect 8988 4274 9044 4284
rect 9548 3668 9604 3678
rect 9660 3668 9716 5180
rect 10332 5234 10388 5292
rect 10332 5182 10334 5234
rect 10386 5182 10388 5234
rect 10332 5170 10388 5182
rect 10556 4564 10612 5740
rect 10556 4498 10612 4508
rect 12012 4338 12068 6076
rect 12012 4286 12014 4338
rect 12066 4286 12068 4338
rect 12012 4274 12068 4286
rect 9548 3666 9716 3668
rect 9548 3614 9550 3666
rect 9602 3614 9716 3666
rect 9548 3612 9716 3614
rect 10108 4114 10164 4126
rect 10108 4062 10110 4114
rect 10162 4062 10164 4114
rect 9548 3602 9604 3612
rect 8652 3502 8654 3554
rect 8706 3502 8708 3554
rect 8652 3490 8708 3502
rect 10108 3388 10164 4062
rect 9884 3332 10164 3388
rect 11228 3666 11284 3678
rect 11228 3614 11230 3666
rect 11282 3614 11284 3666
rect 9884 800 9940 3332
rect 11228 800 11284 3614
rect 12124 3668 12180 8428
rect 12348 8372 12404 11116
rect 12460 11172 12516 11182
rect 12684 11172 12740 11228
rect 12460 11170 12740 11172
rect 12460 11118 12462 11170
rect 12514 11118 12740 11170
rect 12460 11116 12740 11118
rect 12460 11106 12516 11116
rect 13020 10610 13076 10622
rect 13020 10558 13022 10610
rect 13074 10558 13076 10610
rect 13020 10164 13076 10558
rect 13244 10164 13300 10174
rect 13020 10108 13244 10164
rect 13244 10098 13300 10108
rect 13804 9940 13860 12124
rect 13692 9884 13860 9940
rect 13580 9826 13636 9838
rect 13580 9774 13582 9826
rect 13634 9774 13636 9826
rect 13244 9604 13300 9614
rect 13244 9042 13300 9548
rect 13244 8990 13246 9042
rect 13298 8990 13300 9042
rect 13244 8978 13300 8990
rect 13356 9602 13412 9614
rect 13356 9550 13358 9602
rect 13410 9550 13412 9602
rect 12460 8596 12516 8606
rect 12516 8540 12628 8596
rect 12460 8530 12516 8540
rect 12460 8372 12516 8382
rect 12348 8370 12516 8372
rect 12348 8318 12462 8370
rect 12514 8318 12516 8370
rect 12348 8316 12516 8318
rect 12460 8306 12516 8316
rect 12236 8258 12292 8270
rect 12236 8206 12238 8258
rect 12290 8206 12292 8258
rect 12236 8148 12292 8206
rect 12236 8082 12292 8092
rect 12572 6132 12628 8540
rect 12684 8372 12740 8382
rect 12684 8258 12740 8316
rect 12684 8206 12686 8258
rect 12738 8206 12740 8258
rect 12684 8194 12740 8206
rect 12908 8146 12964 8158
rect 12908 8094 12910 8146
rect 12962 8094 12964 8146
rect 12908 6804 12964 8094
rect 13356 7252 13412 9550
rect 13580 8482 13636 9774
rect 13580 8430 13582 8482
rect 13634 8430 13636 8482
rect 13580 8418 13636 8430
rect 13692 8260 13748 9884
rect 13692 8194 13748 8204
rect 13804 9716 13860 9726
rect 13580 8036 13636 8046
rect 13580 7474 13636 7980
rect 13580 7422 13582 7474
rect 13634 7422 13636 7474
rect 13580 7410 13636 7422
rect 13692 7476 13748 7486
rect 13356 7196 13524 7252
rect 13468 7140 13524 7196
rect 13468 7084 13636 7140
rect 12908 6738 12964 6748
rect 13468 6692 13524 6702
rect 12684 6468 12740 6478
rect 12684 6374 12740 6412
rect 12684 6132 12740 6142
rect 12572 6130 12740 6132
rect 12572 6078 12686 6130
rect 12738 6078 12740 6130
rect 12572 6076 12740 6078
rect 12460 6020 12516 6030
rect 12460 5234 12516 5964
rect 12460 5182 12462 5234
rect 12514 5182 12516 5234
rect 12460 5170 12516 5182
rect 12684 5012 12740 6076
rect 13132 6132 13188 6142
rect 13132 5906 13188 6076
rect 13468 6130 13524 6636
rect 13468 6078 13470 6130
rect 13522 6078 13524 6130
rect 13468 6066 13524 6078
rect 13132 5854 13134 5906
rect 13186 5854 13188 5906
rect 13132 5842 13188 5854
rect 12908 5796 12964 5806
rect 12908 5702 12964 5740
rect 12796 5348 12852 5358
rect 12796 5254 12852 5292
rect 13580 5122 13636 7084
rect 13692 6916 13748 7420
rect 13804 7474 13860 9660
rect 13916 9714 13972 9726
rect 13916 9662 13918 9714
rect 13970 9662 13972 9714
rect 13916 9154 13972 9662
rect 13916 9102 13918 9154
rect 13970 9102 13972 9154
rect 13916 9090 13972 9102
rect 13916 8260 13972 8270
rect 13916 8166 13972 8204
rect 13804 7422 13806 7474
rect 13858 7422 13860 7474
rect 13804 7410 13860 7422
rect 13692 6802 13748 6860
rect 13692 6750 13694 6802
rect 13746 6750 13748 6802
rect 13692 6738 13748 6750
rect 13916 6132 13972 6142
rect 13916 6038 13972 6076
rect 13580 5070 13582 5122
rect 13634 5070 13636 5122
rect 13580 5058 13636 5070
rect 12908 5012 12964 5022
rect 12684 5010 12964 5012
rect 12684 4958 12910 5010
rect 12962 4958 12964 5010
rect 12684 4956 12964 4958
rect 12908 4946 12964 4956
rect 13804 4898 13860 4910
rect 13804 4846 13806 4898
rect 13858 4846 13860 4898
rect 13804 4340 13860 4846
rect 13804 4274 13860 4284
rect 12124 3554 12180 3612
rect 12124 3502 12126 3554
rect 12178 3502 12180 3554
rect 12124 3490 12180 3502
rect 13020 4114 13076 4126
rect 13020 4062 13022 4114
rect 13074 4062 13076 4114
rect 13020 3388 13076 4062
rect 13132 3668 13188 3678
rect 13188 3612 13300 3668
rect 13132 3602 13188 3612
rect 13244 3554 13300 3612
rect 13244 3502 13246 3554
rect 13298 3502 13300 3554
rect 13244 3490 13300 3502
rect 14028 3554 14084 17612
rect 14140 15986 14196 15998
rect 14140 15934 14142 15986
rect 14194 15934 14196 15986
rect 14140 9826 14196 15934
rect 14140 9774 14142 9826
rect 14194 9774 14196 9826
rect 14140 9762 14196 9774
rect 14252 9826 14308 18956
rect 14476 18676 14532 19964
rect 14812 19954 14868 19964
rect 14812 19460 14868 19470
rect 14588 19348 14644 19358
rect 14588 19254 14644 19292
rect 14812 19122 14868 19404
rect 14812 19070 14814 19122
rect 14866 19070 14868 19122
rect 14812 19058 14868 19070
rect 14588 19012 14644 19022
rect 14588 19010 14756 19012
rect 14588 18958 14590 19010
rect 14642 18958 14756 19010
rect 14588 18956 14756 18958
rect 14588 18946 14644 18956
rect 14588 18676 14644 18686
rect 14476 18674 14644 18676
rect 14476 18622 14590 18674
rect 14642 18622 14644 18674
rect 14476 18620 14644 18622
rect 14588 18610 14644 18620
rect 14700 18564 14756 18956
rect 15148 19010 15204 19022
rect 15148 18958 15150 19010
rect 15202 18958 15204 19010
rect 14700 18508 14868 18564
rect 14700 18338 14756 18350
rect 14700 18286 14702 18338
rect 14754 18286 14756 18338
rect 14700 18004 14756 18286
rect 14812 18228 14868 18508
rect 15148 18340 15204 18958
rect 14812 18162 14868 18172
rect 15036 18284 15204 18340
rect 15036 18004 15092 18284
rect 14700 17948 15092 18004
rect 14364 16212 14420 16222
rect 14364 15986 14420 16156
rect 14364 15934 14366 15986
rect 14418 15934 14420 15986
rect 14364 15922 14420 15934
rect 14588 15988 14644 15998
rect 14588 15894 14644 15932
rect 14476 15874 14532 15886
rect 14476 15822 14478 15874
rect 14530 15822 14532 15874
rect 14476 15540 14532 15822
rect 14924 15876 14980 15886
rect 14924 15782 14980 15820
rect 14476 15484 14868 15540
rect 14812 15426 14868 15484
rect 14812 15374 14814 15426
rect 14866 15374 14868 15426
rect 14812 15362 14868 15374
rect 15036 15148 15092 17948
rect 14252 9774 14254 9826
rect 14306 9774 14308 9826
rect 14140 8932 14196 8942
rect 14140 8146 14196 8876
rect 14140 8094 14142 8146
rect 14194 8094 14196 8146
rect 14140 8082 14196 8094
rect 14140 6690 14196 6702
rect 14140 6638 14142 6690
rect 14194 6638 14196 6690
rect 14140 6580 14196 6638
rect 14140 6514 14196 6524
rect 14140 6356 14196 6366
rect 14140 5234 14196 6300
rect 14252 6018 14308 9774
rect 14364 15092 15092 15148
rect 15260 16100 15316 16110
rect 15260 15874 15316 16044
rect 15260 15822 15262 15874
rect 15314 15822 15316 15874
rect 14364 6692 14420 15092
rect 15260 14868 15316 15822
rect 15260 14802 15316 14812
rect 15148 14530 15204 14542
rect 15148 14478 15150 14530
rect 15202 14478 15204 14530
rect 14588 14308 14644 14318
rect 14588 14214 14644 14252
rect 15148 13972 15204 14478
rect 15148 13906 15204 13916
rect 15036 13636 15092 13646
rect 15036 13542 15092 13580
rect 14700 11508 14756 11518
rect 14700 9826 14756 11452
rect 14700 9774 14702 9826
rect 14754 9774 14756 9826
rect 14700 9762 14756 9774
rect 15036 11172 15092 11182
rect 15036 9714 15092 11116
rect 15036 9662 15038 9714
rect 15090 9662 15092 9714
rect 15036 9650 15092 9662
rect 15372 9492 15428 20076
rect 15484 20066 15540 20076
rect 15484 19796 15540 19806
rect 15484 19012 15540 19740
rect 15484 18918 15540 18956
rect 15708 16212 15764 21420
rect 15932 20132 15988 20142
rect 15932 20018 15988 20076
rect 16380 20132 16436 20142
rect 16380 20038 16436 20076
rect 15932 19966 15934 20018
rect 15986 19966 15988 20018
rect 15932 19954 15988 19966
rect 15932 19460 15988 19470
rect 15932 19346 15988 19404
rect 15932 19294 15934 19346
rect 15986 19294 15988 19346
rect 15932 19282 15988 19294
rect 16604 18116 16660 21980
rect 17164 21028 17220 29708
rect 17388 29650 17444 30046
rect 17500 29876 17556 30158
rect 17500 29810 17556 29820
rect 17388 29598 17390 29650
rect 17442 29598 17444 29650
rect 17388 29586 17444 29598
rect 17612 29538 17668 30268
rect 17836 30380 18228 30436
rect 18284 32508 18452 32564
rect 17724 30212 17780 30222
rect 17724 29988 17780 30156
rect 17724 29922 17780 29932
rect 17612 29486 17614 29538
rect 17666 29486 17668 29538
rect 16828 20972 17220 21028
rect 17276 29316 17332 29326
rect 16716 20130 16772 20142
rect 16716 20078 16718 20130
rect 16770 20078 16772 20130
rect 16716 20020 16772 20078
rect 16716 18900 16772 19964
rect 16716 18834 16772 18844
rect 16604 18050 16660 18060
rect 15820 17668 15876 17678
rect 16156 17668 16212 17678
rect 15820 17666 16212 17668
rect 15820 17614 15822 17666
rect 15874 17614 16158 17666
rect 16210 17614 16212 17666
rect 15820 17612 16212 17614
rect 15820 17602 15876 17612
rect 15708 16118 15764 16156
rect 16044 15540 16100 17612
rect 16156 17602 16212 17612
rect 15596 15538 16100 15540
rect 15596 15486 16046 15538
rect 16098 15486 16100 15538
rect 15596 15484 16100 15486
rect 15596 15314 15652 15484
rect 16044 15474 16100 15484
rect 15596 15262 15598 15314
rect 15650 15262 15652 15314
rect 15596 13636 15652 15262
rect 15596 13570 15652 13580
rect 16156 15204 16212 15214
rect 15820 12404 15876 12414
rect 15820 11506 15876 12348
rect 15820 11454 15822 11506
rect 15874 11454 15876 11506
rect 15820 11442 15876 11454
rect 15372 9426 15428 9436
rect 15932 8372 15988 8382
rect 15260 8260 15316 8270
rect 15260 8166 15316 8204
rect 15932 8258 15988 8316
rect 15932 8206 15934 8258
rect 15986 8206 15988 8258
rect 15932 8194 15988 8206
rect 16044 8370 16100 8382
rect 16044 8318 16046 8370
rect 16098 8318 16100 8370
rect 16044 8260 16100 8318
rect 14700 8148 14756 8158
rect 15148 8148 15204 8158
rect 14476 8092 14700 8148
rect 14476 7586 14532 8092
rect 14700 8054 14756 8092
rect 14812 8146 15204 8148
rect 14812 8094 15150 8146
rect 15202 8094 15204 8146
rect 14812 8092 15204 8094
rect 14476 7534 14478 7586
rect 14530 7534 14532 7586
rect 14476 7522 14532 7534
rect 14812 7364 14868 8092
rect 15148 8082 15204 8092
rect 15372 8148 15428 8158
rect 15372 8054 15428 8092
rect 16044 8036 16100 8204
rect 15820 7980 16100 8036
rect 15820 7700 15876 7980
rect 16156 7924 16212 15148
rect 16828 15148 16884 20972
rect 17052 20132 17108 20142
rect 17052 19234 17108 20076
rect 17052 19182 17054 19234
rect 17106 19182 17108 19234
rect 17052 19170 17108 19182
rect 17276 17892 17332 29260
rect 17612 29092 17668 29486
rect 17724 29540 17780 29550
rect 17724 29446 17780 29484
rect 17612 29026 17668 29036
rect 17836 26908 17892 30380
rect 18284 30324 18340 32508
rect 18620 31668 18676 31678
rect 18620 31554 18676 31612
rect 18620 31502 18622 31554
rect 18674 31502 18676 31554
rect 18620 30996 18676 31502
rect 18732 31108 18788 33292
rect 18844 31332 18900 34076
rect 19180 34020 19236 34078
rect 19180 33954 19236 33964
rect 19628 34132 19684 34142
rect 19628 33460 19684 34076
rect 19628 33366 19684 33404
rect 19852 34130 19908 34142
rect 19852 34078 19854 34130
rect 19906 34078 19908 34130
rect 19068 33348 19124 33358
rect 19068 33254 19124 33292
rect 19852 33236 19908 34078
rect 20076 33346 20132 34300
rect 20972 34020 21028 34030
rect 20972 33926 21028 33964
rect 20300 33460 20356 33470
rect 20076 33294 20078 33346
rect 20130 33294 20132 33346
rect 20076 33282 20132 33294
rect 20188 33348 20244 33358
rect 19852 33170 19908 33180
rect 19516 33124 19572 33134
rect 19516 32564 19572 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32788 19684 32798
rect 19628 32694 19684 32732
rect 19852 32564 19908 32574
rect 19516 32562 19908 32564
rect 19516 32510 19854 32562
rect 19906 32510 19908 32562
rect 19516 32508 19908 32510
rect 19292 32450 19348 32462
rect 19292 32398 19294 32450
rect 19346 32398 19348 32450
rect 19292 32340 19348 32398
rect 19516 32340 19572 32350
rect 19292 32284 19516 32340
rect 19516 32246 19572 32284
rect 19852 32228 19908 32508
rect 20188 32452 20244 33292
rect 20300 33346 20356 33404
rect 20300 33294 20302 33346
rect 20354 33294 20356 33346
rect 20300 33282 20356 33294
rect 20524 33348 20580 33358
rect 20524 33254 20580 33292
rect 20636 33236 20692 33246
rect 20636 33142 20692 33180
rect 20188 32450 20580 32452
rect 20188 32398 20190 32450
rect 20242 32398 20580 32450
rect 20188 32396 20580 32398
rect 20188 32386 20244 32396
rect 19852 32172 20356 32228
rect 20300 31666 20356 32172
rect 20524 31778 20580 32396
rect 20524 31726 20526 31778
rect 20578 31726 20580 31778
rect 20524 31714 20580 31726
rect 20300 31614 20302 31666
rect 20354 31614 20356 31666
rect 20300 31602 20356 31614
rect 18956 31556 19012 31566
rect 19012 31500 19124 31556
rect 18956 31462 19012 31500
rect 18844 31276 19012 31332
rect 18844 31108 18900 31118
rect 18732 31106 18900 31108
rect 18732 31054 18846 31106
rect 18898 31054 18900 31106
rect 18732 31052 18900 31054
rect 18844 31042 18900 31052
rect 18508 30940 18620 30996
rect 17948 30268 18340 30324
rect 18396 30324 18452 30334
rect 17948 28084 18004 30268
rect 18396 30210 18452 30268
rect 18396 30158 18398 30210
rect 18450 30158 18452 30210
rect 18396 30146 18452 30158
rect 18172 30100 18228 30110
rect 18060 30098 18228 30100
rect 18060 30046 18174 30098
rect 18226 30046 18228 30098
rect 18060 30044 18228 30046
rect 18060 29988 18116 30044
rect 18172 30034 18228 30044
rect 18060 29922 18116 29932
rect 18396 29988 18452 29998
rect 18396 29894 18452 29932
rect 18172 29540 18228 29550
rect 18508 29540 18564 30940
rect 18620 30930 18676 30940
rect 18732 30772 18788 30782
rect 18620 30770 18788 30772
rect 18620 30718 18734 30770
rect 18786 30718 18788 30770
rect 18620 30716 18788 30718
rect 18620 30212 18676 30716
rect 18732 30706 18788 30716
rect 18620 30146 18676 30156
rect 18732 30100 18788 30110
rect 18732 30006 18788 30044
rect 18228 29484 18564 29540
rect 18172 29446 18228 29484
rect 17948 28018 18004 28028
rect 18844 27188 18900 27198
rect 18956 27188 19012 31276
rect 19068 31108 19124 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19180 31108 19236 31118
rect 19068 31052 19180 31108
rect 19180 31042 19236 31052
rect 20412 30212 20468 30222
rect 19068 29988 19124 29998
rect 19068 29538 19124 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19068 29486 19070 29538
rect 19122 29486 19124 29538
rect 19068 29474 19124 29486
rect 19180 29540 19236 29550
rect 19180 29446 19236 29484
rect 18844 27186 19012 27188
rect 18844 27134 18846 27186
rect 18898 27134 19012 27186
rect 18844 27132 19012 27134
rect 19404 29426 19460 29438
rect 19404 29374 19406 29426
rect 19458 29374 19460 29426
rect 18844 27122 18900 27132
rect 19404 26908 19460 29374
rect 20188 28644 20244 28654
rect 20188 28550 20244 28588
rect 20412 28530 20468 30156
rect 20636 29428 20692 29438
rect 20636 29334 20692 29372
rect 21196 29316 21252 35532
rect 21308 33908 21364 37886
rect 21644 36932 21700 38444
rect 22428 38722 22484 38734
rect 22428 38670 22430 38722
rect 22482 38670 22484 38722
rect 21868 38164 21924 38174
rect 22316 38164 22372 38174
rect 21868 38162 22372 38164
rect 21868 38110 21870 38162
rect 21922 38110 22318 38162
rect 22370 38110 22372 38162
rect 21868 38108 22372 38110
rect 21868 38098 21924 38108
rect 22316 38098 22372 38108
rect 21868 37940 21924 37950
rect 21868 37846 21924 37884
rect 21756 37828 21812 37838
rect 21756 37156 21812 37772
rect 22428 37828 22484 38670
rect 22652 38274 22708 39452
rect 23436 39442 23492 39452
rect 22876 38948 22932 38958
rect 22876 38854 22932 38892
rect 22652 38222 22654 38274
rect 22706 38222 22708 38274
rect 22652 38210 22708 38222
rect 22428 37762 22484 37772
rect 22652 38050 22708 38062
rect 22652 37998 22654 38050
rect 22706 37998 22708 38050
rect 22652 37380 22708 37998
rect 24108 37940 24164 37950
rect 24164 37884 24276 37940
rect 24108 37874 24164 37884
rect 23100 37828 23156 37838
rect 23100 37734 23156 37772
rect 22652 37314 22708 37324
rect 21756 37090 21812 37100
rect 22204 37154 22260 37166
rect 22204 37102 22206 37154
rect 22258 37102 22260 37154
rect 21420 36876 21700 36932
rect 22204 37044 22260 37102
rect 23548 37156 23604 37166
rect 23548 37154 24164 37156
rect 23548 37102 23550 37154
rect 23602 37102 24164 37154
rect 23548 37100 24164 37102
rect 23548 37090 23604 37100
rect 21420 36594 21476 36876
rect 22204 36708 22260 36988
rect 21420 36542 21422 36594
rect 21474 36542 21476 36594
rect 21420 35700 21476 36542
rect 21868 36652 22260 36708
rect 22428 36932 22484 36942
rect 21420 35634 21476 35644
rect 21644 36484 21700 36494
rect 21868 36484 21924 36652
rect 21644 36482 21924 36484
rect 21644 36430 21646 36482
rect 21698 36430 21924 36482
rect 21644 36428 21924 36430
rect 21980 36484 22036 36494
rect 22316 36484 22372 36494
rect 21980 36482 22372 36484
rect 21980 36430 21982 36482
rect 22034 36430 22318 36482
rect 22370 36430 22372 36482
rect 21980 36428 22372 36430
rect 21644 35588 21700 36428
rect 21980 36418 22036 36428
rect 22316 36418 22372 36428
rect 22428 36258 22484 36876
rect 22428 36206 22430 36258
rect 22482 36206 22484 36258
rect 22428 36194 22484 36206
rect 22764 36484 22820 36494
rect 22764 35810 22820 36428
rect 23436 36484 23492 36494
rect 23884 36484 23940 36494
rect 24108 36484 24164 37100
rect 23492 36482 23940 36484
rect 23492 36430 23886 36482
rect 23938 36430 23940 36482
rect 23492 36428 23940 36430
rect 23436 36390 23492 36428
rect 23884 36418 23940 36428
rect 23996 36482 24164 36484
rect 23996 36430 24110 36482
rect 24162 36430 24164 36482
rect 23996 36428 24164 36430
rect 22764 35758 22766 35810
rect 22818 35758 22820 35810
rect 22764 35746 22820 35758
rect 23324 36370 23380 36382
rect 23324 36318 23326 36370
rect 23378 36318 23380 36370
rect 22204 35700 22260 35710
rect 22204 35606 22260 35644
rect 21868 35588 21924 35598
rect 21644 35532 21868 35588
rect 21868 35494 21924 35532
rect 23212 35588 23268 35598
rect 23212 35494 23268 35532
rect 22876 35028 22932 35038
rect 21308 33842 21364 33852
rect 21644 34020 21700 34030
rect 21308 33348 21364 33358
rect 21532 33348 21588 33358
rect 21364 33346 21588 33348
rect 21364 33294 21534 33346
rect 21586 33294 21588 33346
rect 21364 33292 21588 33294
rect 21308 33282 21364 33292
rect 21532 33282 21588 33292
rect 21308 33122 21364 33134
rect 21308 33070 21310 33122
rect 21362 33070 21364 33122
rect 21308 32788 21364 33070
rect 21420 33124 21476 33134
rect 21644 33124 21700 33964
rect 21756 33908 21812 33918
rect 21756 33348 21812 33852
rect 21756 33292 21924 33348
rect 21756 33124 21812 33134
rect 21420 33030 21476 33068
rect 21532 33122 21812 33124
rect 21532 33070 21758 33122
rect 21810 33070 21812 33122
rect 21532 33068 21812 33070
rect 21308 32722 21364 32732
rect 21196 29250 21252 29260
rect 21308 29314 21364 29326
rect 21308 29262 21310 29314
rect 21362 29262 21364 29314
rect 21308 28756 21364 29262
rect 21308 28690 21364 28700
rect 20748 28644 20804 28654
rect 20748 28550 20804 28588
rect 20412 28478 20414 28530
rect 20466 28478 20468 28530
rect 20412 28466 20468 28478
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 21532 26908 21588 33068
rect 21756 33058 21812 33068
rect 21868 32900 21924 33292
rect 21756 32844 21924 32900
rect 22316 33124 22372 33134
rect 21644 32340 21700 32350
rect 21644 27972 21700 32284
rect 21756 31666 21812 32844
rect 22316 32674 22372 33068
rect 22316 32622 22318 32674
rect 22370 32622 22372 32674
rect 22316 32610 22372 32622
rect 21756 31614 21758 31666
rect 21810 31614 21812 31666
rect 21756 31602 21812 31614
rect 22092 31554 22148 31566
rect 22092 31502 22094 31554
rect 22146 31502 22148 31554
rect 22092 30996 22148 31502
rect 22652 30996 22708 31006
rect 22092 30994 22708 30996
rect 22092 30942 22654 30994
rect 22706 30942 22708 30994
rect 22092 30940 22708 30942
rect 22652 30324 22708 30940
rect 21756 28532 21812 28542
rect 22652 28532 22708 30268
rect 22764 28756 22820 28766
rect 22764 28662 22820 28700
rect 22652 28476 22820 28532
rect 21756 28082 21812 28476
rect 22652 28084 22708 28094
rect 21756 28030 21758 28082
rect 21810 28030 21812 28082
rect 21756 28018 21812 28030
rect 21980 28028 22652 28084
rect 21644 27878 21700 27916
rect 21980 27970 22036 28028
rect 22652 27990 22708 28028
rect 21980 27918 21982 27970
rect 22034 27918 22036 27970
rect 17836 26852 18340 26908
rect 19404 26852 19684 26908
rect 18284 26516 18340 26852
rect 17500 26180 17556 26190
rect 17500 25844 17556 26124
rect 17500 25778 17556 25788
rect 17948 25506 18004 25518
rect 17948 25454 17950 25506
rect 18002 25454 18004 25506
rect 17500 25284 17556 25294
rect 17500 25190 17556 25228
rect 17948 25284 18004 25454
rect 17948 25218 18004 25228
rect 18284 24722 18340 26460
rect 18844 26180 18900 26190
rect 18732 26124 18844 26180
rect 18284 24670 18286 24722
rect 18338 24670 18340 24722
rect 18284 24658 18340 24670
rect 18620 25394 18676 25406
rect 18620 25342 18622 25394
rect 18674 25342 18676 25394
rect 17500 23380 17556 23390
rect 17500 23286 17556 23324
rect 18172 23380 18228 23390
rect 17612 23268 17668 23278
rect 17388 23154 17444 23166
rect 17388 23102 17390 23154
rect 17442 23102 17444 23154
rect 17388 22820 17444 23102
rect 17388 22754 17444 22764
rect 17388 20132 17444 20142
rect 17388 20038 17444 20076
rect 17612 19908 17668 23212
rect 17724 23154 17780 23166
rect 17724 23102 17726 23154
rect 17778 23102 17780 23154
rect 17724 22372 17780 23102
rect 18172 23154 18228 23324
rect 18620 23378 18676 25342
rect 18620 23326 18622 23378
rect 18674 23326 18676 23378
rect 18620 23314 18676 23326
rect 18172 23102 18174 23154
rect 18226 23102 18228 23154
rect 17948 22932 18004 22942
rect 17948 22838 18004 22876
rect 18172 22484 18228 23102
rect 18508 23156 18564 23166
rect 18172 22418 18228 22428
rect 18396 22932 18452 22942
rect 17948 22372 18004 22382
rect 17724 22370 18004 22372
rect 17724 22318 17950 22370
rect 18002 22318 18004 22370
rect 17724 22316 18004 22318
rect 17948 22306 18004 22316
rect 18284 22372 18340 22382
rect 18284 22278 18340 22316
rect 17836 22148 17892 22158
rect 18172 22148 18228 22158
rect 17836 22146 18228 22148
rect 17836 22094 17838 22146
rect 17890 22094 18174 22146
rect 18226 22094 18228 22146
rect 17836 22092 18228 22094
rect 17836 22082 17892 22092
rect 17836 19908 17892 19918
rect 17612 19906 17892 19908
rect 17612 19854 17838 19906
rect 17890 19854 17892 19906
rect 17612 19852 17892 19854
rect 17276 17826 17332 17836
rect 17388 19010 17444 19022
rect 17388 18958 17390 19010
rect 17442 18958 17444 19010
rect 17388 18564 17444 18958
rect 17388 17668 17444 18508
rect 17388 17612 17780 17668
rect 16940 17554 16996 17566
rect 16940 17502 16942 17554
rect 16994 17502 16996 17554
rect 16940 17108 16996 17502
rect 17612 17108 17668 17118
rect 16940 17106 17668 17108
rect 16940 17054 17614 17106
rect 17666 17054 17668 17106
rect 16940 17052 17668 17054
rect 17612 17042 17668 17052
rect 17388 16884 17444 16894
rect 17388 15148 17444 16828
rect 17724 16324 17780 17612
rect 17836 17108 17892 19852
rect 17836 16884 17892 17052
rect 17836 16790 17892 16828
rect 17948 18452 18004 18462
rect 17948 16882 18004 18396
rect 17948 16830 17950 16882
rect 18002 16830 18004 16882
rect 17948 16818 18004 16830
rect 18060 16436 18116 22092
rect 18172 22082 18228 22092
rect 18396 19908 18452 22876
rect 18396 19842 18452 19852
rect 18508 21586 18564 23100
rect 18732 22036 18788 26124
rect 18844 26114 18900 26124
rect 18844 24724 18900 24734
rect 18844 24630 18900 24668
rect 19292 24724 19348 24734
rect 19292 24630 19348 24668
rect 18956 24050 19012 24062
rect 18956 23998 18958 24050
rect 19010 23998 19012 24050
rect 18732 21970 18788 21980
rect 18844 23154 18900 23166
rect 18844 23102 18846 23154
rect 18898 23102 18900 23154
rect 18844 21924 18900 23102
rect 18956 22372 19012 23998
rect 19516 23714 19572 23726
rect 19516 23662 19518 23714
rect 19570 23662 19572 23714
rect 19516 23604 19572 23662
rect 19516 23538 19572 23548
rect 19516 23380 19572 23390
rect 19068 23378 19572 23380
rect 19068 23326 19518 23378
rect 19570 23326 19572 23378
rect 19068 23324 19572 23326
rect 19628 23380 19684 26852
rect 20636 26852 21588 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20076 26290 20132 26302
rect 20076 26238 20078 26290
rect 20130 26238 20132 26290
rect 20076 25284 20132 26238
rect 20076 25228 20244 25284
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 23940 20244 25228
rect 20300 23940 20356 23950
rect 20188 23884 20300 23940
rect 20300 23874 20356 23884
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23324 19908 23380
rect 19068 23266 19124 23324
rect 19516 23314 19572 23324
rect 19068 23214 19070 23266
rect 19122 23214 19124 23266
rect 19068 23202 19124 23214
rect 19180 23156 19236 23166
rect 19404 23156 19460 23166
rect 19236 23154 19460 23156
rect 19236 23102 19406 23154
rect 19458 23102 19460 23154
rect 19236 23100 19460 23102
rect 19180 23090 19236 23100
rect 19404 23090 19460 23100
rect 19628 23154 19684 23166
rect 19628 23102 19630 23154
rect 19682 23102 19684 23154
rect 18956 22306 19012 22316
rect 19516 23044 19572 23054
rect 19068 22260 19124 22270
rect 18956 22148 19012 22158
rect 18956 22054 19012 22092
rect 19068 21924 19124 22204
rect 18844 21868 19124 21924
rect 18508 21534 18510 21586
rect 18562 21534 18564 21586
rect 18284 18676 18340 18686
rect 18284 18582 18340 18620
rect 18396 18450 18452 18462
rect 18396 18398 18398 18450
rect 18450 18398 18452 18450
rect 18284 18226 18340 18238
rect 18284 18174 18286 18226
rect 18338 18174 18340 18226
rect 18284 16996 18340 18174
rect 18396 17780 18452 18398
rect 18508 18452 18564 21534
rect 18732 21810 18788 21822
rect 18732 21758 18734 21810
rect 18786 21758 18788 21810
rect 18732 21476 18788 21758
rect 18844 21586 18900 21868
rect 18844 21534 18846 21586
rect 18898 21534 18900 21586
rect 18844 21522 18900 21534
rect 19068 21588 19124 21598
rect 18732 21410 18788 21420
rect 18844 21026 18900 21038
rect 18844 20974 18846 21026
rect 18898 20974 18900 21026
rect 18844 20914 18900 20974
rect 18844 20862 18846 20914
rect 18898 20862 18900 20914
rect 18844 20580 18900 20862
rect 18844 20514 18900 20524
rect 19068 20244 19124 21532
rect 19404 21586 19460 21598
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 19404 21026 19460 21534
rect 19404 20974 19406 21026
rect 19458 20974 19460 21026
rect 19404 20962 19460 20974
rect 19068 20178 19124 20188
rect 19292 20578 19348 20590
rect 19292 20526 19294 20578
rect 19346 20526 19348 20578
rect 18956 20018 19012 20030
rect 18956 19966 18958 20018
rect 19010 19966 19012 20018
rect 18844 19348 18900 19358
rect 18844 18676 18900 19292
rect 18956 19012 19012 19966
rect 19292 20020 19348 20526
rect 19292 19954 19348 19964
rect 19404 20020 19460 20030
rect 19516 20020 19572 22988
rect 19628 22260 19684 23102
rect 19628 22194 19684 22204
rect 19852 22258 19908 23324
rect 19964 23154 20020 23166
rect 19964 23102 19966 23154
rect 20018 23102 20020 23154
rect 19964 23044 20020 23102
rect 19964 22978 20020 22988
rect 20412 23044 20468 23054
rect 20412 22950 20468 22988
rect 19852 22206 19854 22258
rect 19906 22206 19908 22258
rect 19852 22194 19908 22206
rect 20076 22370 20132 22382
rect 20076 22318 20078 22370
rect 20130 22318 20132 22370
rect 20076 22148 20132 22318
rect 20412 22260 20468 22270
rect 20412 22166 20468 22204
rect 20076 22092 20244 22148
rect 19628 22036 19684 22046
rect 19628 21026 19684 21980
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 22092
rect 20076 21756 20244 21812
rect 20076 21588 20132 21756
rect 20076 21522 20132 21532
rect 19628 20974 19630 21026
rect 19682 20974 19684 21026
rect 19628 20962 19684 20974
rect 19964 21476 20020 21486
rect 19964 21026 20020 21420
rect 19964 20974 19966 21026
rect 20018 20974 20020 21026
rect 19964 20962 20020 20974
rect 19740 20804 19796 20814
rect 19404 20018 19572 20020
rect 19404 19966 19406 20018
rect 19458 19966 19572 20018
rect 19404 19964 19572 19966
rect 19628 20802 19796 20804
rect 19628 20750 19742 20802
rect 19794 20750 19796 20802
rect 19628 20748 19796 20750
rect 19628 20020 19684 20748
rect 19740 20738 19796 20748
rect 20076 20802 20132 20814
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20580 20132 20750
rect 20076 20524 20244 20580
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19404 19954 19460 19964
rect 19628 19954 19684 19964
rect 19740 20244 19796 20254
rect 19740 20018 19796 20188
rect 20188 20188 20244 20524
rect 20188 20132 20580 20188
rect 20524 20038 20580 20076
rect 19740 19966 19742 20018
rect 19794 19966 19796 20018
rect 19740 19954 19796 19966
rect 19964 20018 20020 20030
rect 19964 19966 19966 20018
rect 20018 19966 20020 20018
rect 19964 19796 20020 19966
rect 19516 19740 20020 19796
rect 20076 20018 20132 20030
rect 20076 19966 20078 20018
rect 20130 19966 20132 20018
rect 19516 19236 19572 19740
rect 18956 18946 19012 18956
rect 19292 19010 19348 19022
rect 19292 18958 19294 19010
rect 19346 18958 19348 19010
rect 18844 18452 18900 18620
rect 18508 18386 18564 18396
rect 18620 18450 18900 18452
rect 18620 18398 18846 18450
rect 18898 18398 18900 18450
rect 18620 18396 18900 18398
rect 18620 18228 18676 18396
rect 18844 18386 18900 18396
rect 19292 18452 19348 18958
rect 19516 18676 19572 19180
rect 20076 19236 20132 19966
rect 20636 19684 20692 26852
rect 20748 26180 20804 26190
rect 20748 26086 20804 26124
rect 20748 25620 20804 25630
rect 20748 25526 20804 25564
rect 21756 23940 21812 23950
rect 21756 23846 21812 23884
rect 21644 23828 21700 23838
rect 21532 23772 21644 23828
rect 20748 22146 20804 22158
rect 20748 22094 20750 22146
rect 20802 22094 20804 22146
rect 20748 20580 20804 22094
rect 21308 20580 21364 20590
rect 20748 20578 21364 20580
rect 20748 20526 21310 20578
rect 21362 20526 21364 20578
rect 20748 20524 21364 20526
rect 20636 19346 20692 19628
rect 20636 19294 20638 19346
rect 20690 19294 20692 19346
rect 20636 19282 20692 19294
rect 21196 19908 21252 19918
rect 20076 19180 20356 19236
rect 19628 19124 19684 19134
rect 19628 19030 19684 19068
rect 20076 19124 20132 19180
rect 20076 19058 20132 19068
rect 20188 19012 20244 19022
rect 20188 18918 20244 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 18676 19796 18686
rect 19516 18674 19796 18676
rect 19516 18622 19742 18674
rect 19794 18622 19796 18674
rect 19516 18620 19796 18622
rect 19740 18610 19796 18620
rect 19852 18676 19908 18686
rect 19852 18562 19908 18620
rect 19852 18510 19854 18562
rect 19906 18510 19908 18562
rect 19852 18498 19908 18510
rect 19292 18386 19348 18396
rect 19628 18340 19684 18350
rect 19068 18228 19124 18238
rect 18396 17714 18452 17724
rect 18508 18172 18676 18228
rect 18956 18172 19068 18228
rect 18396 16996 18452 17006
rect 18284 16994 18452 16996
rect 18284 16942 18398 16994
rect 18450 16942 18452 16994
rect 18284 16940 18452 16942
rect 18396 16930 18452 16940
rect 18172 16884 18228 16894
rect 18172 16790 18228 16828
rect 18508 16548 18564 18172
rect 18396 16492 18564 16548
rect 18732 17780 18788 17790
rect 18172 16436 18228 16446
rect 18060 16380 18172 16436
rect 18172 16370 18228 16380
rect 17724 16268 18116 16324
rect 17836 15988 17892 15998
rect 17724 15876 17780 15886
rect 17724 15538 17780 15820
rect 17724 15486 17726 15538
rect 17778 15486 17780 15538
rect 17724 15474 17780 15486
rect 17836 15538 17892 15932
rect 17836 15486 17838 15538
rect 17890 15486 17892 15538
rect 17836 15474 17892 15486
rect 16828 15092 17220 15148
rect 16268 14308 16324 14318
rect 16268 13970 16324 14252
rect 16268 13918 16270 13970
rect 16322 13918 16324 13970
rect 16268 13748 16324 13918
rect 16268 13682 16324 13692
rect 16604 11394 16660 11406
rect 16604 11342 16606 11394
rect 16658 11342 16660 11394
rect 16604 11172 16660 11342
rect 17052 11172 17108 11182
rect 16604 11170 17108 11172
rect 16604 11118 17054 11170
rect 17106 11118 17108 11170
rect 16604 11116 17108 11118
rect 16604 10724 16660 11116
rect 17052 11106 17108 11116
rect 16156 7858 16212 7868
rect 16380 10722 16660 10724
rect 16380 10670 16606 10722
rect 16658 10670 16660 10722
rect 16380 10668 16660 10670
rect 14364 6626 14420 6636
rect 14588 7308 14868 7364
rect 15260 7698 15876 7700
rect 15260 7646 15822 7698
rect 15874 7646 15876 7698
rect 15260 7644 15876 7646
rect 14588 6690 14644 7308
rect 15260 6692 15316 7644
rect 15820 7634 15876 7644
rect 15820 6916 15876 6926
rect 15484 6804 15540 6814
rect 14588 6638 14590 6690
rect 14642 6638 14644 6690
rect 14588 6626 14644 6638
rect 15148 6636 15316 6692
rect 15372 6692 15428 6730
rect 15148 6578 15204 6636
rect 15372 6626 15428 6636
rect 15148 6526 15150 6578
rect 15202 6526 15204 6578
rect 15148 6514 15204 6526
rect 14252 5966 14254 6018
rect 14306 5966 14308 6018
rect 14252 5954 14308 5966
rect 15036 6466 15092 6478
rect 15036 6414 15038 6466
rect 15090 6414 15092 6466
rect 15036 6020 15092 6414
rect 15260 6468 15316 6478
rect 15484 6468 15540 6748
rect 15596 6692 15652 6702
rect 15596 6598 15652 6636
rect 15260 6466 15540 6468
rect 15260 6414 15262 6466
rect 15314 6414 15540 6466
rect 15260 6412 15540 6414
rect 15260 6402 15316 6412
rect 15372 6244 15428 6254
rect 15036 5954 15092 5964
rect 15148 6018 15204 6030
rect 15148 5966 15150 6018
rect 15202 5966 15204 6018
rect 14140 5182 14142 5234
rect 14194 5182 14196 5234
rect 14140 5170 14196 5182
rect 14364 5682 14420 5694
rect 14364 5630 14366 5682
rect 14418 5630 14420 5682
rect 14028 3502 14030 3554
rect 14082 3502 14084 3554
rect 14028 3490 14084 3502
rect 14364 3556 14420 5630
rect 15148 5684 15204 5966
rect 15372 5906 15428 6188
rect 15372 5854 15374 5906
rect 15426 5854 15428 5906
rect 15372 5842 15428 5854
rect 15820 6018 15876 6860
rect 16380 6690 16436 10668
rect 16604 10658 16660 10668
rect 16940 10052 16996 10062
rect 16940 9602 16996 9996
rect 16940 9550 16942 9602
rect 16994 9550 16996 9602
rect 16940 9044 16996 9550
rect 16940 8978 16996 8988
rect 16492 8372 16548 8382
rect 16492 8278 16548 8316
rect 17052 7700 17108 7710
rect 16380 6638 16382 6690
rect 16434 6638 16436 6690
rect 15820 5966 15822 6018
rect 15874 5966 15876 6018
rect 15820 5684 15876 5966
rect 16156 6580 16212 6590
rect 16156 5906 16212 6524
rect 16380 6468 16436 6638
rect 16716 6916 16772 6926
rect 16716 6690 16772 6860
rect 16716 6638 16718 6690
rect 16770 6638 16772 6690
rect 16716 6626 16772 6638
rect 17052 6690 17108 7644
rect 17052 6638 17054 6690
rect 17106 6638 17108 6690
rect 17052 6626 17108 6638
rect 16940 6580 16996 6590
rect 16940 6486 16996 6524
rect 16380 6402 16436 6412
rect 17164 6356 17220 15092
rect 17276 15092 17444 15148
rect 17612 15314 17668 15326
rect 17612 15262 17614 15314
rect 17666 15262 17668 15314
rect 17612 15148 17668 15262
rect 17948 15314 18004 15326
rect 17948 15262 17950 15314
rect 18002 15262 18004 15314
rect 17612 15092 17892 15148
rect 17276 8260 17332 15092
rect 17612 14980 17668 14990
rect 17612 14308 17668 14924
rect 17612 14306 17780 14308
rect 17612 14254 17614 14306
rect 17666 14254 17780 14306
rect 17612 14252 17780 14254
rect 17612 14242 17668 14252
rect 17612 13972 17668 13982
rect 17724 13972 17780 14252
rect 17836 14196 17892 15092
rect 17948 14756 18004 15262
rect 17948 14690 18004 14700
rect 17836 14130 17892 14140
rect 17948 14306 18004 14318
rect 17948 14254 17950 14306
rect 18002 14254 18004 14306
rect 17948 13972 18004 14254
rect 17724 13916 18004 13972
rect 17612 13878 17668 13916
rect 17948 13748 18004 13916
rect 17948 13654 18004 13692
rect 17948 12964 18004 12974
rect 17948 12290 18004 12908
rect 17948 12238 17950 12290
rect 18002 12238 18004 12290
rect 17948 12226 18004 12238
rect 17612 12178 17668 12190
rect 17612 12126 17614 12178
rect 17666 12126 17668 12178
rect 17612 11396 17668 12126
rect 18060 12180 18116 16268
rect 18172 16212 18228 16222
rect 18228 16156 18340 16212
rect 18172 16118 18228 16156
rect 18172 15314 18228 15326
rect 18172 15262 18174 15314
rect 18226 15262 18228 15314
rect 18172 13970 18228 15262
rect 18284 14756 18340 16156
rect 18396 15764 18452 16492
rect 18396 15698 18452 15708
rect 18508 16324 18564 16334
rect 18508 15428 18564 16268
rect 18620 16212 18676 16222
rect 18620 15986 18676 16156
rect 18732 16212 18788 17724
rect 18956 17220 19012 18172
rect 19068 18162 19124 18172
rect 19068 17778 19124 17790
rect 19068 17726 19070 17778
rect 19122 17726 19124 17778
rect 19068 17668 19124 17726
rect 19628 17668 19684 18284
rect 19740 18228 19796 18238
rect 19740 18134 19796 18172
rect 20188 17892 20244 17902
rect 20300 17892 20356 19180
rect 20188 17890 20356 17892
rect 20188 17838 20190 17890
rect 20242 17838 20356 17890
rect 20188 17836 20356 17838
rect 20188 17826 20244 17836
rect 19068 17612 19572 17668
rect 19516 17554 19572 17612
rect 19628 17574 19684 17612
rect 19740 17780 19796 17790
rect 19740 17666 19796 17724
rect 19740 17614 19742 17666
rect 19794 17614 19796 17666
rect 19740 17602 19796 17614
rect 19516 17502 19518 17554
rect 19570 17502 19572 17554
rect 18956 17164 19460 17220
rect 18844 17108 18900 17118
rect 18844 17014 18900 17052
rect 19292 16884 19348 16894
rect 19292 16770 19348 16828
rect 19292 16718 19294 16770
rect 19346 16718 19348 16770
rect 19292 16324 19348 16718
rect 18732 16210 19236 16212
rect 18732 16158 18734 16210
rect 18786 16158 19236 16210
rect 18732 16156 19236 16158
rect 18732 16146 18788 16156
rect 18620 15934 18622 15986
rect 18674 15934 18676 15986
rect 18620 15922 18676 15934
rect 18844 15986 18900 15998
rect 18844 15934 18846 15986
rect 18898 15934 18900 15986
rect 18508 15362 18564 15372
rect 18620 15652 18676 15662
rect 18396 15204 18452 15242
rect 18620 15148 18676 15596
rect 18844 15540 18900 15934
rect 18396 15138 18452 15148
rect 18508 15092 18676 15148
rect 18732 15484 18900 15540
rect 18956 15988 19012 15998
rect 18284 14700 18452 14756
rect 18172 13918 18174 13970
rect 18226 13918 18228 13970
rect 18172 13906 18228 13918
rect 18284 14306 18340 14318
rect 18284 14254 18286 14306
rect 18338 14254 18340 14306
rect 18284 14196 18340 14254
rect 18284 13300 18340 14140
rect 18396 13972 18452 14700
rect 18508 13972 18564 15092
rect 18620 14756 18676 14766
rect 18732 14756 18788 15484
rect 18844 15092 18900 15102
rect 18844 14998 18900 15036
rect 18732 14700 18900 14756
rect 18620 14662 18676 14700
rect 18732 14530 18788 14542
rect 18732 14478 18734 14530
rect 18786 14478 18788 14530
rect 18732 14196 18788 14478
rect 18732 14130 18788 14140
rect 18508 13916 18676 13972
rect 18396 13878 18452 13916
rect 18508 13746 18564 13758
rect 18508 13694 18510 13746
rect 18562 13694 18564 13746
rect 18508 13412 18564 13694
rect 18620 13636 18676 13916
rect 18620 13570 18676 13580
rect 18844 13412 18900 14700
rect 18956 14530 19012 15932
rect 19068 15874 19124 15886
rect 19068 15822 19070 15874
rect 19122 15822 19124 15874
rect 19068 15540 19124 15822
rect 19068 15314 19124 15484
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 19068 15250 19124 15262
rect 18956 14478 18958 14530
rect 19010 14478 19012 14530
rect 18956 14308 19012 14478
rect 19180 14530 19236 16156
rect 19292 15986 19348 16268
rect 19404 16212 19460 17164
rect 19516 16996 19572 17502
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19516 16940 19684 16996
rect 19404 16156 19572 16212
rect 19292 15934 19294 15986
rect 19346 15934 19348 15986
rect 19292 15922 19348 15934
rect 19404 15986 19460 15998
rect 19404 15934 19406 15986
rect 19458 15934 19460 15986
rect 19404 15876 19460 15934
rect 19404 15810 19460 15820
rect 19516 15652 19572 16156
rect 19292 15596 19572 15652
rect 19292 15314 19348 15596
rect 19292 15262 19294 15314
rect 19346 15262 19348 15314
rect 19292 15250 19348 15262
rect 19404 15316 19460 15326
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 19180 14466 19236 14478
rect 18956 14252 19348 14308
rect 19180 13858 19236 13870
rect 19180 13806 19182 13858
rect 19234 13806 19236 13858
rect 19180 13748 19236 13806
rect 19292 13860 19348 14252
rect 19404 14196 19460 15260
rect 19516 15204 19572 15242
rect 19516 15138 19572 15148
rect 19516 14532 19572 14542
rect 19628 14532 19684 16940
rect 20748 16548 20804 16558
rect 19852 16324 19908 16334
rect 19852 16210 19908 16268
rect 19852 16158 19854 16210
rect 19906 16158 19908 16210
rect 19852 16146 19908 16158
rect 20188 16212 20244 16222
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19740 15538 19796 15550
rect 19740 15486 19742 15538
rect 19794 15486 19796 15538
rect 19740 15428 19796 15486
rect 20076 15540 20132 15550
rect 20076 15446 20132 15484
rect 19740 15362 19796 15372
rect 19852 15426 19908 15438
rect 19852 15374 19854 15426
rect 19906 15374 19908 15426
rect 19852 14642 19908 15374
rect 20188 14756 20244 16156
rect 20748 15538 20804 16492
rect 20748 15486 20750 15538
rect 20802 15486 20804 15538
rect 20300 15316 20356 15326
rect 20300 15222 20356 15260
rect 20748 15204 20804 15486
rect 20748 15138 20804 15148
rect 21196 15148 21252 19852
rect 21308 19236 21364 20524
rect 21532 20130 21588 23772
rect 21644 23762 21700 23772
rect 21980 23156 22036 27918
rect 22204 27860 22260 27870
rect 22204 27858 22372 27860
rect 22204 27806 22206 27858
rect 22258 27806 22372 27858
rect 22204 27804 22372 27806
rect 22204 27794 22260 27804
rect 22316 27634 22372 27804
rect 22316 27582 22318 27634
rect 22370 27582 22372 27634
rect 22316 27570 22372 27582
rect 22764 25508 22820 28476
rect 22876 28196 22932 34972
rect 23324 34692 23380 36318
rect 23996 35028 24052 36428
rect 24108 36418 24164 36428
rect 24220 36260 24276 37884
rect 24108 35924 24164 35934
rect 24220 35924 24276 36204
rect 24108 35922 24276 35924
rect 24108 35870 24110 35922
rect 24162 35870 24276 35922
rect 24108 35868 24276 35870
rect 24444 37380 24500 37390
rect 24108 35858 24164 35868
rect 24332 35812 24388 35822
rect 24332 35698 24388 35756
rect 24332 35646 24334 35698
rect 24386 35646 24388 35698
rect 24332 35634 24388 35646
rect 23996 34962 24052 34972
rect 23324 34690 23492 34692
rect 23324 34638 23326 34690
rect 23378 34638 23492 34690
rect 23324 34636 23492 34638
rect 23324 34626 23380 34636
rect 23100 32788 23156 32798
rect 23100 32562 23156 32732
rect 23100 32510 23102 32562
rect 23154 32510 23156 32562
rect 23100 32498 23156 32510
rect 23212 31108 23268 31118
rect 23212 31014 23268 31052
rect 23436 29314 23492 34636
rect 24444 33124 24500 37324
rect 24668 37380 24724 39564
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 24668 37314 24724 37324
rect 28252 37380 28308 37390
rect 28252 37266 28308 37324
rect 28812 37380 28868 37390
rect 28812 37286 28868 37324
rect 28252 37214 28254 37266
rect 28306 37214 28308 37266
rect 24556 37156 24612 37166
rect 24556 37062 24612 37100
rect 25340 37154 25396 37166
rect 25340 37102 25342 37154
rect 25394 37102 25396 37154
rect 24668 37044 24724 37054
rect 25340 37044 25396 37102
rect 27580 37156 27636 37166
rect 27580 37062 27636 37100
rect 24668 37042 25172 37044
rect 24668 36990 24670 37042
rect 24722 36990 25172 37042
rect 24668 36988 25172 36990
rect 24668 36978 24724 36988
rect 25116 36596 25172 36988
rect 25228 36596 25284 36606
rect 25116 36594 25284 36596
rect 25116 36542 25230 36594
rect 25282 36542 25284 36594
rect 25116 36540 25284 36542
rect 25228 36530 25284 36540
rect 25340 36482 25396 36988
rect 26236 37044 26292 37054
rect 26236 36594 26292 36988
rect 26236 36542 26238 36594
rect 26290 36542 26292 36594
rect 26236 36530 26292 36542
rect 25340 36430 25342 36482
rect 25394 36430 25396 36482
rect 25340 36418 25396 36430
rect 24780 36372 24836 36382
rect 24780 36278 24836 36316
rect 25564 36372 25620 36382
rect 25564 36278 25620 36316
rect 25788 36370 25844 36382
rect 25788 36318 25790 36370
rect 25842 36318 25844 36370
rect 24892 36260 24948 36270
rect 25228 36260 25284 36270
rect 24948 36258 25284 36260
rect 24948 36206 25230 36258
rect 25282 36206 25284 36258
rect 24948 36204 25284 36206
rect 24892 36194 24948 36204
rect 25228 36194 25284 36204
rect 25004 35812 25060 35822
rect 25788 35812 25844 36318
rect 25060 35756 25172 35812
rect 25004 35746 25060 35756
rect 24444 33058 24500 33068
rect 23548 32788 23604 32798
rect 23548 32694 23604 32732
rect 25116 32788 25172 35756
rect 25788 35746 25844 35756
rect 26684 35812 26740 35822
rect 25340 35028 25396 35038
rect 25340 34130 25396 34972
rect 25340 34078 25342 34130
rect 25394 34078 25396 34130
rect 25228 32788 25284 32798
rect 25116 32786 25284 32788
rect 25116 32734 25230 32786
rect 25282 32734 25284 32786
rect 25116 32732 25284 32734
rect 23660 32676 23716 32686
rect 23660 30994 23716 32620
rect 25116 32676 25172 32732
rect 25228 32722 25284 32732
rect 25340 32788 25396 34078
rect 26012 34020 26068 34030
rect 25564 34018 26068 34020
rect 25564 33966 26014 34018
rect 26066 33966 26068 34018
rect 25564 33964 26068 33966
rect 25564 33458 25620 33964
rect 26012 33954 26068 33964
rect 25564 33406 25566 33458
rect 25618 33406 25620 33458
rect 25564 33394 25620 33406
rect 25676 33460 25732 33470
rect 26124 33460 26180 33470
rect 25676 33458 26180 33460
rect 25676 33406 25678 33458
rect 25730 33406 26126 33458
rect 26178 33406 26180 33458
rect 25676 33404 26180 33406
rect 25676 33394 25732 33404
rect 26124 33394 26180 33404
rect 26684 33346 26740 35756
rect 28252 35700 28308 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 33068 36260 33124 36270
rect 33068 36166 33124 36204
rect 33404 36258 33460 36270
rect 33404 36206 33406 36258
rect 33458 36206 33460 36258
rect 33404 35812 33460 36206
rect 33404 35746 33460 35756
rect 33740 36260 33796 36270
rect 28252 35698 28420 35700
rect 28252 35646 28254 35698
rect 28306 35646 28420 35698
rect 28252 35644 28420 35646
rect 28252 35634 28308 35644
rect 28364 35028 28420 35644
rect 28364 34934 28420 34972
rect 28924 35586 28980 35598
rect 28924 35534 28926 35586
rect 28978 35534 28980 35586
rect 28924 34354 28980 35534
rect 31052 35586 31108 35598
rect 31052 35534 31054 35586
rect 31106 35534 31108 35586
rect 29372 34692 29428 34702
rect 28924 34302 28926 34354
rect 28978 34302 28980 34354
rect 28924 34290 28980 34302
rect 29148 34690 29428 34692
rect 29148 34638 29374 34690
rect 29426 34638 29428 34690
rect 29148 34636 29428 34638
rect 29148 34356 29204 34636
rect 29372 34626 29428 34636
rect 29148 34262 29204 34300
rect 29596 34242 29652 34254
rect 30828 34244 30884 34254
rect 29596 34190 29598 34242
rect 29650 34190 29652 34242
rect 29260 34130 29316 34142
rect 29260 34078 29262 34130
rect 29314 34078 29316 34130
rect 28140 34020 28196 34030
rect 26684 33294 26686 33346
rect 26738 33294 26740 33346
rect 26684 33282 26740 33294
rect 28028 34018 28196 34020
rect 28028 33966 28142 34018
rect 28194 33966 28196 34018
rect 28028 33964 28196 33966
rect 25340 32722 25396 32732
rect 25452 33124 25508 33134
rect 26124 33124 26180 33134
rect 25116 32610 25172 32620
rect 25452 32452 25508 33068
rect 26012 33122 26180 33124
rect 26012 33070 26126 33122
rect 26178 33070 26180 33122
rect 26012 33068 26180 33070
rect 25564 32676 25620 32686
rect 26012 32676 26068 33068
rect 26124 33058 26180 33068
rect 26236 33124 26292 33134
rect 26460 33124 26516 33134
rect 26236 33122 26404 33124
rect 26236 33070 26238 33122
rect 26290 33070 26404 33122
rect 26236 33068 26404 33070
rect 26236 33058 26292 33068
rect 25564 32674 26068 32676
rect 25564 32622 25566 32674
rect 25618 32622 26068 32674
rect 25564 32620 26068 32622
rect 25564 32610 25620 32620
rect 23660 30942 23662 30994
rect 23714 30942 23716 30994
rect 23660 30322 23716 30942
rect 25116 32396 25508 32452
rect 24108 30884 24164 30894
rect 24108 30790 24164 30828
rect 23660 30270 23662 30322
rect 23714 30270 23716 30322
rect 23660 30258 23716 30270
rect 23996 30324 24052 30334
rect 23996 30230 24052 30268
rect 24220 30212 24276 30222
rect 25004 30212 25060 30222
rect 25116 30212 25172 32396
rect 26012 31444 26068 32620
rect 26012 31378 26068 31388
rect 26124 32676 26180 32686
rect 26348 32676 26404 33068
rect 26460 33122 26628 33124
rect 26460 33070 26462 33122
rect 26514 33070 26628 33122
rect 26460 33068 26628 33070
rect 26460 33058 26516 33068
rect 26572 32788 26628 33068
rect 26572 32732 26852 32788
rect 26124 32674 26404 32676
rect 26124 32622 26126 32674
rect 26178 32622 26404 32674
rect 26124 32620 26404 32622
rect 26796 32674 26852 32732
rect 26796 32622 26798 32674
rect 26850 32622 26852 32674
rect 26124 31220 26180 32620
rect 26796 32610 26852 32622
rect 26460 32564 26516 32574
rect 26124 31164 26292 31220
rect 24220 30210 24948 30212
rect 24220 30158 24222 30210
rect 24274 30158 24948 30210
rect 24220 30156 24948 30158
rect 24220 30146 24276 30156
rect 24892 29986 24948 30156
rect 25060 30156 25172 30212
rect 25788 30660 25844 30670
rect 25004 30146 25060 30156
rect 24892 29934 24894 29986
rect 24946 29934 24948 29986
rect 23436 29262 23438 29314
rect 23490 29262 23492 29314
rect 23436 29250 23492 29262
rect 23548 29428 23604 29438
rect 22876 28130 22932 28140
rect 23100 27972 23156 27982
rect 23100 27878 23156 27916
rect 22876 27636 22932 27646
rect 22876 27634 23044 27636
rect 22876 27582 22878 27634
rect 22930 27582 23044 27634
rect 22876 27580 23044 27582
rect 22876 27570 22932 27580
rect 22988 27524 23044 27580
rect 22988 27468 23156 27524
rect 22876 26180 22932 26190
rect 22876 26086 22932 26124
rect 23100 26068 23156 27468
rect 23548 26908 23604 29372
rect 23996 29428 24052 29438
rect 23996 29334 24052 29372
rect 23772 28532 23828 28542
rect 23772 28438 23828 28476
rect 22988 26012 23156 26068
rect 23324 26852 23604 26908
rect 23324 26178 23380 26852
rect 23324 26126 23326 26178
rect 23378 26126 23380 26178
rect 22092 25452 22932 25508
rect 22092 24946 22148 25452
rect 22764 25284 22820 25294
rect 22092 24894 22094 24946
rect 22146 24894 22148 24946
rect 22092 24882 22148 24894
rect 22652 25282 22820 25284
rect 22652 25230 22766 25282
rect 22818 25230 22820 25282
rect 22652 25228 22820 25230
rect 22428 24724 22484 24734
rect 22652 24724 22708 25228
rect 22764 25218 22820 25228
rect 22484 24668 22708 24724
rect 22428 24630 22484 24668
rect 22428 23828 22484 23838
rect 22428 23734 22484 23772
rect 21644 20690 21700 20702
rect 21644 20638 21646 20690
rect 21698 20638 21700 20690
rect 21644 20356 21700 20638
rect 21644 20290 21700 20300
rect 21532 20078 21534 20130
rect 21586 20078 21588 20130
rect 21532 20066 21588 20078
rect 21644 19908 21700 19918
rect 21644 19814 21700 19852
rect 21868 19908 21924 19918
rect 21868 19814 21924 19852
rect 21308 19142 21364 19180
rect 21868 19460 21924 19470
rect 21532 19122 21588 19134
rect 21532 19070 21534 19122
rect 21586 19070 21588 19122
rect 21532 18676 21588 19070
rect 21644 19124 21700 19134
rect 21644 19030 21700 19068
rect 21868 18788 21924 19404
rect 21868 18722 21924 18732
rect 21532 18610 21588 18620
rect 21868 18004 21924 18014
rect 21980 18004 22036 23100
rect 22540 23266 22596 23278
rect 22540 23214 22542 23266
rect 22594 23214 22596 23266
rect 22092 23044 22148 23054
rect 22540 23044 22596 23214
rect 22148 22988 22596 23044
rect 22092 22950 22148 22988
rect 22540 22932 22596 22988
rect 22540 22866 22596 22876
rect 22652 20356 22708 24668
rect 22876 24722 22932 25452
rect 22876 24670 22878 24722
rect 22930 24670 22932 24722
rect 22876 24658 22932 24670
rect 22876 23380 22932 23390
rect 22988 23380 23044 26012
rect 22876 23378 23044 23380
rect 22876 23326 22878 23378
rect 22930 23326 23044 23378
rect 22876 23324 23044 23326
rect 23100 25844 23156 25854
rect 22876 23314 22932 23324
rect 22764 23156 22820 23166
rect 22764 23062 22820 23100
rect 22988 23156 23044 23166
rect 22988 23062 23044 23100
rect 22988 21476 23044 21486
rect 23100 21476 23156 25788
rect 23324 25284 23380 26126
rect 23324 25228 23604 25284
rect 23324 24610 23380 24622
rect 23324 24558 23326 24610
rect 23378 24558 23380 24610
rect 23324 23156 23380 24558
rect 23548 23940 23604 25228
rect 24668 24724 24724 24734
rect 24556 24164 24612 24174
rect 24556 24050 24612 24108
rect 24556 23998 24558 24050
rect 24610 23998 24612 24050
rect 24556 23986 24612 23998
rect 23548 23874 23604 23884
rect 23660 23380 23716 23390
rect 23436 23156 23492 23166
rect 23324 23100 23436 23156
rect 23436 23042 23492 23100
rect 23436 22990 23438 23042
rect 23490 22990 23492 23042
rect 23436 22036 23492 22990
rect 23436 21970 23492 21980
rect 22988 21474 23156 21476
rect 22988 21422 22990 21474
rect 23042 21422 23156 21474
rect 22988 21420 23156 21422
rect 22876 20804 22932 20814
rect 22876 20710 22932 20748
rect 22652 20300 22932 20356
rect 22652 20132 22708 20142
rect 22092 20018 22148 20030
rect 22092 19966 22094 20018
rect 22146 19966 22148 20018
rect 22092 19460 22148 19966
rect 22652 19906 22708 20076
rect 22652 19854 22654 19906
rect 22706 19854 22708 19906
rect 22652 19842 22708 19854
rect 22092 19458 22820 19460
rect 22092 19406 22094 19458
rect 22146 19406 22820 19458
rect 22092 19404 22820 19406
rect 22092 19394 22148 19404
rect 22764 19122 22820 19404
rect 22764 19070 22766 19122
rect 22818 19070 22820 19122
rect 22764 19058 22820 19070
rect 22876 18116 22932 20300
rect 21924 17948 22036 18004
rect 22652 18060 22932 18116
rect 21868 17938 21924 17948
rect 22540 17668 22596 17678
rect 22540 17574 22596 17612
rect 22540 16772 22596 16782
rect 22092 16436 22148 16446
rect 21196 15092 21364 15148
rect 19852 14590 19854 14642
rect 19906 14590 19908 14642
rect 19852 14578 19908 14590
rect 19964 14700 20356 14756
rect 19572 14476 19684 14532
rect 19964 14530 20020 14700
rect 19964 14478 19966 14530
rect 20018 14478 20020 14530
rect 19516 14438 19572 14476
rect 19964 14466 20020 14478
rect 20188 14530 20244 14542
rect 20188 14478 20190 14530
rect 20242 14478 20244 14530
rect 19740 14308 19796 14318
rect 19404 14130 19460 14140
rect 19516 14306 19796 14308
rect 19516 14254 19742 14306
rect 19794 14254 19796 14306
rect 19516 14252 19796 14254
rect 19404 13860 19460 13870
rect 19292 13858 19460 13860
rect 19292 13806 19406 13858
rect 19458 13806 19460 13858
rect 19292 13804 19460 13806
rect 19404 13794 19460 13804
rect 19180 13682 19236 13692
rect 19068 13522 19124 13534
rect 19068 13470 19070 13522
rect 19122 13470 19124 13522
rect 18508 13356 19012 13412
rect 18284 13244 18564 13300
rect 18284 12404 18340 12442
rect 18284 12338 18340 12348
rect 18284 12180 18340 12190
rect 18060 12178 18452 12180
rect 18060 12126 18286 12178
rect 18338 12126 18452 12178
rect 18060 12124 18452 12126
rect 18284 12114 18340 12124
rect 17836 12066 17892 12078
rect 17836 12014 17838 12066
rect 17890 12014 17892 12066
rect 17612 11330 17668 11340
rect 17724 11844 17780 11854
rect 17724 11394 17780 11788
rect 17836 11620 17892 12014
rect 17836 11554 17892 11564
rect 17724 11342 17726 11394
rect 17778 11342 17780 11394
rect 17724 11330 17780 11342
rect 18060 11396 18116 11406
rect 18396 11396 18452 12124
rect 18508 11844 18564 13244
rect 18732 13076 18788 13086
rect 18620 13074 18788 13076
rect 18620 13022 18734 13074
rect 18786 13022 18788 13074
rect 18620 13020 18788 13022
rect 18620 12178 18676 13020
rect 18732 13010 18788 13020
rect 18620 12126 18622 12178
rect 18674 12126 18676 12178
rect 18620 12114 18676 12126
rect 18732 12738 18788 12750
rect 18732 12686 18734 12738
rect 18786 12686 18788 12738
rect 18620 11844 18676 11854
rect 18732 11844 18788 12686
rect 18844 12738 18900 12750
rect 18844 12686 18846 12738
rect 18898 12686 18900 12738
rect 18844 12404 18900 12686
rect 18956 12740 19012 13356
rect 19068 12964 19124 13470
rect 19068 12870 19124 12908
rect 19292 12850 19348 12862
rect 19292 12798 19294 12850
rect 19346 12798 19348 12850
rect 19292 12740 19348 12798
rect 18956 12684 19348 12740
rect 18844 12338 18900 12348
rect 18956 12516 19012 12526
rect 18844 12180 18900 12190
rect 18956 12180 19012 12460
rect 19292 12402 19348 12684
rect 19516 12852 19572 14252
rect 19740 14242 19796 14252
rect 19836 14140 20100 14150
rect 19628 14084 19684 14094
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13188 19684 14028
rect 19964 13972 20020 13982
rect 19964 13878 20020 13916
rect 20188 13636 20244 14478
rect 20300 13972 20356 14700
rect 20300 13906 20356 13916
rect 20188 13570 20244 13580
rect 19740 13188 19796 13198
rect 19628 13186 19796 13188
rect 19628 13134 19742 13186
rect 19794 13134 19796 13186
rect 19628 13132 19796 13134
rect 19740 13122 19796 13132
rect 19292 12350 19294 12402
rect 19346 12350 19348 12402
rect 19292 12338 19348 12350
rect 19404 12404 19460 12414
rect 19404 12310 19460 12348
rect 18844 12178 19012 12180
rect 18844 12126 18846 12178
rect 18898 12126 19012 12178
rect 18844 12124 19012 12126
rect 19068 12180 19124 12190
rect 19068 12178 19236 12180
rect 19068 12126 19070 12178
rect 19122 12126 19236 12178
rect 19068 12124 19236 12126
rect 18844 12114 18900 12124
rect 19068 12114 19124 12124
rect 18508 11788 18620 11844
rect 18676 11788 18788 11844
rect 19068 11956 19124 11966
rect 18620 11778 18676 11788
rect 18844 11620 18900 11630
rect 19068 11620 19124 11900
rect 19180 11732 19236 12124
rect 19516 11956 19572 12796
rect 19628 12850 19684 12862
rect 19628 12798 19630 12850
rect 19682 12798 19684 12850
rect 19628 12180 19684 12798
rect 19740 12740 19796 12778
rect 19740 12674 19796 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19964 12180 20020 12190
rect 19628 12178 19796 12180
rect 19628 12126 19630 12178
rect 19682 12126 19796 12178
rect 19628 12124 19796 12126
rect 19628 12114 19684 12124
rect 19516 11890 19572 11900
rect 19180 11676 19684 11732
rect 19068 11564 19236 11620
rect 18844 11526 18900 11564
rect 18732 11508 18788 11518
rect 18620 11396 18676 11406
rect 18396 11394 18676 11396
rect 18396 11342 18622 11394
rect 18674 11342 18676 11394
rect 18396 11340 18676 11342
rect 17948 11284 18004 11294
rect 17948 11190 18004 11228
rect 17836 11170 17892 11182
rect 17836 11118 17838 11170
rect 17890 11118 17892 11170
rect 17836 10724 17892 11118
rect 17948 10724 18004 10734
rect 17836 10722 18004 10724
rect 17836 10670 17950 10722
rect 18002 10670 18004 10722
rect 17836 10668 18004 10670
rect 17948 10658 18004 10668
rect 17724 10610 17780 10622
rect 17724 10558 17726 10610
rect 17778 10558 17780 10610
rect 17388 9604 17444 9614
rect 17724 9604 17780 10558
rect 18060 9714 18116 11340
rect 18620 11330 18676 11340
rect 18172 11170 18228 11182
rect 18172 11118 18174 11170
rect 18226 11118 18228 11170
rect 18172 11060 18228 11118
rect 18172 10994 18228 11004
rect 18620 10724 18676 10734
rect 18732 10724 18788 11452
rect 19068 11396 19124 11406
rect 18844 11340 19068 11396
rect 18844 10834 18900 11340
rect 19068 11302 19124 11340
rect 18844 10782 18846 10834
rect 18898 10782 18900 10834
rect 18844 10770 18900 10782
rect 18956 11170 19012 11182
rect 18956 11118 18958 11170
rect 19010 11118 19012 11170
rect 18620 10722 18788 10724
rect 18620 10670 18622 10722
rect 18674 10670 18788 10722
rect 18620 10668 18788 10670
rect 18620 10658 18676 10668
rect 18396 10610 18452 10622
rect 18396 10558 18398 10610
rect 18450 10558 18452 10610
rect 18172 10500 18228 10510
rect 18172 10498 18340 10500
rect 18172 10446 18174 10498
rect 18226 10446 18340 10498
rect 18172 10444 18340 10446
rect 18172 10434 18228 10444
rect 18060 9662 18062 9714
rect 18114 9662 18116 9714
rect 18060 9650 18116 9662
rect 17388 9602 17780 9604
rect 17388 9550 17390 9602
rect 17442 9550 17780 9602
rect 17388 9548 17780 9550
rect 17388 9492 17444 9548
rect 17388 9426 17444 9436
rect 18284 9044 18340 10444
rect 18396 10388 18452 10558
rect 18732 10388 18788 10398
rect 18396 10386 18788 10388
rect 18396 10334 18734 10386
rect 18786 10334 18788 10386
rect 18396 10332 18788 10334
rect 18732 10322 18788 10332
rect 18396 9716 18452 9726
rect 18396 9622 18452 9660
rect 18732 9602 18788 9614
rect 18732 9550 18734 9602
rect 18786 9550 18788 9602
rect 18284 8988 18676 9044
rect 18620 8370 18676 8988
rect 18620 8318 18622 8370
rect 18674 8318 18676 8370
rect 18620 8306 18676 8318
rect 18732 8372 18788 9550
rect 18732 8306 18788 8316
rect 17276 8204 18004 8260
rect 17724 7700 17780 7710
rect 17724 7606 17780 7644
rect 17948 7588 18004 8204
rect 18956 7700 19012 11118
rect 19068 10836 19124 10846
rect 19180 10836 19236 11564
rect 19068 10834 19236 10836
rect 19068 10782 19070 10834
rect 19122 10782 19236 10834
rect 19068 10780 19236 10782
rect 19404 11508 19460 11518
rect 19404 11394 19460 11452
rect 19404 11342 19406 11394
rect 19458 11342 19460 11394
rect 19404 10836 19460 11342
rect 19628 11394 19684 11676
rect 19628 11342 19630 11394
rect 19682 11342 19684 11394
rect 19628 11330 19684 11342
rect 19740 11172 19796 12124
rect 19964 12178 20132 12180
rect 19964 12126 19966 12178
rect 20018 12126 20132 12178
rect 19964 12124 20132 12126
rect 19964 12114 20020 12124
rect 19964 11396 20020 11406
rect 19964 11302 20020 11340
rect 19852 11172 19908 11182
rect 19628 11170 19908 11172
rect 19628 11118 19854 11170
rect 19906 11118 19908 11170
rect 19628 11116 19908 11118
rect 20076 11172 20132 12124
rect 20748 11396 20804 11406
rect 20076 11116 20244 11172
rect 19068 10770 19124 10780
rect 19404 10770 19460 10780
rect 19516 11060 19572 11070
rect 19628 11060 19684 11116
rect 19852 11106 19908 11116
rect 19572 11004 19684 11060
rect 20188 11060 20244 11116
rect 19836 11004 20100 11014
rect 20188 11004 20356 11060
rect 19068 9716 19124 9726
rect 19516 9716 19572 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19740 10836 19796 10846
rect 19740 10742 19796 10780
rect 20188 10836 20244 10846
rect 20188 10742 20244 10780
rect 19068 9714 19572 9716
rect 19068 9662 19070 9714
rect 19122 9662 19572 9714
rect 19068 9660 19572 9662
rect 19628 10612 19684 10622
rect 20300 10612 20356 11004
rect 19068 9650 19124 9660
rect 19628 8484 19684 10556
rect 20076 10556 20356 10612
rect 20076 9716 20132 10556
rect 20076 9650 20132 9660
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19404 8428 19908 8484
rect 19404 8258 19460 8428
rect 19852 8370 19908 8428
rect 19852 8318 19854 8370
rect 19906 8318 19908 8370
rect 19852 8306 19908 8318
rect 19404 8206 19406 8258
rect 19458 8206 19460 8258
rect 19404 8194 19460 8206
rect 20748 8260 20804 11340
rect 21196 10612 21252 10622
rect 21196 10518 21252 10556
rect 20748 8194 20804 8204
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 17836 6690 17892 6702
rect 17836 6638 17838 6690
rect 17890 6638 17892 6690
rect 16940 6300 17220 6356
rect 17500 6466 17556 6478
rect 17836 6468 17892 6638
rect 17500 6414 17502 6466
rect 17554 6414 17556 6466
rect 16940 6132 16996 6300
rect 16156 5854 16158 5906
rect 16210 5854 16212 5906
rect 16156 5842 16212 5854
rect 16492 6130 16996 6132
rect 16492 6078 16942 6130
rect 16994 6078 16996 6130
rect 16492 6076 16996 6078
rect 16492 5906 16548 6076
rect 16940 6066 16996 6076
rect 16492 5854 16494 5906
rect 16546 5854 16548 5906
rect 16492 5842 16548 5854
rect 17388 5908 17444 5918
rect 17500 5908 17556 6414
rect 17444 5852 17556 5908
rect 17724 6412 17836 6468
rect 17388 5814 17444 5852
rect 16268 5796 16324 5806
rect 16268 5702 16324 5740
rect 17612 5796 17668 5806
rect 17612 5702 17668 5740
rect 15148 5628 15876 5684
rect 16268 5236 16324 5246
rect 16268 5142 16324 5180
rect 17612 5236 17668 5246
rect 17724 5236 17780 6412
rect 17836 6402 17892 6412
rect 17948 6132 18004 7532
rect 18620 7644 19012 7700
rect 20748 7700 20804 7710
rect 21308 7700 21364 15092
rect 21420 13636 21476 13646
rect 21420 12404 21476 13580
rect 21420 12310 21476 12348
rect 21980 12964 22036 12974
rect 21756 12178 21812 12190
rect 21756 12126 21758 12178
rect 21810 12126 21812 12178
rect 21644 11284 21700 11294
rect 21532 11228 21644 11284
rect 21420 7700 21476 7710
rect 20748 7698 21476 7700
rect 20748 7646 20750 7698
rect 20802 7646 21422 7698
rect 21474 7646 21476 7698
rect 20748 7644 21476 7646
rect 18620 6690 18676 7644
rect 20748 7634 20804 7644
rect 21420 7634 21476 7644
rect 20972 7476 21028 7486
rect 20860 7420 20972 7476
rect 20748 6804 20804 6814
rect 20860 6804 20916 7420
rect 20972 7382 21028 7420
rect 21084 7476 21140 7486
rect 21532 7476 21588 11228
rect 21644 11190 21700 11228
rect 21756 11172 21812 12126
rect 21868 11396 21924 11406
rect 21980 11396 22036 12908
rect 21924 11340 22036 11396
rect 22092 11396 22148 16380
rect 22540 16100 22596 16716
rect 22204 15988 22260 15998
rect 22204 15540 22260 15932
rect 22428 15988 22484 15998
rect 22428 15894 22484 15932
rect 22204 15474 22260 15484
rect 22540 14530 22596 16044
rect 22540 14478 22542 14530
rect 22594 14478 22596 14530
rect 22540 14466 22596 14478
rect 22652 16322 22708 18060
rect 22876 17892 22932 17902
rect 22876 17554 22932 17836
rect 22876 17502 22878 17554
rect 22930 17502 22932 17554
rect 22876 17490 22932 17502
rect 22876 17108 22932 17118
rect 22876 17014 22932 17052
rect 22652 16270 22654 16322
rect 22706 16270 22708 16322
rect 22652 13860 22708 16270
rect 22540 13804 22708 13860
rect 22876 15876 22932 15886
rect 22876 14306 22932 15820
rect 22876 14254 22878 14306
rect 22930 14254 22932 14306
rect 22876 13860 22932 14254
rect 22988 14308 23044 21420
rect 23548 20692 23604 20702
rect 23436 20690 23604 20692
rect 23436 20638 23550 20690
rect 23602 20638 23604 20690
rect 23436 20636 23604 20638
rect 23100 20020 23156 20030
rect 23100 19926 23156 19964
rect 23212 19794 23268 19806
rect 23212 19742 23214 19794
rect 23266 19742 23268 19794
rect 23212 19458 23268 19742
rect 23212 19406 23214 19458
rect 23266 19406 23268 19458
rect 23212 19394 23268 19406
rect 23436 19346 23492 20636
rect 23548 20626 23604 20636
rect 23660 19460 23716 23324
rect 23884 23044 23940 23054
rect 23884 22950 23940 22988
rect 23772 20132 23828 20142
rect 23772 20018 23828 20076
rect 23772 19966 23774 20018
rect 23826 19966 23828 20018
rect 23772 19954 23828 19966
rect 24220 20018 24276 20030
rect 24220 19966 24222 20018
rect 24274 19966 24276 20018
rect 23996 19908 24052 19918
rect 23996 19814 24052 19852
rect 24220 19908 24276 19966
rect 24444 20020 24500 20030
rect 24444 19926 24500 19964
rect 24220 19842 24276 19852
rect 23660 19394 23716 19404
rect 23436 19294 23438 19346
rect 23490 19294 23492 19346
rect 23436 19282 23492 19294
rect 23548 19234 23604 19246
rect 23548 19182 23550 19234
rect 23602 19182 23604 19234
rect 23100 19124 23156 19134
rect 23100 19122 23380 19124
rect 23100 19070 23102 19122
rect 23154 19070 23380 19122
rect 23100 19068 23380 19070
rect 23100 19058 23156 19068
rect 23212 18788 23268 18798
rect 23100 17668 23156 17678
rect 23100 16772 23156 17612
rect 23212 17666 23268 18732
rect 23212 17614 23214 17666
rect 23266 17614 23268 17666
rect 23212 17220 23268 17614
rect 23212 17154 23268 17164
rect 23324 17892 23380 19068
rect 23548 18564 23604 19182
rect 23548 18498 23604 18508
rect 24556 18564 24612 18574
rect 23436 17892 23492 17902
rect 23324 17890 23492 17892
rect 23324 17838 23438 17890
rect 23490 17838 23492 17890
rect 23324 17836 23492 17838
rect 23212 16996 23268 17006
rect 23324 16996 23380 17836
rect 23436 17826 23492 17836
rect 23772 17892 23828 17902
rect 23772 17666 23828 17836
rect 23772 17614 23774 17666
rect 23826 17614 23828 17666
rect 23772 17602 23828 17614
rect 23436 17556 23492 17566
rect 23436 17106 23492 17500
rect 23996 17554 24052 17566
rect 23996 17502 23998 17554
rect 24050 17502 24052 17554
rect 23436 17054 23438 17106
rect 23490 17054 23492 17106
rect 23436 17042 23492 17054
rect 23660 17442 23716 17454
rect 23660 17390 23662 17442
rect 23714 17390 23716 17442
rect 23212 16994 23380 16996
rect 23212 16942 23214 16994
rect 23266 16942 23380 16994
rect 23212 16940 23380 16942
rect 23548 16996 23604 17006
rect 23212 16930 23268 16940
rect 23548 16902 23604 16940
rect 23660 16882 23716 17390
rect 23660 16830 23662 16882
rect 23714 16830 23716 16882
rect 23660 16818 23716 16830
rect 23996 16772 24052 17502
rect 24332 17556 24388 17566
rect 24332 17462 24388 17500
rect 24556 17554 24612 18508
rect 24556 17502 24558 17554
rect 24610 17502 24612 17554
rect 24556 17490 24612 17502
rect 24444 17444 24500 17454
rect 24444 17350 24500 17388
rect 24556 16994 24612 17006
rect 24556 16942 24558 16994
rect 24610 16942 24612 16994
rect 24108 16884 24164 16894
rect 24108 16790 24164 16828
rect 24332 16882 24388 16894
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 23100 16716 23268 16772
rect 23212 16098 23268 16716
rect 23212 16046 23214 16098
rect 23266 16046 23268 16098
rect 23212 16034 23268 16046
rect 23772 16716 24052 16772
rect 23772 16100 23828 16716
rect 24220 16660 24276 16670
rect 23100 15986 23156 15998
rect 23100 15934 23102 15986
rect 23154 15934 23156 15986
rect 23100 15876 23156 15934
rect 23324 15988 23380 15998
rect 23324 15894 23380 15932
rect 23100 15810 23156 15820
rect 23436 15876 23492 15886
rect 23100 15540 23156 15550
rect 23100 15446 23156 15484
rect 23436 15538 23492 15820
rect 23436 15486 23438 15538
rect 23490 15486 23492 15538
rect 23436 15474 23492 15486
rect 23772 15540 23828 16044
rect 23884 16658 24276 16660
rect 23884 16606 24222 16658
rect 24274 16606 24276 16658
rect 23884 16604 24276 16606
rect 23884 15986 23940 16604
rect 24220 16594 24276 16604
rect 23884 15934 23886 15986
rect 23938 15934 23940 15986
rect 23884 15922 23940 15934
rect 23996 15876 24052 15886
rect 23996 15782 24052 15820
rect 23772 15474 23828 15484
rect 24332 15538 24388 16830
rect 24556 16884 24612 16942
rect 24556 16818 24612 16828
rect 24668 16324 24724 24668
rect 24892 17108 24948 29934
rect 25228 27074 25284 27086
rect 25228 27022 25230 27074
rect 25282 27022 25284 27074
rect 25228 26180 25284 27022
rect 25676 27076 25732 27086
rect 25004 23940 25060 23950
rect 25004 23846 25060 23884
rect 25228 21812 25284 26124
rect 25452 26290 25508 26302
rect 25452 26238 25454 26290
rect 25506 26238 25508 26290
rect 25452 25620 25508 26238
rect 25340 21812 25396 21822
rect 25228 21810 25396 21812
rect 25228 21758 25342 21810
rect 25394 21758 25396 21810
rect 25228 21756 25396 21758
rect 25228 21364 25284 21374
rect 25228 20804 25284 21308
rect 25116 20748 25284 20804
rect 25116 17780 25172 20748
rect 25228 20580 25284 20590
rect 25228 19348 25284 20524
rect 25340 20244 25396 21756
rect 25340 20178 25396 20188
rect 25452 20356 25508 25564
rect 25564 24724 25620 24734
rect 25564 24630 25620 24668
rect 25452 20020 25508 20300
rect 25564 24164 25620 24174
rect 25564 20244 25620 24108
rect 25676 21364 25732 27020
rect 25788 26178 25844 30604
rect 26124 30210 26180 30222
rect 26124 30158 26126 30210
rect 26178 30158 26180 30210
rect 25900 28644 25956 28654
rect 25900 27186 25956 28588
rect 26124 28532 26180 30158
rect 26236 29988 26292 31164
rect 26460 30322 26516 32508
rect 27468 32562 27524 32574
rect 27468 32510 27470 32562
rect 27522 32510 27524 32562
rect 27468 30772 27524 32510
rect 28028 32564 28084 33964
rect 28140 33954 28196 33964
rect 28812 34018 28868 34030
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 28812 33348 28868 33966
rect 29148 33348 29204 33358
rect 28812 33346 29204 33348
rect 28812 33294 29150 33346
rect 29202 33294 29204 33346
rect 28812 33292 29204 33294
rect 28588 33234 28644 33246
rect 28588 33182 28590 33234
rect 28642 33182 28644 33234
rect 28140 33122 28196 33134
rect 28140 33070 28142 33122
rect 28194 33070 28196 33122
rect 28140 32900 28196 33070
rect 28252 33124 28308 33134
rect 28252 33030 28308 33068
rect 28476 33122 28532 33134
rect 28476 33070 28478 33122
rect 28530 33070 28532 33122
rect 28476 32900 28532 33070
rect 28140 32844 28532 32900
rect 28140 32564 28196 32574
rect 28028 32508 28140 32564
rect 28140 32470 28196 32508
rect 27468 30706 27524 30716
rect 27580 32452 27636 32462
rect 26460 30270 26462 30322
rect 26514 30270 26516 30322
rect 26460 30258 26516 30270
rect 26236 29922 26292 29932
rect 26348 30212 26404 30222
rect 26348 29538 26404 30156
rect 27468 30212 27524 30222
rect 27468 30118 27524 30156
rect 27020 30098 27076 30110
rect 27020 30046 27022 30098
rect 27074 30046 27076 30098
rect 26348 29486 26350 29538
rect 26402 29486 26404 29538
rect 26348 29474 26404 29486
rect 26460 29988 26516 29998
rect 26460 29538 26516 29932
rect 26796 29652 26852 29662
rect 26796 29558 26852 29596
rect 26460 29486 26462 29538
rect 26514 29486 26516 29538
rect 26460 29474 26516 29486
rect 26572 29538 26628 29550
rect 26572 29486 26574 29538
rect 26626 29486 26628 29538
rect 26572 29428 26628 29486
rect 26684 29540 26740 29550
rect 26684 29446 26740 29484
rect 27020 29540 27076 30046
rect 27356 30100 27412 30110
rect 27356 30006 27412 30044
rect 27132 29988 27188 29998
rect 27188 29932 27300 29988
rect 27132 29922 27188 29932
rect 27020 29474 27076 29484
rect 26572 28644 26628 29372
rect 27132 29428 27188 29438
rect 27132 29334 27188 29372
rect 26572 28578 26628 28588
rect 25900 27134 25902 27186
rect 25954 27134 25956 27186
rect 25900 27122 25956 27134
rect 26012 28476 26180 28532
rect 27132 28532 27188 28542
rect 27244 28532 27300 29932
rect 27132 28530 27300 28532
rect 27132 28478 27134 28530
rect 27186 28478 27300 28530
rect 27132 28476 27300 28478
rect 27356 29652 27412 29662
rect 27356 29426 27412 29596
rect 27356 29374 27358 29426
rect 27410 29374 27412 29426
rect 25788 26126 25790 26178
rect 25842 26126 25844 26178
rect 25788 26114 25844 26126
rect 25788 25508 25844 25518
rect 25788 24610 25844 25452
rect 25788 24558 25790 24610
rect 25842 24558 25844 24610
rect 25788 24546 25844 24558
rect 26012 24164 26068 28476
rect 27132 28466 27188 28476
rect 26796 28420 26852 28430
rect 26684 28418 26852 28420
rect 26684 28366 26798 28418
rect 26850 28366 26852 28418
rect 26684 28364 26852 28366
rect 26236 27746 26292 27758
rect 26236 27694 26238 27746
rect 26290 27694 26292 27746
rect 26236 27076 26292 27694
rect 26684 27186 26740 28364
rect 26796 28354 26852 28364
rect 26908 28420 26964 28430
rect 26908 28326 26964 28364
rect 26684 27134 26686 27186
rect 26738 27134 26740 27186
rect 26684 27122 26740 27134
rect 26908 27860 26964 27870
rect 26236 27010 26292 27020
rect 26796 27076 26852 27086
rect 26796 26982 26852 27020
rect 26124 26962 26180 26974
rect 26124 26910 26126 26962
rect 26178 26910 26180 26962
rect 26124 26908 26180 26910
rect 26124 26852 26628 26908
rect 26572 26628 26628 26852
rect 26236 26292 26292 26302
rect 26012 24098 26068 24108
rect 26124 26066 26180 26078
rect 26124 26014 26126 26066
rect 26178 26014 26180 26066
rect 26124 25506 26180 26014
rect 26236 25618 26292 26236
rect 26236 25566 26238 25618
rect 26290 25566 26292 25618
rect 26236 25554 26292 25566
rect 26124 25454 26126 25506
rect 26178 25454 26180 25506
rect 26124 23940 26180 25454
rect 26572 25172 26628 26572
rect 26796 26290 26852 26302
rect 26796 26238 26798 26290
rect 26850 26238 26852 26290
rect 26684 25956 26740 25966
rect 26684 25394 26740 25900
rect 26796 25620 26852 26238
rect 26908 25844 26964 27804
rect 27356 27188 27412 29374
rect 27580 29428 27636 32396
rect 28476 31108 28532 32844
rect 28588 32004 28644 33182
rect 28588 31938 28644 31948
rect 28700 32674 28756 32686
rect 28700 32622 28702 32674
rect 28754 32622 28756 32674
rect 28700 31220 28756 32622
rect 28700 31154 28756 31164
rect 27804 30996 27860 31006
rect 27804 30434 27860 30940
rect 27804 30382 27806 30434
rect 27858 30382 27860 30434
rect 27804 30370 27860 30382
rect 27692 30322 27748 30334
rect 27692 30270 27694 30322
rect 27746 30270 27748 30322
rect 27692 29988 27748 30270
rect 28252 30212 28308 30222
rect 28308 30156 28420 30212
rect 28252 30146 28308 30156
rect 27692 29922 27748 29932
rect 28252 29650 28308 29662
rect 28252 29598 28254 29650
rect 28306 29598 28308 29650
rect 27580 29362 27636 29372
rect 27916 29426 27972 29438
rect 27916 29374 27918 29426
rect 27970 29374 27972 29426
rect 27692 29204 27748 29214
rect 27916 29204 27972 29374
rect 27692 29202 27972 29204
rect 27692 29150 27694 29202
rect 27746 29150 27972 29202
rect 27692 29148 27972 29150
rect 27468 28644 27524 28654
rect 27692 28644 27748 29148
rect 27468 28642 27748 28644
rect 27468 28590 27470 28642
rect 27522 28590 27748 28642
rect 27468 28588 27748 28590
rect 28028 28644 28084 28654
rect 27468 28532 27524 28588
rect 27468 28466 27524 28476
rect 27356 27132 27972 27188
rect 27356 26908 27412 27132
rect 27244 26852 27412 26908
rect 27468 26964 27524 26974
rect 27468 26962 27636 26964
rect 27468 26910 27470 26962
rect 27522 26910 27636 26962
rect 27468 26908 27636 26910
rect 27468 26898 27524 26908
rect 27580 26852 27748 26908
rect 27244 26514 27300 26852
rect 27244 26462 27246 26514
rect 27298 26462 27300 26514
rect 27244 26450 27300 26462
rect 27468 26628 27524 26638
rect 27468 26514 27524 26572
rect 27468 26462 27470 26514
rect 27522 26462 27524 26514
rect 27468 26450 27524 26462
rect 27020 26292 27076 26302
rect 27020 26198 27076 26236
rect 26908 25778 26964 25788
rect 27244 26178 27300 26190
rect 27244 26126 27246 26178
rect 27298 26126 27300 26178
rect 26796 25564 27076 25620
rect 26684 25342 26686 25394
rect 26738 25342 26740 25394
rect 26684 25330 26740 25342
rect 26572 25116 26740 25172
rect 26236 24724 26292 24734
rect 26236 24630 26292 24668
rect 26572 23940 26628 23950
rect 26124 23938 26628 23940
rect 26124 23886 26574 23938
rect 26626 23886 26628 23938
rect 26124 23884 26628 23886
rect 26572 23874 26628 23884
rect 26684 23826 26740 25116
rect 27020 24724 27076 25564
rect 27244 25506 27300 26126
rect 27244 25454 27246 25506
rect 27298 25454 27300 25506
rect 27244 25442 27300 25454
rect 27692 25506 27748 26852
rect 27804 26628 27860 26638
rect 27804 26402 27860 26572
rect 27916 26514 27972 27132
rect 27916 26462 27918 26514
rect 27970 26462 27972 26514
rect 27916 26450 27972 26462
rect 27804 26350 27806 26402
rect 27858 26350 27860 26402
rect 27804 26338 27860 26350
rect 27692 25454 27694 25506
rect 27746 25454 27748 25506
rect 27692 25442 27748 25454
rect 26908 24668 27076 24724
rect 27244 25282 27300 25294
rect 27244 25230 27246 25282
rect 27298 25230 27300 25282
rect 26908 24164 26964 24668
rect 26684 23774 26686 23826
rect 26738 23774 26740 23826
rect 26684 23762 26740 23774
rect 26796 24108 26964 24164
rect 27020 24498 27076 24510
rect 27020 24446 27022 24498
rect 27074 24446 27076 24498
rect 26796 21924 26852 24108
rect 26908 23828 26964 23838
rect 26908 23734 26964 23772
rect 27020 23492 27076 24446
rect 27132 24498 27188 24510
rect 27132 24446 27134 24498
rect 27186 24446 27188 24498
rect 27132 23828 27188 24446
rect 27244 24052 27300 25230
rect 27356 25172 27412 25182
rect 27356 24722 27412 25116
rect 27804 24836 27860 24846
rect 27356 24670 27358 24722
rect 27410 24670 27412 24722
rect 27356 24658 27412 24670
rect 27580 24834 27860 24836
rect 27580 24782 27806 24834
rect 27858 24782 27860 24834
rect 27580 24780 27860 24782
rect 27580 24722 27636 24780
rect 27804 24770 27860 24780
rect 27916 24836 27972 24846
rect 28028 24836 28084 28588
rect 28140 28642 28196 28654
rect 28140 28590 28142 28642
rect 28194 28590 28196 28642
rect 28140 28532 28196 28590
rect 28140 27188 28196 28476
rect 28252 28084 28308 29598
rect 28364 29538 28420 30156
rect 28476 30100 28532 31052
rect 28476 30034 28532 30044
rect 28364 29486 28366 29538
rect 28418 29486 28420 29538
rect 28364 29474 28420 29486
rect 28476 29540 28532 29550
rect 28476 29426 28532 29484
rect 28476 29374 28478 29426
rect 28530 29374 28532 29426
rect 28364 28644 28420 28654
rect 28476 28644 28532 29374
rect 28420 28588 28532 28644
rect 28364 28550 28420 28588
rect 28700 28532 28756 28542
rect 28700 28438 28756 28476
rect 28588 28420 28644 28430
rect 28588 28326 28644 28364
rect 28252 28028 28420 28084
rect 28252 27860 28308 27870
rect 28252 27766 28308 27804
rect 28140 27122 28196 27132
rect 28140 26290 28196 26302
rect 28140 26238 28142 26290
rect 28194 26238 28196 26290
rect 28140 25060 28196 26238
rect 28252 26068 28308 26078
rect 28252 25974 28308 26012
rect 28140 24994 28196 25004
rect 28252 25844 28308 25854
rect 27916 24834 28084 24836
rect 27916 24782 27918 24834
rect 27970 24782 28084 24834
rect 27916 24780 28084 24782
rect 28140 24836 28196 24846
rect 28252 24836 28308 25788
rect 28364 25394 28420 28028
rect 29148 27860 29204 33292
rect 29260 32788 29316 34078
rect 29260 32722 29316 32732
rect 29484 32564 29540 32574
rect 29484 32470 29540 32508
rect 29596 32452 29652 34190
rect 30268 34188 30548 34244
rect 29932 34130 29988 34142
rect 29932 34078 29934 34130
rect 29986 34078 29988 34130
rect 29932 34020 29988 34078
rect 30268 34130 30324 34188
rect 30268 34078 30270 34130
rect 30322 34078 30324 34130
rect 30268 34066 30324 34078
rect 29932 33954 29988 33964
rect 30380 34018 30436 34030
rect 30380 33966 30382 34018
rect 30434 33966 30436 34018
rect 30380 33684 30436 33966
rect 30156 33628 30436 33684
rect 29820 33124 29876 33134
rect 29820 32562 29876 33068
rect 29820 32510 29822 32562
rect 29874 32510 29876 32562
rect 29820 32498 29876 32510
rect 30156 32562 30212 33628
rect 30492 32900 30548 34188
rect 30828 34150 30884 34188
rect 30604 34132 30660 34142
rect 30604 34130 30772 34132
rect 30604 34078 30606 34130
rect 30658 34078 30772 34130
rect 30604 34076 30772 34078
rect 30604 34066 30660 34076
rect 30492 32844 30660 32900
rect 30380 32788 30436 32798
rect 30380 32694 30436 32732
rect 30604 32788 30660 32844
rect 30156 32510 30158 32562
rect 30210 32510 30212 32562
rect 30156 32498 30212 32510
rect 30268 32562 30324 32574
rect 30268 32510 30270 32562
rect 30322 32510 30324 32562
rect 29596 32386 29652 32396
rect 30268 32452 30324 32510
rect 30268 32386 30324 32396
rect 30492 32564 30548 32574
rect 29708 31220 29764 31230
rect 29708 31126 29764 31164
rect 29932 31108 29988 31118
rect 30268 31108 30324 31118
rect 29932 31106 30324 31108
rect 29932 31054 29934 31106
rect 29986 31054 30270 31106
rect 30322 31054 30324 31106
rect 29932 31052 30324 31054
rect 29932 31042 29988 31052
rect 30268 31042 30324 31052
rect 29596 30994 29652 31006
rect 29596 30942 29598 30994
rect 29650 30942 29652 30994
rect 29596 30212 29652 30942
rect 30380 30994 30436 31006
rect 30380 30942 30382 30994
rect 30434 30942 30436 30994
rect 30268 30772 30324 30782
rect 30268 30678 30324 30716
rect 30156 30324 30212 30334
rect 29932 30212 29988 30222
rect 29596 30210 30100 30212
rect 29596 30158 29934 30210
rect 29986 30158 30100 30210
rect 29596 30156 30100 30158
rect 29932 30146 29988 30156
rect 29820 28868 29876 28878
rect 29148 27794 29204 27804
rect 29260 28866 29876 28868
rect 29260 28814 29822 28866
rect 29874 28814 29876 28866
rect 29260 28812 29876 28814
rect 29260 27300 29316 28812
rect 29820 28802 29876 28812
rect 29708 28532 29764 28542
rect 29708 28438 29764 28476
rect 29820 28420 29876 28430
rect 30044 28420 30100 30156
rect 30156 30098 30212 30268
rect 30380 30212 30436 30942
rect 30380 30146 30436 30156
rect 30156 30046 30158 30098
rect 30210 30046 30212 30098
rect 30156 30034 30212 30046
rect 30492 29988 30548 32508
rect 30604 31780 30660 32732
rect 30604 31714 30660 31724
rect 30716 31556 30772 34076
rect 31052 34020 31108 35534
rect 31500 35586 31556 35598
rect 31500 35534 31502 35586
rect 31554 35534 31556 35586
rect 31052 33954 31108 33964
rect 31164 35028 31220 35038
rect 31500 35028 31556 35534
rect 31220 34972 31556 35028
rect 33740 35028 33796 36204
rect 35084 35812 35140 35822
rect 33740 34972 34356 35028
rect 31164 34132 31220 34972
rect 31164 33458 31220 34076
rect 31724 34916 31780 34926
rect 31724 34130 31780 34860
rect 34076 34804 34132 34814
rect 33964 34802 34132 34804
rect 33964 34750 34078 34802
rect 34130 34750 34132 34802
rect 33964 34748 34132 34750
rect 31724 34078 31726 34130
rect 31778 34078 31780 34130
rect 31724 34066 31780 34078
rect 32172 34244 32228 34254
rect 31164 33406 31166 33458
rect 31218 33406 31220 33458
rect 31164 33394 31220 33406
rect 31276 34020 31332 34030
rect 31276 32562 31332 33964
rect 31276 32510 31278 32562
rect 31330 32510 31332 32562
rect 31276 32498 31332 32510
rect 31836 32564 31892 32574
rect 31836 32470 31892 32508
rect 32060 32564 32116 32574
rect 32172 32564 32228 34188
rect 33180 33348 33236 33358
rect 32956 32788 33012 32798
rect 32956 32694 33012 32732
rect 33180 32786 33236 33292
rect 33180 32734 33182 32786
rect 33234 32734 33236 32786
rect 32060 32562 32228 32564
rect 32060 32510 32062 32562
rect 32114 32510 32228 32562
rect 32060 32508 32228 32510
rect 31500 32452 31556 32462
rect 31388 32450 31556 32452
rect 31388 32398 31502 32450
rect 31554 32398 31556 32450
rect 31388 32396 31556 32398
rect 30940 32338 30996 32350
rect 30940 32286 30942 32338
rect 30994 32286 30996 32338
rect 30828 32004 30884 32042
rect 30828 31938 30884 31948
rect 30940 31948 30996 32286
rect 31388 32116 31444 32396
rect 31500 32386 31556 32396
rect 32060 32228 32116 32508
rect 31388 32050 31444 32060
rect 31500 32172 32116 32228
rect 32284 32452 32340 32462
rect 30940 31892 31332 31948
rect 30940 31780 30996 31790
rect 31164 31780 31220 31790
rect 30996 31778 31220 31780
rect 30996 31726 31166 31778
rect 31218 31726 31220 31778
rect 30996 31724 31220 31726
rect 30940 31714 30996 31724
rect 31164 31714 31220 31724
rect 31276 31780 31332 31892
rect 31276 31714 31332 31724
rect 31500 31778 31556 32172
rect 31500 31726 31502 31778
rect 31554 31726 31556 31778
rect 31500 31714 31556 31726
rect 31724 31780 31780 31790
rect 30940 31556 30996 31566
rect 31612 31556 31668 31566
rect 30716 31554 31668 31556
rect 30716 31502 30942 31554
rect 30994 31502 31614 31554
rect 31666 31502 31668 31554
rect 30716 31500 31668 31502
rect 30940 31490 30996 31500
rect 31612 31490 31668 31500
rect 30940 31332 30996 31342
rect 30940 30210 30996 31276
rect 31724 30996 31780 31724
rect 31948 31780 32004 31790
rect 31836 31554 31892 31566
rect 31836 31502 31838 31554
rect 31890 31502 31892 31554
rect 31836 31220 31892 31502
rect 31836 31154 31892 31164
rect 31836 30996 31892 31006
rect 31724 30940 31836 30996
rect 31836 30902 31892 30940
rect 31948 30660 32004 31724
rect 32284 31218 32340 32396
rect 33180 32452 33236 32734
rect 33292 32564 33348 32574
rect 33964 32564 34020 34748
rect 34076 34738 34132 34748
rect 34076 34132 34132 34142
rect 34076 33572 34132 34076
rect 34076 33506 34132 33516
rect 34076 32564 34132 32574
rect 33964 32508 34076 32564
rect 33292 32470 33348 32508
rect 34076 32498 34132 32508
rect 33180 32386 33236 32396
rect 32284 31166 32286 31218
rect 32338 31166 32340 31218
rect 32284 31154 32340 31166
rect 32396 32338 32452 32350
rect 32396 32286 32398 32338
rect 32450 32286 32452 32338
rect 32060 30996 32116 31006
rect 32060 30902 32116 30940
rect 32396 30994 32452 32286
rect 34188 32338 34244 32350
rect 34188 32286 34190 32338
rect 34242 32286 34244 32338
rect 34076 31668 34132 31678
rect 33180 31220 33236 31230
rect 33180 31126 33236 31164
rect 32396 30942 32398 30994
rect 32450 30942 32452 30994
rect 32396 30930 32452 30942
rect 33404 30996 33460 31006
rect 33404 30902 33460 30940
rect 31948 30594 32004 30604
rect 32172 30882 32228 30894
rect 32172 30830 32174 30882
rect 32226 30830 32228 30882
rect 32172 30436 32228 30830
rect 31612 30434 32228 30436
rect 31612 30382 32174 30434
rect 32226 30382 32228 30434
rect 31612 30380 32228 30382
rect 30940 30158 30942 30210
rect 30994 30158 30996 30210
rect 30940 30146 30996 30158
rect 31164 30324 31220 30334
rect 31164 30210 31220 30268
rect 31164 30158 31166 30210
rect 31218 30158 31220 30210
rect 31164 30146 31220 30158
rect 31388 30212 31444 30222
rect 31388 30118 31444 30156
rect 31500 30210 31556 30222
rect 31500 30158 31502 30210
rect 31554 30158 31556 30210
rect 29820 28418 29988 28420
rect 29820 28366 29822 28418
rect 29874 28366 29988 28418
rect 29820 28364 29988 28366
rect 29820 28354 29876 28364
rect 29932 27748 29988 28364
rect 30044 28354 30100 28364
rect 30380 29932 30548 29988
rect 31276 29986 31332 29998
rect 31276 29934 31278 29986
rect 31330 29934 31332 29986
rect 30268 27972 30324 27982
rect 30380 27972 30436 29932
rect 31164 29540 31220 29550
rect 30940 29426 30996 29438
rect 30940 29374 30942 29426
rect 30994 29374 30996 29426
rect 30604 29316 30660 29326
rect 30940 29316 30996 29374
rect 30604 29314 30996 29316
rect 30604 29262 30606 29314
rect 30658 29262 30996 29314
rect 30604 29260 30996 29262
rect 30492 28420 30548 28430
rect 30492 28326 30548 28364
rect 30324 27916 30436 27972
rect 30268 27906 30324 27916
rect 29932 27692 30212 27748
rect 28924 27244 29316 27300
rect 30044 27300 30100 27310
rect 28924 26290 28980 27244
rect 29372 27188 29428 27198
rect 29372 27094 29428 27132
rect 28924 26238 28926 26290
rect 28978 26238 28980 26290
rect 28924 26226 28980 26238
rect 29484 27074 29540 27086
rect 29484 27022 29486 27074
rect 29538 27022 29540 27074
rect 29148 26178 29204 26190
rect 29148 26126 29150 26178
rect 29202 26126 29204 26178
rect 28364 25342 28366 25394
rect 28418 25342 28420 25394
rect 28364 25330 28420 25342
rect 28700 26066 28756 26078
rect 28700 26014 28702 26066
rect 28754 26014 28756 26066
rect 28700 25284 28756 26014
rect 28700 25228 29092 25284
rect 28924 25060 28980 25070
rect 28140 24834 28308 24836
rect 28140 24782 28142 24834
rect 28194 24782 28308 24834
rect 28140 24780 28308 24782
rect 28364 24836 28420 24846
rect 27916 24770 27972 24780
rect 28140 24770 28196 24780
rect 28364 24742 28420 24780
rect 28924 24834 28980 25004
rect 28924 24782 28926 24834
rect 28978 24782 28980 24834
rect 28924 24770 28980 24782
rect 27580 24670 27582 24722
rect 27634 24670 27636 24722
rect 27580 24658 27636 24670
rect 28588 24724 28644 24734
rect 28588 24630 28644 24668
rect 29036 24610 29092 25228
rect 29148 25172 29204 26126
rect 29484 25844 29540 27022
rect 30044 26908 30100 27244
rect 30156 27186 30212 27692
rect 30156 27134 30158 27186
rect 30210 27134 30212 27186
rect 30156 27122 30212 27134
rect 30380 26908 30436 27916
rect 30044 26852 30212 26908
rect 30380 26852 30548 26908
rect 29484 25778 29540 25788
rect 29708 26178 29764 26190
rect 29708 26126 29710 26178
rect 29762 26126 29764 26178
rect 29708 25508 29764 26126
rect 30156 25618 30212 26852
rect 30156 25566 30158 25618
rect 30210 25566 30212 25618
rect 30156 25554 30212 25566
rect 30044 25508 30100 25518
rect 29708 25506 30100 25508
rect 29708 25454 30046 25506
rect 30098 25454 30100 25506
rect 29708 25452 30100 25454
rect 29148 25106 29204 25116
rect 29372 25394 29428 25406
rect 29372 25342 29374 25394
rect 29426 25342 29428 25394
rect 29372 24836 29428 25342
rect 30044 24948 30100 25452
rect 30044 24892 30212 24948
rect 29372 24742 29428 24780
rect 29148 24724 29204 24734
rect 29708 24724 29764 24734
rect 29148 24722 29316 24724
rect 29148 24670 29150 24722
rect 29202 24670 29316 24722
rect 29148 24668 29316 24670
rect 29148 24658 29204 24668
rect 29036 24558 29038 24610
rect 29090 24558 29092 24610
rect 29036 24546 29092 24558
rect 29260 24612 29316 24668
rect 29708 24630 29764 24668
rect 30044 24722 30100 24734
rect 30044 24670 30046 24722
rect 30098 24670 30100 24722
rect 29260 24556 29652 24612
rect 29596 24500 29652 24556
rect 29820 24610 29876 24622
rect 29820 24558 29822 24610
rect 29874 24558 29876 24610
rect 29820 24500 29876 24558
rect 29596 24444 29876 24500
rect 27244 23996 27748 24052
rect 27132 23762 27188 23772
rect 27020 23436 27412 23492
rect 26908 23268 26964 23278
rect 26964 23212 27300 23268
rect 26908 23174 26964 23212
rect 27244 23154 27300 23212
rect 27244 23102 27246 23154
rect 27298 23102 27300 23154
rect 27244 23090 27300 23102
rect 26572 21868 26852 21924
rect 25900 21588 25956 21598
rect 26348 21588 26404 21598
rect 25900 21494 25956 21532
rect 26012 21586 26404 21588
rect 26012 21534 26350 21586
rect 26402 21534 26404 21586
rect 26012 21532 26404 21534
rect 25676 21298 25732 21308
rect 26012 21028 26068 21532
rect 25676 20972 26068 21028
rect 26124 21140 26180 21150
rect 25676 20914 25732 20972
rect 25676 20862 25678 20914
rect 25730 20862 25732 20914
rect 25676 20850 25732 20862
rect 26012 20692 26068 20702
rect 26012 20598 26068 20636
rect 25900 20356 25956 20366
rect 26124 20356 26180 21084
rect 25564 20188 25844 20244
rect 25228 19282 25284 19292
rect 25340 19964 25508 20020
rect 25116 17778 25284 17780
rect 25116 17726 25118 17778
rect 25170 17726 25284 17778
rect 25116 17724 25284 17726
rect 25116 17714 25172 17724
rect 24892 17042 24948 17052
rect 25228 16996 25284 17724
rect 25228 16902 25284 16940
rect 24332 15486 24334 15538
rect 24386 15486 24388 15538
rect 23884 15316 23940 15326
rect 23772 15260 23884 15316
rect 23772 15202 23828 15260
rect 23884 15250 23940 15260
rect 23772 15150 23774 15202
rect 23826 15150 23828 15202
rect 23772 15138 23828 15150
rect 24332 15148 24388 15486
rect 23884 15092 24388 15148
rect 24444 16098 24500 16110
rect 24444 16046 24446 16098
rect 24498 16046 24500 16098
rect 23884 14754 23940 15092
rect 23884 14702 23886 14754
rect 23938 14702 23940 14754
rect 23884 14690 23940 14702
rect 23884 14532 23940 14542
rect 23772 14420 23828 14430
rect 23772 14326 23828 14364
rect 22988 14242 23044 14252
rect 22876 13804 23156 13860
rect 22316 12964 22372 12974
rect 22316 12870 22372 12908
rect 22540 12852 22596 13804
rect 22652 13636 22708 13646
rect 22652 13542 22708 13580
rect 22876 13636 22932 13646
rect 22764 13524 22820 13534
rect 22764 13430 22820 13468
rect 22764 12964 22820 12974
rect 22876 12964 22932 13580
rect 22820 12908 22932 12964
rect 22764 12870 22820 12908
rect 22988 12852 23044 12862
rect 22540 12796 22708 12852
rect 22204 12180 22260 12190
rect 22204 12086 22260 12124
rect 22204 11956 22260 11966
rect 22204 11618 22260 11900
rect 22652 11788 22708 12796
rect 22988 12758 23044 12796
rect 23100 12516 23156 13804
rect 23884 13524 23940 14476
rect 23100 12450 23156 12460
rect 23436 13074 23492 13086
rect 23436 13022 23438 13074
rect 23490 13022 23492 13074
rect 23436 12740 23492 13022
rect 23884 12962 23940 13468
rect 23884 12910 23886 12962
rect 23938 12910 23940 12962
rect 23884 12898 23940 12910
rect 22764 12180 22820 12190
rect 22820 12124 22932 12180
rect 22764 12114 22820 12124
rect 22428 11676 22708 11788
rect 22204 11566 22206 11618
rect 22258 11566 22260 11618
rect 22204 11554 22260 11566
rect 21868 11302 21924 11340
rect 22092 11330 22148 11340
rect 22428 11506 22484 11518
rect 22428 11454 22430 11506
rect 22482 11454 22484 11506
rect 21756 11106 21812 11116
rect 22092 11172 22148 11182
rect 22092 11078 22148 11116
rect 21868 10500 21924 10510
rect 21868 10498 22372 10500
rect 21868 10446 21870 10498
rect 21922 10446 22372 10498
rect 21868 10444 22372 10446
rect 21868 10434 21924 10444
rect 22316 10050 22372 10444
rect 22316 9998 22318 10050
rect 22370 9998 22372 10050
rect 22316 9986 22372 9998
rect 22428 9938 22484 11454
rect 22428 9886 22430 9938
rect 22482 9886 22484 9938
rect 22428 9874 22484 9886
rect 22540 9716 22596 9726
rect 21084 7474 21588 7476
rect 21084 7422 21086 7474
rect 21138 7422 21588 7474
rect 21084 7420 21588 7422
rect 21756 7586 21812 7598
rect 21756 7534 21758 7586
rect 21810 7534 21812 7586
rect 20748 6802 20916 6804
rect 20748 6750 20750 6802
rect 20802 6750 20916 6802
rect 20748 6748 20916 6750
rect 20748 6738 20804 6748
rect 18620 6638 18622 6690
rect 18674 6638 18676 6690
rect 18620 6626 18676 6638
rect 21084 6692 21140 7420
rect 21084 6626 21140 6636
rect 19628 6580 19684 6590
rect 18396 6132 18452 6142
rect 17948 6130 18452 6132
rect 17948 6078 18398 6130
rect 18450 6078 18452 6130
rect 17948 6076 18452 6078
rect 17836 5908 17892 5918
rect 17948 5908 18004 6076
rect 18396 6066 18452 6076
rect 17836 5906 18004 5908
rect 17836 5854 17838 5906
rect 17890 5854 18004 5906
rect 17836 5852 18004 5854
rect 19628 5908 19684 6524
rect 21756 6580 21812 7534
rect 22092 7476 22148 7486
rect 22092 7382 22148 7420
rect 22540 7362 22596 9660
rect 22652 7700 22708 11676
rect 22764 11282 22820 11294
rect 22764 11230 22766 11282
rect 22818 11230 22820 11282
rect 22764 10836 22820 11230
rect 22876 11282 22932 12124
rect 23212 11508 23268 11518
rect 22876 11230 22878 11282
rect 22930 11230 22932 11282
rect 22876 11218 22932 11230
rect 22988 11396 23044 11406
rect 22988 11282 23044 11340
rect 23212 11394 23268 11452
rect 23212 11342 23214 11394
rect 23266 11342 23268 11394
rect 23212 11330 23268 11342
rect 23436 11396 23492 12684
rect 24444 11956 24500 16046
rect 24668 15316 24724 16268
rect 24668 15250 24724 15260
rect 25228 14420 25284 14430
rect 24780 13748 24836 13758
rect 24780 12068 24836 13692
rect 24780 11974 24836 12012
rect 24892 13074 24948 13086
rect 24892 13022 24894 13074
rect 24946 13022 24948 13074
rect 24444 11890 24500 11900
rect 23436 11330 23492 11340
rect 22988 11230 22990 11282
rect 23042 11230 23044 11282
rect 22988 11218 23044 11230
rect 23660 11284 23716 11294
rect 23660 11190 23716 11228
rect 24108 11284 24164 11294
rect 22764 10780 23156 10836
rect 22652 7634 22708 7644
rect 22876 10612 22932 10622
rect 22540 7310 22542 7362
rect 22594 7310 22596 7362
rect 22540 7298 22596 7310
rect 22876 6692 22932 10556
rect 23100 10500 23156 10780
rect 23100 9938 23156 10444
rect 23996 10500 24052 10510
rect 23996 10406 24052 10444
rect 23100 9886 23102 9938
rect 23154 9886 23156 9938
rect 23100 9874 23156 9886
rect 23996 9940 24052 9950
rect 24108 9940 24164 11228
rect 24556 10612 24612 10622
rect 24556 10518 24612 10556
rect 24892 10164 24948 13022
rect 25228 12962 25284 14364
rect 25340 13858 25396 19964
rect 25452 19794 25508 19806
rect 25452 19742 25454 19794
rect 25506 19742 25508 19794
rect 25452 19236 25508 19742
rect 25452 16548 25508 19180
rect 25788 18452 25844 20188
rect 25900 20018 25956 20300
rect 25900 19966 25902 20018
rect 25954 19966 25956 20018
rect 25900 19954 25956 19966
rect 26012 20300 26180 20356
rect 26012 19796 26068 20300
rect 26124 20132 26180 20142
rect 26124 20018 26180 20076
rect 26124 19966 26126 20018
rect 26178 19966 26180 20018
rect 26124 19954 26180 19966
rect 26236 20020 26292 21532
rect 26348 21522 26404 21532
rect 26572 20916 26628 21868
rect 26348 20860 26628 20916
rect 26348 20802 26404 20860
rect 26348 20750 26350 20802
rect 26402 20750 26404 20802
rect 26348 20738 26404 20750
rect 26348 20020 26404 20030
rect 26236 20018 26404 20020
rect 26236 19966 26350 20018
rect 26402 19966 26404 20018
rect 26236 19964 26404 19966
rect 26348 19954 26404 19964
rect 26012 19740 26404 19796
rect 26348 19458 26404 19740
rect 26348 19406 26350 19458
rect 26402 19406 26404 19458
rect 26348 19394 26404 19406
rect 26460 18562 26516 18574
rect 26460 18510 26462 18562
rect 26514 18510 26516 18562
rect 26124 18452 26180 18462
rect 25788 18450 26180 18452
rect 25788 18398 26126 18450
rect 26178 18398 26180 18450
rect 25788 18396 26180 18398
rect 25564 16882 25620 16894
rect 25564 16830 25566 16882
rect 25618 16830 25620 16882
rect 25564 16772 25620 16830
rect 25564 16706 25620 16716
rect 25452 16492 25620 16548
rect 25564 16098 25620 16492
rect 25564 16046 25566 16098
rect 25618 16046 25620 16098
rect 25564 16034 25620 16046
rect 25452 15986 25508 15998
rect 25452 15934 25454 15986
rect 25506 15934 25508 15986
rect 25452 15876 25508 15934
rect 25788 15876 25844 18396
rect 26124 18386 26180 18396
rect 26460 18340 26516 18510
rect 26460 18274 26516 18284
rect 26572 17892 26628 20860
rect 26684 21698 26740 21710
rect 26684 21646 26686 21698
rect 26738 21646 26740 21698
rect 26684 20580 26740 21646
rect 27020 21586 27076 21598
rect 27020 21534 27022 21586
rect 27074 21534 27076 21586
rect 27020 21476 27076 21534
rect 26796 20804 26852 20814
rect 27020 20804 27076 21420
rect 26852 20748 27076 20804
rect 27244 20804 27300 20814
rect 27356 20804 27412 23436
rect 27580 23378 27636 23390
rect 27580 23326 27582 23378
rect 27634 23326 27636 23378
rect 27244 20802 27412 20804
rect 27244 20750 27246 20802
rect 27298 20750 27412 20802
rect 27244 20748 27412 20750
rect 27468 22930 27524 22942
rect 27468 22878 27470 22930
rect 27522 22878 27524 22930
rect 26796 20710 26852 20748
rect 27244 20738 27300 20748
rect 26684 20524 26964 20580
rect 26908 20244 26964 20524
rect 27468 20578 27524 22878
rect 27580 22148 27636 23326
rect 27692 23154 27748 23996
rect 27692 23102 27694 23154
rect 27746 23102 27748 23154
rect 27692 23090 27748 23102
rect 28588 23154 28644 23166
rect 28588 23102 28590 23154
rect 28642 23102 28644 23154
rect 28476 23044 28532 23054
rect 28476 22950 28532 22988
rect 27692 22932 27748 22942
rect 28252 22932 28308 22942
rect 27692 22482 27748 22876
rect 27692 22430 27694 22482
rect 27746 22430 27748 22482
rect 27692 22418 27748 22430
rect 28140 22930 28308 22932
rect 28140 22878 28254 22930
rect 28306 22878 28308 22930
rect 28140 22876 28308 22878
rect 27580 22092 27860 22148
rect 27692 21812 27748 21822
rect 27692 20802 27748 21756
rect 27804 21698 27860 22092
rect 27804 21646 27806 21698
rect 27858 21646 27860 21698
rect 27804 21634 27860 21646
rect 28028 21252 28084 21262
rect 28028 20916 28084 21196
rect 28140 21140 28196 22876
rect 28252 22866 28308 22876
rect 28588 22372 28644 23102
rect 29932 23156 29988 23166
rect 29260 22372 29316 22382
rect 28588 22316 29260 22372
rect 29260 22278 29316 22316
rect 29932 22370 29988 23100
rect 29932 22318 29934 22370
rect 29986 22318 29988 22370
rect 29932 22306 29988 22318
rect 30044 22372 30100 24670
rect 30044 22278 30100 22316
rect 29372 22258 29428 22270
rect 29372 22206 29374 22258
rect 29426 22206 29428 22258
rect 28252 22148 28308 22158
rect 28252 22054 28308 22092
rect 28140 21074 28196 21084
rect 28700 22036 28756 22046
rect 28028 20860 28196 20916
rect 27692 20750 27694 20802
rect 27746 20750 27748 20802
rect 27692 20738 27748 20750
rect 27580 20692 27636 20702
rect 27580 20598 27636 20636
rect 27468 20526 27470 20578
rect 27522 20526 27524 20578
rect 27468 20514 27524 20526
rect 27916 20580 27972 20590
rect 26908 20130 26964 20188
rect 26908 20078 26910 20130
rect 26962 20078 26964 20130
rect 26908 20066 26964 20078
rect 27020 20132 27076 20142
rect 27020 20038 27076 20076
rect 26684 20020 26740 20030
rect 26684 19908 26740 19964
rect 26684 19852 26908 19908
rect 26852 19796 26908 19852
rect 27468 19796 27524 19806
rect 27804 19796 27860 19806
rect 26852 19740 26964 19796
rect 26796 19346 26852 19358
rect 26796 19294 26798 19346
rect 26850 19294 26852 19346
rect 26684 19236 26740 19246
rect 26796 19236 26852 19294
rect 26740 19180 26852 19236
rect 26908 19236 26964 19740
rect 27468 19794 27860 19796
rect 27468 19742 27470 19794
rect 27522 19742 27806 19794
rect 27858 19742 27860 19794
rect 27468 19740 27860 19742
rect 27020 19236 27076 19246
rect 26908 19234 27076 19236
rect 26908 19182 27022 19234
rect 27074 19182 27076 19234
rect 26908 19180 27076 19182
rect 26684 19170 26740 19180
rect 26908 18452 26964 19180
rect 27020 19170 27076 19180
rect 27244 19234 27300 19246
rect 27244 19182 27246 19234
rect 27298 19182 27300 19234
rect 27244 19012 27300 19182
rect 26796 18396 26964 18452
rect 27132 18788 27188 18798
rect 26796 18340 26852 18396
rect 26796 18274 26852 18284
rect 26628 17836 26852 17892
rect 26572 17798 26628 17836
rect 26796 17780 26852 17836
rect 26796 17724 27076 17780
rect 26796 16884 26852 16894
rect 26796 16790 26852 16828
rect 26684 16100 26740 16110
rect 26684 16006 26740 16044
rect 27020 16098 27076 17724
rect 27020 16046 27022 16098
rect 27074 16046 27076 16098
rect 27020 16034 27076 16046
rect 25452 15820 25844 15876
rect 27132 14532 27188 18732
rect 27244 16548 27300 18956
rect 27468 18676 27524 19740
rect 27804 19730 27860 19740
rect 27692 19012 27748 19022
rect 27692 18918 27748 18956
rect 27468 18610 27524 18620
rect 27468 17444 27524 17454
rect 27468 16994 27524 17388
rect 27468 16942 27470 16994
rect 27522 16942 27524 16994
rect 27468 16930 27524 16942
rect 27244 16482 27300 16492
rect 27244 15988 27300 15998
rect 27244 15894 27300 15932
rect 27804 15988 27860 15998
rect 27356 15876 27412 15886
rect 27356 15782 27412 15820
rect 27132 14466 27188 14476
rect 26012 14308 26068 14318
rect 25340 13806 25342 13858
rect 25394 13806 25396 13858
rect 25340 13794 25396 13806
rect 25900 13858 25956 13870
rect 25900 13806 25902 13858
rect 25954 13806 25956 13858
rect 25788 13746 25844 13758
rect 25788 13694 25790 13746
rect 25842 13694 25844 13746
rect 25228 12910 25230 12962
rect 25282 12910 25284 12962
rect 25228 12898 25284 12910
rect 25452 13522 25508 13534
rect 25452 13470 25454 13522
rect 25506 13470 25508 13522
rect 25340 12852 25396 12862
rect 25340 12290 25396 12796
rect 25340 12238 25342 12290
rect 25394 12238 25396 12290
rect 25340 12226 25396 12238
rect 25452 11844 25508 13470
rect 25564 12964 25620 12974
rect 25564 12290 25620 12908
rect 25564 12238 25566 12290
rect 25618 12238 25620 12290
rect 25564 12226 25620 12238
rect 25676 12850 25732 12862
rect 25676 12798 25678 12850
rect 25730 12798 25732 12850
rect 25676 12180 25732 12798
rect 25788 12402 25844 13694
rect 25788 12350 25790 12402
rect 25842 12350 25844 12402
rect 25788 12338 25844 12350
rect 25788 12180 25844 12190
rect 25676 12178 25844 12180
rect 25676 12126 25790 12178
rect 25842 12126 25844 12178
rect 25676 12124 25844 12126
rect 25788 12114 25844 12124
rect 25452 11778 25508 11788
rect 25788 11396 25844 11406
rect 25788 11302 25844 11340
rect 25228 11172 25284 11182
rect 25900 11172 25956 13806
rect 26012 13748 26068 14252
rect 26124 13972 26180 13982
rect 26124 13970 26516 13972
rect 26124 13918 26126 13970
rect 26178 13918 26516 13970
rect 26124 13916 26516 13918
rect 26124 13906 26180 13916
rect 26348 13748 26404 13758
rect 26012 13746 26404 13748
rect 26012 13694 26350 13746
rect 26402 13694 26404 13746
rect 26012 13692 26404 13694
rect 26012 12962 26068 12974
rect 26012 12910 26014 12962
rect 26066 12910 26068 12962
rect 26012 12852 26068 12910
rect 26236 12964 26292 12974
rect 26236 12870 26292 12908
rect 26012 12786 26068 12796
rect 26236 12516 26292 12526
rect 26012 12404 26068 12414
rect 26012 12178 26068 12348
rect 26236 12290 26292 12460
rect 26236 12238 26238 12290
rect 26290 12238 26292 12290
rect 26236 12226 26292 12238
rect 26012 12126 26014 12178
rect 26066 12126 26068 12178
rect 26012 12114 26068 12126
rect 26348 11956 26404 13692
rect 26460 12292 26516 13916
rect 27132 12962 27188 12974
rect 27132 12910 27134 12962
rect 27186 12910 27188 12962
rect 26796 12740 26852 12750
rect 26572 12292 26628 12302
rect 26460 12290 26628 12292
rect 26460 12238 26574 12290
rect 26626 12238 26628 12290
rect 26460 12236 26628 12238
rect 26572 12226 26628 12236
rect 25228 11170 25956 11172
rect 25228 11118 25230 11170
rect 25282 11118 25956 11170
rect 25228 11116 25956 11118
rect 26236 11900 26404 11956
rect 26796 11956 26852 12684
rect 27132 12516 27188 12910
rect 27692 12962 27748 12974
rect 27692 12910 27694 12962
rect 27746 12910 27748 12962
rect 27132 12450 27188 12460
rect 27468 12850 27524 12862
rect 27468 12798 27470 12850
rect 27522 12798 27524 12850
rect 27468 12180 27524 12798
rect 27692 12404 27748 12910
rect 27804 12628 27860 15932
rect 27916 13636 27972 20524
rect 28140 20244 28196 20860
rect 28252 20692 28308 20702
rect 28252 20598 28308 20636
rect 28028 20130 28084 20142
rect 28028 20078 28030 20130
rect 28082 20078 28084 20130
rect 28028 20020 28084 20078
rect 28028 19012 28084 19964
rect 28140 19906 28196 20188
rect 28588 20020 28644 20030
rect 28588 19926 28644 19964
rect 28140 19854 28142 19906
rect 28194 19854 28196 19906
rect 28140 19842 28196 19854
rect 28028 18946 28084 18956
rect 28588 16098 28644 16110
rect 28588 16046 28590 16098
rect 28642 16046 28644 16098
rect 28028 15876 28084 15886
rect 28028 15782 28084 15820
rect 28588 14308 28644 16046
rect 28700 15148 28756 21980
rect 29372 21812 29428 22206
rect 29708 22148 29764 22158
rect 29372 21746 29428 21756
rect 29484 21924 29540 21934
rect 29484 21588 29540 21868
rect 29372 21532 29540 21588
rect 28700 15092 29092 15148
rect 28700 14308 28756 14318
rect 28588 14306 28700 14308
rect 28588 14254 28590 14306
rect 28642 14254 28700 14306
rect 28588 14252 28700 14254
rect 28588 14242 28644 14252
rect 27916 13570 27972 13580
rect 28140 12964 28196 12974
rect 28140 12870 28196 12908
rect 28476 12964 28532 12974
rect 28476 12850 28532 12908
rect 28476 12798 28478 12850
rect 28530 12798 28532 12850
rect 28476 12786 28532 12798
rect 27804 12562 27860 12572
rect 27748 12348 28308 12404
rect 27692 12310 27748 12348
rect 28140 12180 28196 12190
rect 27468 12114 27524 12124
rect 28028 12178 28196 12180
rect 28028 12126 28142 12178
rect 28194 12126 28196 12178
rect 28028 12124 28196 12126
rect 25228 11106 25284 11116
rect 24892 10098 24948 10108
rect 26012 10164 26068 10174
rect 23996 9938 24164 9940
rect 23996 9886 23998 9938
rect 24050 9886 24164 9938
rect 23996 9884 24164 9886
rect 23996 9874 24052 9884
rect 23548 9826 23604 9838
rect 23548 9774 23550 9826
rect 23602 9774 23604 9826
rect 23548 9716 23604 9774
rect 23548 9650 23604 9660
rect 24668 9044 24724 9054
rect 24668 8950 24724 8988
rect 25340 9044 25396 9054
rect 25340 8950 25396 8988
rect 26012 8260 26068 10108
rect 26124 9044 26180 9054
rect 26236 9044 26292 11900
rect 26796 11890 26852 11900
rect 26908 11956 26964 11966
rect 26460 11396 26516 11406
rect 26348 11172 26404 11182
rect 26348 9940 26404 11116
rect 26460 10612 26516 11340
rect 26684 11394 26740 11406
rect 26684 11342 26686 11394
rect 26738 11342 26740 11394
rect 26572 11284 26628 11294
rect 26572 11190 26628 11228
rect 26572 10612 26628 10622
rect 26460 10610 26628 10612
rect 26460 10558 26574 10610
rect 26626 10558 26628 10610
rect 26460 10556 26628 10558
rect 26572 10546 26628 10556
rect 26684 9940 26740 11342
rect 26348 9938 26628 9940
rect 26348 9886 26350 9938
rect 26402 9886 26628 9938
rect 26348 9884 26628 9886
rect 26348 9874 26404 9884
rect 26572 9826 26628 9884
rect 26684 9874 26740 9884
rect 26572 9774 26574 9826
rect 26626 9774 26628 9826
rect 26572 9762 26628 9774
rect 26180 8988 26292 9044
rect 26796 9602 26852 9614
rect 26796 9550 26798 9602
rect 26850 9550 26852 9602
rect 26124 8978 26180 8988
rect 26236 8260 26292 8270
rect 25788 8258 26292 8260
rect 25788 8206 26238 8258
rect 26290 8206 26292 8258
rect 25788 8204 26292 8206
rect 25564 8148 25620 8158
rect 24444 7924 24500 7934
rect 24220 7586 24276 7598
rect 24220 7534 24222 7586
rect 24274 7534 24276 7586
rect 23772 7476 23828 7486
rect 24220 7476 24276 7534
rect 24444 7586 24500 7868
rect 24444 7534 24446 7586
rect 24498 7534 24500 7586
rect 24444 7522 24500 7534
rect 23772 7474 24276 7476
rect 23772 7422 23774 7474
rect 23826 7422 24276 7474
rect 23772 7420 24276 7422
rect 23772 7410 23828 7420
rect 24108 7252 24164 7262
rect 23884 7250 24164 7252
rect 23884 7198 24110 7250
rect 24162 7198 24164 7250
rect 23884 7196 24164 7198
rect 23884 6916 23940 7196
rect 24108 7186 24164 7196
rect 23548 6860 23940 6916
rect 23548 6802 23604 6860
rect 23548 6750 23550 6802
rect 23602 6750 23604 6802
rect 23548 6738 23604 6750
rect 23884 6692 23940 6702
rect 22932 6636 23044 6692
rect 22876 6598 22932 6636
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 17836 5842 17892 5852
rect 17612 5234 17780 5236
rect 17612 5182 17614 5234
rect 17666 5182 17780 5234
rect 17612 5180 17780 5182
rect 17948 5682 18004 5694
rect 17948 5630 17950 5682
rect 18002 5630 18004 5682
rect 17948 5236 18004 5630
rect 16940 5124 16996 5134
rect 16940 5030 16996 5068
rect 17612 5124 17668 5180
rect 17948 5170 18004 5180
rect 17612 5058 17668 5068
rect 16604 4452 16660 4462
rect 14924 4340 14980 4350
rect 14924 4246 14980 4284
rect 14364 3490 14420 3500
rect 12572 3332 13076 3388
rect 13916 3444 13972 3454
rect 12572 800 12628 3332
rect 13916 800 13972 3388
rect 14812 3444 14868 3454
rect 14812 3330 14868 3388
rect 14812 3278 14814 3330
rect 14866 3278 14868 3330
rect 14812 3266 14868 3278
rect 15260 3444 15316 3454
rect 15260 800 15316 3388
rect 16604 800 16660 4396
rect 17388 4452 17444 4462
rect 17388 4358 17444 4396
rect 18172 4450 18228 4462
rect 18172 4398 18174 4450
rect 18226 4398 18228 4450
rect 16940 3556 16996 3566
rect 16940 3462 16996 3500
rect 18172 3388 18228 4398
rect 19628 4226 19684 5852
rect 21420 5796 21476 5806
rect 21420 5794 21700 5796
rect 21420 5742 21422 5794
rect 21474 5742 21700 5794
rect 21420 5740 21700 5742
rect 21420 5730 21476 5740
rect 21308 5348 21364 5358
rect 21308 5122 21364 5292
rect 21644 5346 21700 5740
rect 21644 5294 21646 5346
rect 21698 5294 21700 5346
rect 21644 5282 21700 5294
rect 21756 5348 21812 6524
rect 22876 6356 22932 6366
rect 22876 6132 22932 6300
rect 22316 6130 22932 6132
rect 22316 6078 22878 6130
rect 22930 6078 22932 6130
rect 22316 6076 22932 6078
rect 21868 5908 21924 5918
rect 21868 5814 21924 5852
rect 22316 5906 22372 6076
rect 22876 6066 22932 6076
rect 22316 5854 22318 5906
rect 22370 5854 22372 5906
rect 22316 5842 22372 5854
rect 21756 5282 21812 5292
rect 22092 5348 22148 5358
rect 22092 5234 22148 5292
rect 22092 5182 22094 5234
rect 22146 5182 22148 5234
rect 22092 5170 22148 5182
rect 21308 5070 21310 5122
rect 21362 5070 21364 5122
rect 21308 5058 21364 5070
rect 21532 4898 21588 4910
rect 21532 4846 21534 4898
rect 21586 4846 21588 4898
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 21532 4564 21588 4846
rect 22988 4564 23044 6636
rect 23884 5124 23940 6636
rect 24220 6580 24276 7420
rect 24276 6524 24724 6580
rect 24220 6514 24276 6524
rect 24668 6130 24724 6524
rect 24668 6078 24670 6130
rect 24722 6078 24724 6130
rect 24668 6020 24724 6078
rect 24668 5954 24724 5964
rect 25340 6020 25396 6030
rect 25340 5926 25396 5964
rect 25564 6018 25620 8092
rect 25676 7588 25732 7598
rect 25676 7494 25732 7532
rect 25676 6804 25732 6814
rect 25788 6804 25844 8204
rect 26236 8194 26292 8204
rect 26572 8034 26628 8046
rect 26572 7982 26574 8034
rect 26626 7982 26628 8034
rect 26572 7812 26628 7982
rect 26572 7746 26628 7756
rect 26348 7700 26404 7710
rect 26124 7588 26180 7598
rect 26124 7474 26180 7532
rect 26124 7422 26126 7474
rect 26178 7422 26180 7474
rect 26124 7410 26180 7422
rect 26348 7474 26404 7644
rect 26348 7422 26350 7474
rect 26402 7422 26404 7474
rect 26348 7410 26404 7422
rect 26572 7476 26628 7486
rect 26796 7476 26852 9550
rect 26572 7474 26852 7476
rect 26572 7422 26574 7474
rect 26626 7422 26852 7474
rect 26572 7420 26852 7422
rect 26908 7476 26964 11900
rect 27468 11844 27524 11854
rect 27244 11508 27300 11518
rect 27020 10612 27076 10622
rect 27020 9826 27076 10556
rect 27020 9774 27022 9826
rect 27074 9774 27076 9826
rect 27020 9762 27076 9774
rect 27244 9714 27300 11452
rect 27468 11396 27524 11788
rect 27468 11394 27748 11396
rect 27468 11342 27470 11394
rect 27522 11342 27748 11394
rect 27468 11340 27748 11342
rect 27468 11330 27524 11340
rect 27356 11282 27412 11294
rect 27356 11230 27358 11282
rect 27410 11230 27412 11282
rect 27356 9828 27412 11230
rect 27692 10610 27748 11340
rect 28028 10722 28084 12124
rect 28140 12114 28196 12124
rect 28252 11618 28308 12348
rect 28588 12180 28644 12190
rect 28588 12086 28644 12124
rect 28252 11566 28254 11618
rect 28306 11566 28308 11618
rect 28252 11554 28308 11566
rect 28028 10670 28030 10722
rect 28082 10670 28084 10722
rect 28028 10658 28084 10670
rect 28364 11282 28420 11294
rect 28364 11230 28366 11282
rect 28418 11230 28420 11282
rect 27692 10558 27694 10610
rect 27746 10558 27748 10610
rect 27692 10546 27748 10558
rect 27916 10612 27972 10622
rect 27356 9762 27412 9772
rect 27580 9940 27636 9950
rect 27580 9826 27636 9884
rect 27580 9774 27582 9826
rect 27634 9774 27636 9826
rect 27244 9662 27246 9714
rect 27298 9662 27300 9714
rect 27244 8372 27300 9662
rect 27244 8306 27300 8316
rect 27020 7476 27076 7486
rect 27468 7476 27524 7486
rect 27580 7476 27636 9774
rect 27916 9714 27972 10556
rect 28364 10612 28420 11230
rect 28588 10612 28644 10622
rect 28364 10610 28644 10612
rect 28364 10558 28590 10610
rect 28642 10558 28644 10610
rect 28364 10556 28644 10558
rect 27916 9662 27918 9714
rect 27970 9662 27972 9714
rect 27916 9650 27972 9662
rect 28140 10498 28196 10510
rect 28140 10446 28142 10498
rect 28194 10446 28196 10498
rect 28140 9716 28196 10446
rect 28364 10164 28420 10556
rect 28588 10546 28644 10556
rect 28140 9650 28196 9660
rect 28252 9828 28308 9838
rect 28252 9492 28308 9772
rect 28252 9426 28308 9436
rect 26908 7474 27412 7476
rect 26908 7422 27022 7474
rect 27074 7422 27412 7474
rect 26908 7420 27412 7422
rect 26572 7410 26628 7420
rect 27020 7410 27076 7420
rect 25676 6802 25844 6804
rect 25676 6750 25678 6802
rect 25730 6750 25844 6802
rect 25676 6748 25844 6750
rect 26012 7250 26068 7262
rect 26012 7198 26014 7250
rect 26066 7198 26068 7250
rect 25676 6738 25732 6748
rect 25564 5966 25566 6018
rect 25618 5966 25620 6018
rect 25564 5954 25620 5966
rect 25228 5684 25284 5694
rect 24780 5682 25284 5684
rect 24780 5630 25230 5682
rect 25282 5630 25284 5682
rect 24780 5628 25284 5630
rect 24668 5236 24724 5246
rect 24780 5236 24836 5628
rect 25228 5618 25284 5628
rect 24668 5234 24836 5236
rect 24668 5182 24670 5234
rect 24722 5182 24836 5234
rect 24668 5180 24836 5182
rect 24668 5170 24724 5180
rect 23884 5030 23940 5068
rect 25452 5124 25508 5134
rect 21532 4508 21812 4564
rect 21756 4450 21812 4508
rect 21756 4398 21758 4450
rect 21810 4398 21812 4450
rect 21756 4386 21812 4398
rect 22540 4562 23044 4564
rect 22540 4510 22990 4562
rect 23042 4510 23044 4562
rect 22540 4508 23044 4510
rect 22540 4338 22596 4508
rect 22988 4498 23044 4508
rect 22540 4286 22542 4338
rect 22594 4286 22596 4338
rect 22540 4274 22596 4286
rect 25452 4338 25508 5068
rect 26012 4452 26068 7198
rect 26124 6466 26180 6478
rect 26124 6414 26126 6466
rect 26178 6414 26180 6466
rect 26124 5124 26180 6414
rect 27356 6244 27412 7420
rect 27468 7474 27636 7476
rect 27468 7422 27470 7474
rect 27522 7422 27636 7474
rect 27468 7420 27636 7422
rect 27468 7410 27524 7420
rect 27580 6692 27636 7420
rect 27916 7476 27972 7486
rect 27916 7382 27972 7420
rect 27580 6626 27636 6636
rect 28140 6690 28196 6702
rect 28140 6638 28142 6690
rect 28194 6638 28196 6690
rect 28140 6468 28196 6638
rect 28364 6578 28420 10108
rect 28588 9716 28644 9726
rect 28588 9622 28644 9660
rect 28700 9492 28756 14252
rect 29036 11620 29092 15092
rect 29260 13076 29316 13086
rect 29372 13076 29428 21532
rect 29596 16772 29652 16782
rect 29596 16678 29652 16716
rect 29708 16436 29764 22092
rect 29820 22146 29876 22158
rect 29820 22094 29822 22146
rect 29874 22094 29876 22146
rect 29820 20244 29876 22094
rect 29932 21812 29988 21822
rect 29932 21474 29988 21756
rect 29932 21422 29934 21474
rect 29986 21422 29988 21474
rect 29932 21410 29988 21422
rect 29820 20178 29876 20188
rect 29932 17108 29988 17118
rect 29932 17014 29988 17052
rect 30044 16996 30100 17006
rect 30044 16902 30100 16940
rect 29708 16380 30100 16436
rect 30044 16322 30100 16380
rect 30044 16270 30046 16322
rect 30098 16270 30100 16322
rect 30044 16258 30100 16270
rect 30156 16212 30212 24892
rect 30268 23044 30324 23054
rect 30268 22482 30324 22988
rect 30268 22430 30270 22482
rect 30322 22430 30324 22482
rect 30268 22418 30324 22430
rect 30380 23042 30436 23054
rect 30380 22990 30382 23042
rect 30434 22990 30436 23042
rect 30380 22820 30436 22990
rect 30492 22932 30548 26852
rect 30492 22866 30548 22876
rect 30380 21924 30436 22764
rect 30492 22596 30548 22606
rect 30492 22502 30548 22540
rect 30380 21858 30436 21868
rect 30492 21476 30548 21486
rect 30380 21420 30492 21476
rect 30380 17108 30436 21420
rect 30492 21382 30548 21420
rect 30492 20580 30548 20590
rect 30492 20486 30548 20524
rect 30492 17108 30548 17118
rect 30380 17106 30548 17108
rect 30380 17054 30494 17106
rect 30546 17054 30548 17106
rect 30380 17052 30548 17054
rect 30380 16884 30436 17052
rect 30492 17042 30548 17052
rect 30380 16818 30436 16828
rect 30156 16146 30212 16156
rect 30492 16100 30548 16110
rect 30268 16098 30548 16100
rect 30268 16046 30494 16098
rect 30546 16046 30548 16098
rect 30268 16044 30548 16046
rect 29932 15986 29988 15998
rect 29932 15934 29934 15986
rect 29986 15934 29988 15986
rect 29484 15876 29540 15886
rect 29484 14418 29540 15820
rect 29932 15876 29988 15934
rect 29932 15810 29988 15820
rect 30044 15876 30100 15886
rect 30044 15874 30212 15876
rect 30044 15822 30046 15874
rect 30098 15822 30212 15874
rect 30044 15820 30212 15822
rect 30044 15810 30100 15820
rect 29708 15484 30100 15540
rect 29596 15428 29652 15438
rect 29708 15428 29764 15484
rect 29596 15426 29764 15428
rect 29596 15374 29598 15426
rect 29650 15374 29764 15426
rect 29596 15372 29764 15374
rect 29596 15362 29652 15372
rect 29820 15314 29876 15326
rect 29820 15262 29822 15314
rect 29874 15262 29876 15314
rect 29820 15148 29876 15262
rect 29596 15092 29876 15148
rect 29932 15316 29988 15326
rect 29596 14644 29652 15092
rect 29596 14550 29652 14588
rect 29932 14532 29988 15260
rect 30044 15148 30100 15484
rect 30156 15428 30212 15820
rect 30156 15362 30212 15372
rect 30268 15316 30324 16044
rect 30492 16034 30548 16044
rect 30604 15876 30660 29260
rect 31164 28754 31220 29484
rect 31276 29204 31332 29934
rect 31388 29652 31444 29662
rect 31500 29652 31556 30158
rect 31388 29650 31556 29652
rect 31388 29598 31390 29650
rect 31442 29598 31556 29650
rect 31388 29596 31556 29598
rect 31388 29586 31444 29596
rect 31612 29426 31668 30380
rect 32172 30370 32228 30380
rect 34076 30882 34132 31612
rect 34076 30830 34078 30882
rect 34130 30830 34132 30882
rect 31948 30098 32004 30110
rect 31948 30046 31950 30098
rect 32002 30046 32004 30098
rect 31948 29540 32004 30046
rect 32508 29988 32564 29998
rect 32508 29894 32564 29932
rect 31948 29474 32004 29484
rect 32956 29764 33012 29774
rect 31612 29374 31614 29426
rect 31666 29374 31668 29426
rect 31612 29362 31668 29374
rect 31276 29138 31332 29148
rect 32508 29204 32564 29214
rect 31164 28702 31166 28754
rect 31218 28702 31220 28754
rect 31164 28690 31220 28702
rect 31388 28812 31780 28868
rect 31388 28644 31444 28812
rect 31612 28644 31668 28654
rect 31276 28642 31444 28644
rect 31276 28590 31390 28642
rect 31442 28590 31444 28642
rect 31276 28588 31444 28590
rect 30828 28532 30884 28542
rect 31276 28532 31332 28588
rect 31388 28578 31444 28588
rect 31500 28642 31668 28644
rect 31500 28590 31614 28642
rect 31666 28590 31668 28642
rect 31500 28588 31668 28590
rect 30828 28530 31332 28532
rect 30828 28478 30830 28530
rect 30882 28478 31332 28530
rect 30828 28476 31332 28478
rect 30828 28466 30884 28476
rect 31500 27524 31556 28588
rect 31612 28578 31668 28588
rect 31164 27468 31556 27524
rect 31164 26908 31220 27468
rect 31724 27188 31780 28812
rect 32508 28866 32564 29148
rect 32508 28814 32510 28866
rect 32562 28814 32564 28866
rect 32508 28802 32564 28814
rect 32844 28642 32900 28654
rect 32844 28590 32846 28642
rect 32898 28590 32900 28642
rect 32620 28420 32676 28430
rect 32620 28326 32676 28364
rect 32844 27972 32900 28590
rect 32844 27906 32900 27916
rect 31836 27748 31892 27758
rect 31836 27746 32004 27748
rect 31836 27694 31838 27746
rect 31890 27694 32004 27746
rect 31836 27692 32004 27694
rect 31836 27682 31892 27692
rect 31836 27188 31892 27198
rect 31388 27186 31892 27188
rect 31388 27134 31838 27186
rect 31890 27134 31892 27186
rect 31388 27132 31892 27134
rect 31164 26852 31332 26908
rect 30716 26290 30772 26302
rect 30716 26238 30718 26290
rect 30770 26238 30772 26290
rect 30716 25844 30772 26238
rect 30716 25778 30772 25788
rect 31164 26290 31220 26302
rect 31164 26238 31166 26290
rect 31218 26238 31220 26290
rect 31164 23604 31220 26238
rect 30716 23548 31220 23604
rect 30716 20244 30772 23548
rect 31276 23492 31332 26852
rect 31388 26178 31444 27132
rect 31836 27122 31892 27132
rect 31500 26964 31556 26974
rect 31948 26964 32004 27692
rect 31500 26962 31948 26964
rect 31500 26910 31502 26962
rect 31554 26910 31948 26962
rect 31500 26908 31948 26910
rect 31500 26898 31556 26908
rect 31388 26126 31390 26178
rect 31442 26126 31444 26178
rect 31388 26114 31444 26126
rect 31948 23940 32004 26908
rect 32956 26908 33012 29708
rect 33404 28756 33460 28766
rect 33404 27858 33460 28700
rect 33964 28420 34020 28430
rect 33628 27972 33684 27982
rect 33628 27878 33684 27916
rect 33404 27806 33406 27858
rect 33458 27806 33460 27858
rect 32956 26852 33236 26908
rect 31948 23846 32004 23884
rect 32172 25172 32228 25182
rect 31500 23828 31556 23838
rect 31276 23426 31332 23436
rect 31388 23714 31444 23726
rect 31388 23662 31390 23714
rect 31442 23662 31444 23714
rect 31052 23268 31108 23278
rect 30828 23042 30884 23054
rect 30828 22990 30830 23042
rect 30882 22990 30884 23042
rect 30828 22372 30884 22990
rect 31052 22596 31108 23212
rect 31276 23266 31332 23278
rect 31276 23214 31278 23266
rect 31330 23214 31332 23266
rect 31164 23156 31220 23166
rect 31164 23062 31220 23100
rect 31052 22530 31108 22540
rect 31276 22372 31332 23214
rect 31388 23156 31444 23662
rect 31500 23378 31556 23772
rect 31500 23326 31502 23378
rect 31554 23326 31556 23378
rect 31500 23314 31556 23326
rect 31612 23156 31668 23166
rect 31388 23154 31668 23156
rect 31388 23102 31614 23154
rect 31666 23102 31668 23154
rect 31388 23100 31668 23102
rect 31612 22932 31668 23100
rect 32060 23154 32116 23166
rect 32060 23102 32062 23154
rect 32114 23102 32116 23154
rect 31612 22866 31668 22876
rect 31836 23042 31892 23054
rect 31836 22990 31838 23042
rect 31890 22990 31892 23042
rect 31836 22372 31892 22990
rect 30828 22316 31332 22372
rect 30940 22146 30996 22158
rect 30940 22094 30942 22146
rect 30994 22094 30996 22146
rect 30940 22036 30996 22094
rect 30940 21970 30996 21980
rect 31164 21586 31220 21598
rect 31164 21534 31166 21586
rect 31218 21534 31220 21586
rect 31164 20580 31220 21534
rect 31164 20514 31220 20524
rect 30716 20178 30772 20188
rect 31276 19684 31332 22316
rect 31612 22316 31892 22372
rect 31500 22146 31556 22158
rect 31500 22094 31502 22146
rect 31554 22094 31556 22146
rect 31388 22036 31444 22046
rect 31388 21474 31444 21980
rect 31500 21924 31556 22094
rect 31500 21858 31556 21868
rect 31612 21700 31668 22316
rect 31948 22260 32004 22270
rect 31948 22166 32004 22204
rect 31724 22146 31780 22158
rect 31724 22094 31726 22146
rect 31778 22094 31780 22146
rect 31724 22036 31780 22094
rect 31836 22148 31892 22158
rect 31836 22054 31892 22092
rect 31724 21970 31780 21980
rect 32060 22036 32116 23102
rect 32172 22370 32228 25116
rect 32284 23940 32340 23950
rect 32284 23846 32340 23884
rect 32844 23940 32900 23950
rect 32284 23154 32340 23166
rect 32284 23102 32286 23154
rect 32338 23102 32340 23154
rect 32284 23044 32340 23102
rect 32284 22978 32340 22988
rect 32844 22372 32900 23884
rect 33068 23828 33124 23838
rect 33068 23734 33124 23772
rect 32172 22318 32174 22370
rect 32226 22318 32228 22370
rect 32172 22306 32228 22318
rect 32620 22370 32900 22372
rect 32620 22318 32846 22370
rect 32898 22318 32900 22370
rect 32620 22316 32900 22318
rect 32508 22258 32564 22270
rect 32508 22206 32510 22258
rect 32562 22206 32564 22258
rect 32396 22148 32452 22158
rect 32060 21970 32116 21980
rect 32284 22146 32452 22148
rect 32284 22094 32398 22146
rect 32450 22094 32452 22146
rect 32284 22092 32452 22094
rect 31836 21924 31892 21934
rect 31724 21700 31780 21710
rect 31612 21644 31724 21700
rect 31724 21634 31780 21644
rect 31836 21698 31892 21868
rect 31836 21646 31838 21698
rect 31890 21646 31892 21698
rect 31836 21634 31892 21646
rect 31388 21422 31390 21474
rect 31442 21422 31444 21474
rect 31388 21410 31444 21422
rect 31836 21364 31892 21374
rect 31836 20914 31892 21308
rect 31836 20862 31838 20914
rect 31890 20862 31892 20914
rect 31836 20850 31892 20862
rect 32284 20914 32340 22092
rect 32396 22082 32452 22092
rect 32508 21924 32564 22206
rect 32508 21858 32564 21868
rect 32620 21810 32676 22316
rect 32844 22306 32900 22316
rect 33180 22148 33236 26852
rect 32620 21758 32622 21810
rect 32674 21758 32676 21810
rect 32620 21746 32676 21758
rect 32956 22092 33236 22148
rect 32284 20862 32286 20914
rect 32338 20862 32340 20914
rect 32284 20850 32340 20862
rect 32508 21588 32564 21598
rect 31164 19460 31220 19470
rect 31164 19366 31220 19404
rect 31276 17890 31332 19628
rect 31612 20802 31668 20814
rect 31612 20750 31614 20802
rect 31666 20750 31668 20802
rect 31500 19460 31556 19470
rect 31500 19366 31556 19404
rect 31612 18788 31668 20750
rect 31612 18722 31668 18732
rect 31724 19234 31780 19246
rect 31724 19182 31726 19234
rect 31778 19182 31780 19234
rect 31724 18564 31780 19182
rect 32060 19236 32116 19246
rect 31948 18676 32004 18686
rect 32060 18676 32116 19180
rect 31948 18674 32116 18676
rect 31948 18622 31950 18674
rect 32002 18622 32116 18674
rect 31948 18620 32116 18622
rect 32172 19234 32228 19246
rect 32172 19182 32174 19234
rect 32226 19182 32228 19234
rect 31948 18610 32004 18620
rect 31276 17838 31278 17890
rect 31330 17838 31332 17890
rect 31276 17826 31332 17838
rect 31500 18562 31780 18564
rect 31500 18510 31726 18562
rect 31778 18510 31780 18562
rect 31500 18508 31780 18510
rect 30268 15250 30324 15260
rect 30380 15820 30660 15876
rect 30716 17108 30772 17118
rect 30044 15092 30212 15148
rect 29820 14530 29988 14532
rect 29820 14478 29934 14530
rect 29986 14478 29988 14530
rect 29820 14476 29988 14478
rect 29484 14366 29486 14418
rect 29538 14366 29540 14418
rect 29484 14354 29540 14366
rect 29708 14420 29764 14430
rect 29708 14326 29764 14364
rect 29260 13074 29540 13076
rect 29260 13022 29262 13074
rect 29314 13022 29540 13074
rect 29260 13020 29540 13022
rect 29260 13010 29316 13020
rect 29484 12962 29540 13020
rect 29484 12910 29486 12962
rect 29538 12910 29540 12962
rect 29484 12898 29540 12910
rect 29372 12852 29428 12862
rect 29148 12292 29204 12302
rect 29148 12198 29204 12236
rect 28924 11564 29316 11620
rect 28924 9940 28980 11564
rect 29260 11506 29316 11564
rect 29260 11454 29262 11506
rect 29314 11454 29316 11506
rect 29260 11442 29316 11454
rect 29260 10836 29316 10846
rect 29372 10836 29428 12796
rect 29708 11172 29764 11182
rect 29820 11172 29876 14476
rect 29932 14466 29988 14476
rect 29932 12964 29988 12974
rect 29932 12870 29988 12908
rect 30044 12852 30100 12862
rect 30044 12758 30100 12796
rect 30156 12738 30212 15092
rect 30380 14308 30436 15820
rect 30492 15540 30548 15550
rect 30492 14642 30548 15484
rect 30604 15540 30660 15550
rect 30716 15540 30772 17052
rect 30940 16996 30996 17006
rect 30940 16902 30996 16940
rect 31164 16884 31220 16894
rect 31164 16100 31220 16828
rect 31388 16882 31444 16894
rect 31388 16830 31390 16882
rect 31442 16830 31444 16882
rect 31388 16772 31444 16830
rect 31388 16212 31444 16716
rect 31388 16146 31444 16156
rect 30604 15538 30772 15540
rect 30604 15486 30606 15538
rect 30658 15486 30772 15538
rect 30604 15484 30772 15486
rect 30604 15474 30660 15484
rect 30716 15148 30772 15484
rect 31052 15874 31108 15886
rect 31052 15822 31054 15874
rect 31106 15822 31108 15874
rect 31052 15428 31108 15822
rect 31164 15540 31220 16044
rect 31276 15540 31332 15550
rect 31164 15538 31332 15540
rect 31164 15486 31278 15538
rect 31330 15486 31332 15538
rect 31164 15484 31332 15486
rect 31052 15362 31108 15372
rect 30716 15092 31220 15148
rect 30492 14590 30494 14642
rect 30546 14590 30548 14642
rect 30492 14578 30548 14590
rect 30940 14644 30996 14654
rect 30940 14550 30996 14588
rect 30604 14420 30660 14430
rect 30604 14326 30660 14364
rect 31164 14418 31220 15092
rect 31164 14366 31166 14418
rect 31218 14366 31220 14418
rect 31164 14354 31220 14366
rect 30380 14214 30436 14252
rect 31052 14308 31108 14318
rect 31052 14214 31108 14252
rect 31276 13858 31332 15484
rect 31276 13806 31278 13858
rect 31330 13806 31332 13858
rect 31276 13794 31332 13806
rect 31388 15540 31444 15550
rect 30940 12964 30996 12974
rect 30940 12870 30996 12908
rect 31388 12962 31444 15484
rect 31388 12910 31390 12962
rect 31442 12910 31444 12962
rect 31388 12898 31444 12910
rect 30716 12852 30772 12862
rect 30716 12758 30772 12796
rect 30156 12686 30158 12738
rect 30210 12686 30212 12738
rect 30156 11508 30212 12686
rect 31164 12740 31220 12750
rect 31164 12738 31444 12740
rect 31164 12686 31166 12738
rect 31218 12686 31444 12738
rect 31164 12684 31444 12686
rect 31164 12674 31220 12684
rect 30828 12628 30884 12638
rect 30268 12404 30324 12414
rect 30268 12310 30324 12348
rect 30156 11442 30212 11452
rect 29764 11116 29876 11172
rect 29708 11106 29764 11116
rect 29260 10834 30212 10836
rect 29260 10782 29262 10834
rect 29314 10782 30212 10834
rect 29260 10780 30212 10782
rect 29260 10770 29316 10780
rect 30156 10722 30212 10780
rect 30156 10670 30158 10722
rect 30210 10670 30212 10722
rect 30156 10658 30212 10670
rect 29036 10612 29092 10622
rect 29036 10518 29092 10556
rect 29596 10610 29652 10622
rect 29596 10558 29598 10610
rect 29650 10558 29652 10610
rect 29148 10498 29204 10510
rect 29148 10446 29150 10498
rect 29202 10446 29204 10498
rect 29148 10052 29204 10446
rect 29148 9986 29204 9996
rect 29596 10164 29652 10558
rect 29820 10612 29876 10622
rect 29820 10518 29876 10556
rect 30044 10500 30100 10510
rect 30044 10498 30212 10500
rect 30044 10446 30046 10498
rect 30098 10446 30212 10498
rect 30044 10444 30212 10446
rect 30044 10434 30100 10444
rect 29484 9940 29540 9950
rect 28924 9884 29092 9940
rect 29036 9828 29092 9884
rect 29260 9938 29540 9940
rect 29260 9886 29486 9938
rect 29538 9886 29540 9938
rect 29260 9884 29540 9886
rect 29148 9828 29204 9838
rect 29036 9772 29148 9828
rect 29148 9734 29204 9772
rect 28588 9436 28756 9492
rect 28588 8428 28644 9436
rect 28364 6526 28366 6578
rect 28418 6526 28420 6578
rect 28364 6514 28420 6526
rect 28476 8372 28644 8428
rect 28700 9154 28756 9166
rect 28700 9102 28702 9154
rect 28754 9102 28756 9154
rect 28476 7588 28532 8372
rect 28588 7700 28644 7710
rect 28588 7606 28644 7644
rect 28476 7474 28532 7532
rect 28476 7422 28478 7474
rect 28530 7422 28532 7474
rect 28140 6402 28196 6412
rect 28364 6356 28420 6366
rect 28476 6356 28532 7422
rect 28588 7364 28644 7374
rect 28588 7270 28644 7308
rect 28420 6300 28532 6356
rect 28364 6290 28420 6300
rect 27356 6188 28308 6244
rect 28252 6130 28308 6188
rect 28252 6078 28254 6130
rect 28306 6078 28308 6130
rect 28252 6066 28308 6078
rect 28588 5906 28644 5918
rect 28588 5854 28590 5906
rect 28642 5854 28644 5906
rect 28588 5460 28644 5854
rect 28588 5394 28644 5404
rect 26796 5236 26852 5246
rect 26796 5142 26852 5180
rect 27244 5236 27300 5246
rect 27244 5142 27300 5180
rect 28588 5236 28644 5246
rect 28700 5236 28756 9102
rect 29260 8148 29316 9884
rect 29484 9874 29540 9884
rect 29596 9826 29652 10108
rect 29932 10388 29988 10398
rect 29596 9774 29598 9826
rect 29650 9774 29652 9826
rect 29596 9762 29652 9774
rect 29820 9826 29876 9838
rect 29820 9774 29822 9826
rect 29874 9774 29876 9826
rect 29372 9604 29428 9614
rect 29372 9602 29652 9604
rect 29372 9550 29374 9602
rect 29426 9550 29652 9602
rect 29372 9548 29652 9550
rect 29372 9538 29428 9548
rect 29484 8820 29540 8830
rect 29484 8258 29540 8764
rect 29596 8370 29652 9548
rect 29820 9380 29876 9774
rect 29820 9314 29876 9324
rect 29932 8428 29988 10332
rect 30156 9828 30212 10444
rect 30492 10052 30548 10062
rect 30492 9958 30548 9996
rect 30716 9828 30772 9838
rect 30156 9772 30324 9828
rect 30156 9602 30212 9614
rect 30156 9550 30158 9602
rect 30210 9550 30212 9602
rect 30156 8820 30212 9550
rect 30156 8754 30212 8764
rect 30268 8484 30324 9772
rect 29596 8318 29598 8370
rect 29650 8318 29652 8370
rect 29596 8306 29652 8318
rect 29820 8372 29988 8428
rect 30156 8428 30324 8484
rect 30604 9826 30772 9828
rect 30604 9774 30718 9826
rect 30770 9774 30772 9826
rect 30604 9772 30772 9774
rect 29484 8206 29486 8258
rect 29538 8206 29540 8258
rect 29484 8194 29540 8206
rect 29708 8148 29764 8158
rect 29820 8148 29876 8372
rect 30156 8370 30212 8428
rect 30156 8318 30158 8370
rect 30210 8318 30212 8370
rect 30156 8306 30212 8318
rect 30492 8372 30548 8382
rect 29932 8260 29988 8270
rect 29932 8166 29988 8204
rect 30492 8258 30548 8316
rect 30492 8206 30494 8258
rect 30546 8206 30548 8258
rect 30492 8194 30548 8206
rect 29260 8082 29316 8092
rect 29596 8146 29876 8148
rect 29596 8094 29710 8146
rect 29762 8094 29876 8146
rect 29596 8092 29876 8094
rect 29596 7924 29652 8092
rect 29708 8082 29764 8092
rect 29036 7868 29652 7924
rect 29036 7586 29092 7868
rect 29596 7700 29652 7710
rect 29596 7606 29652 7644
rect 29036 7534 29038 7586
rect 29090 7534 29092 7586
rect 29036 7522 29092 7534
rect 30156 7588 30212 7598
rect 30156 7494 30212 7532
rect 28812 7476 28868 7486
rect 28812 7382 28868 7420
rect 29372 7476 29428 7486
rect 29372 7382 29428 7420
rect 29820 7476 29876 7486
rect 29596 7364 29652 7374
rect 29596 7270 29652 7308
rect 29708 6916 29764 6926
rect 29708 6822 29764 6860
rect 29372 6692 29428 6702
rect 29260 6636 29372 6692
rect 29148 6578 29204 6590
rect 29148 6526 29150 6578
rect 29202 6526 29204 6578
rect 28644 5180 28756 5236
rect 28588 5142 28644 5180
rect 26124 5058 26180 5068
rect 26236 4452 26292 4462
rect 26012 4450 26292 4452
rect 26012 4398 26238 4450
rect 26290 4398 26292 4450
rect 26012 4396 26292 4398
rect 26236 4386 26292 4396
rect 25452 4286 25454 4338
rect 25506 4286 25508 4338
rect 25452 4274 25508 4286
rect 28364 4340 28420 4350
rect 19628 4174 19630 4226
rect 19682 4174 19684 4226
rect 19628 4162 19684 4174
rect 28364 4226 28420 4284
rect 28364 4174 28366 4226
rect 28418 4174 28420 4226
rect 28364 4162 28420 4174
rect 28700 3666 28756 5180
rect 28812 6468 28868 6478
rect 28812 5348 28868 6412
rect 28812 4338 28868 5292
rect 28812 4286 28814 4338
rect 28866 4286 28868 4338
rect 28812 4274 28868 4286
rect 29036 5906 29092 5918
rect 29036 5854 29038 5906
rect 29090 5854 29092 5906
rect 29036 4340 29092 5854
rect 29148 5460 29204 6526
rect 29260 6130 29316 6636
rect 29372 6598 29428 6636
rect 29596 6468 29652 6478
rect 29596 6374 29652 6412
rect 29260 6078 29262 6130
rect 29314 6078 29316 6130
rect 29260 6066 29316 6078
rect 29260 5460 29316 5470
rect 29148 5404 29260 5460
rect 29036 4246 29092 4284
rect 29260 5234 29316 5404
rect 29260 5182 29262 5234
rect 29314 5182 29316 5234
rect 29260 4338 29316 5182
rect 29708 4564 29764 4574
rect 29820 4564 29876 7420
rect 30604 7476 30660 9772
rect 30716 9762 30772 9772
rect 30828 9268 30884 12572
rect 31276 9828 31332 9838
rect 31276 9604 31332 9772
rect 31276 9538 31332 9548
rect 30828 9202 30884 9212
rect 31164 9156 31220 9166
rect 31052 9154 31220 9156
rect 31052 9102 31166 9154
rect 31218 9102 31220 9154
rect 31052 9100 31220 9102
rect 31052 8596 31108 9100
rect 31164 9090 31220 9100
rect 31276 9042 31332 9054
rect 31276 8990 31278 9042
rect 31330 8990 31332 9042
rect 31052 8530 31108 8540
rect 31164 8818 31220 8830
rect 31164 8766 31166 8818
rect 31218 8766 31220 8818
rect 30716 8034 30772 8046
rect 30716 7982 30718 8034
rect 30770 7982 30772 8034
rect 30716 7588 30772 7982
rect 30828 8036 30884 8046
rect 30828 7942 30884 7980
rect 30940 8034 30996 8046
rect 30940 7982 30942 8034
rect 30994 7982 30996 8034
rect 30940 7812 30996 7982
rect 31052 8036 31108 8046
rect 31052 7942 31108 7980
rect 30940 7746 30996 7756
rect 30828 7588 30884 7598
rect 30716 7586 30884 7588
rect 30716 7534 30830 7586
rect 30882 7534 30884 7586
rect 30716 7532 30884 7534
rect 30828 7522 30884 7532
rect 30604 7410 30660 7420
rect 31164 7362 31220 8766
rect 31276 7700 31332 8990
rect 31276 7634 31332 7644
rect 31164 7310 31166 7362
rect 31218 7310 31220 7362
rect 31164 7298 31220 7310
rect 31388 5234 31444 12684
rect 31500 12404 31556 18508
rect 31724 18498 31780 18508
rect 31612 18228 31668 18238
rect 31612 18134 31668 18172
rect 31612 17890 31668 17902
rect 31612 17838 31614 17890
rect 31666 17838 31668 17890
rect 31612 17444 31668 17838
rect 32172 17668 32228 19182
rect 32508 19234 32564 21532
rect 32508 19182 32510 19234
rect 32562 19182 32564 19234
rect 32508 19170 32564 19182
rect 32284 18452 32340 18462
rect 32284 18358 32340 18396
rect 32956 18004 33012 22092
rect 33180 21700 33236 21710
rect 33180 21606 33236 21644
rect 33068 20916 33124 20926
rect 33404 20916 33460 27806
rect 33964 27186 34020 28364
rect 33964 27134 33966 27186
rect 34018 27134 34020 27186
rect 33964 27122 34020 27134
rect 34076 25508 34132 30830
rect 34188 29652 34244 32286
rect 34300 31444 34356 34972
rect 34412 35026 34468 35038
rect 34412 34974 34414 35026
rect 34466 34974 34468 35026
rect 34412 34018 34468 34974
rect 34748 34916 34804 34926
rect 34748 34822 34804 34860
rect 34412 33966 34414 34018
rect 34466 33966 34468 34018
rect 34412 32564 34468 33966
rect 34860 33346 34916 33358
rect 34860 33294 34862 33346
rect 34914 33294 34916 33346
rect 34524 32564 34580 32574
rect 34412 32562 34580 32564
rect 34412 32510 34526 32562
rect 34578 32510 34580 32562
rect 34412 32508 34580 32510
rect 34412 31778 34468 32508
rect 34524 32498 34580 32508
rect 34860 32564 34916 33294
rect 34860 32498 34916 32508
rect 35084 32674 35140 35756
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35756 35028 35812 35038
rect 35756 35026 36596 35028
rect 35756 34974 35758 35026
rect 35810 34974 36596 35026
rect 35756 34972 36596 34974
rect 35756 34962 35812 34972
rect 35420 34804 35476 34814
rect 35420 34802 35588 34804
rect 35420 34750 35422 34802
rect 35474 34750 35588 34802
rect 35420 34748 35588 34750
rect 35420 34738 35476 34748
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35532 33572 35588 34748
rect 35644 34692 35700 34702
rect 35644 34690 35924 34692
rect 35644 34638 35646 34690
rect 35698 34638 35924 34690
rect 35644 34636 35924 34638
rect 35644 34626 35700 34636
rect 35084 32622 35086 32674
rect 35138 32622 35140 32674
rect 34748 32452 34804 32462
rect 34748 32358 34804 32396
rect 34412 31726 34414 31778
rect 34466 31726 34468 31778
rect 34412 31714 34468 31726
rect 34748 31780 34804 31790
rect 34748 31666 34804 31724
rect 35084 31778 35140 32622
rect 35196 33516 35588 33572
rect 35196 32564 35252 33516
rect 35308 33348 35364 33358
rect 35308 33254 35364 33292
rect 35756 33234 35812 33246
rect 35756 33182 35758 33234
rect 35810 33182 35812 33234
rect 35756 32900 35812 33182
rect 35308 32844 35812 32900
rect 35308 32786 35364 32844
rect 35308 32734 35310 32786
rect 35362 32734 35364 32786
rect 35308 32722 35364 32734
rect 35420 32564 35476 32574
rect 35196 32562 35476 32564
rect 35196 32510 35422 32562
rect 35474 32510 35476 32562
rect 35196 32508 35476 32510
rect 35420 32498 35476 32508
rect 35532 32564 35588 32574
rect 35532 32562 35700 32564
rect 35532 32510 35534 32562
rect 35586 32510 35700 32562
rect 35532 32508 35700 32510
rect 35532 32498 35588 32508
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35532 31892 35588 31902
rect 35532 31798 35588 31836
rect 35084 31726 35086 31778
rect 35138 31726 35140 31778
rect 35084 31714 35140 31726
rect 35644 31780 35700 32508
rect 35644 31714 35700 31724
rect 35756 32562 35812 32574
rect 35756 32510 35758 32562
rect 35810 32510 35812 32562
rect 34748 31614 34750 31666
rect 34802 31614 34804 31666
rect 34748 31602 34804 31614
rect 35532 31668 35588 31678
rect 35532 31574 35588 31612
rect 35308 31556 35364 31566
rect 35644 31556 35700 31566
rect 35756 31556 35812 32510
rect 35868 32116 35924 34636
rect 36540 34242 36596 34972
rect 36540 34190 36542 34242
rect 36594 34190 36596 34242
rect 36540 34178 36596 34190
rect 37548 34916 37604 34926
rect 37212 34130 37268 34142
rect 37212 34078 37214 34130
rect 37266 34078 37268 34130
rect 36316 33572 36372 33582
rect 36316 32788 36372 33516
rect 37212 33572 37268 34078
rect 37212 33506 37268 33516
rect 37212 33348 37268 33358
rect 36316 32786 36708 32788
rect 36316 32734 36318 32786
rect 36370 32734 36708 32786
rect 36316 32732 36708 32734
rect 36316 32722 36372 32732
rect 36652 32562 36708 32732
rect 36652 32510 36654 32562
rect 36706 32510 36708 32562
rect 36652 32498 36708 32510
rect 35868 32050 35924 32060
rect 37100 32452 37156 32462
rect 36988 31892 37044 31902
rect 36988 31798 37044 31836
rect 35308 31554 35476 31556
rect 35308 31502 35310 31554
rect 35362 31502 35476 31554
rect 35308 31500 35476 31502
rect 35308 31490 35364 31500
rect 34300 31388 34692 31444
rect 34300 31220 34356 31230
rect 34300 31106 34356 31164
rect 34300 31054 34302 31106
rect 34354 31054 34356 31106
rect 34300 31042 34356 31054
rect 34188 29586 34244 29596
rect 34636 26516 34692 31388
rect 35420 31332 35476 31500
rect 35700 31500 35812 31556
rect 36540 31668 36596 31678
rect 35644 31462 35700 31500
rect 35420 31276 35924 31332
rect 35868 31218 35924 31276
rect 35868 31166 35870 31218
rect 35922 31166 35924 31218
rect 35868 31154 35924 31166
rect 35756 30994 35812 31006
rect 35756 30942 35758 30994
rect 35810 30942 35812 30994
rect 35084 30884 35140 30894
rect 35084 27188 35140 30828
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35756 29652 35812 30942
rect 35868 30996 35924 31006
rect 35868 30210 35924 30940
rect 36540 30994 36596 31612
rect 36540 30942 36542 30994
rect 36594 30942 36596 30994
rect 36540 30930 36596 30942
rect 36988 30996 37044 31006
rect 37100 30996 37156 32396
rect 37212 31780 37268 33292
rect 37436 32450 37492 32462
rect 37436 32398 37438 32450
rect 37490 32398 37492 32450
rect 37324 32004 37380 32014
rect 37436 32004 37492 32398
rect 37324 32002 37492 32004
rect 37324 31950 37326 32002
rect 37378 31950 37492 32002
rect 37324 31948 37492 31950
rect 37324 31938 37380 31948
rect 37212 31724 37380 31780
rect 36988 30994 37156 30996
rect 36988 30942 36990 30994
rect 37042 30942 37156 30994
rect 36988 30940 37156 30942
rect 37212 31556 37268 31566
rect 35868 30158 35870 30210
rect 35922 30158 35924 30210
rect 35868 30146 35924 30158
rect 36316 30322 36372 30334
rect 36316 30270 36318 30322
rect 36370 30270 36372 30322
rect 36316 30212 36372 30270
rect 36988 30324 37044 30940
rect 36988 30258 37044 30268
rect 36876 30212 36932 30222
rect 37212 30212 37268 31500
rect 37324 30322 37380 31724
rect 37548 30994 37604 34860
rect 39564 32452 39620 32462
rect 39564 32358 39620 32396
rect 37548 30942 37550 30994
rect 37602 30942 37604 30994
rect 37548 30436 37604 30942
rect 37772 31106 37828 31118
rect 37772 31054 37774 31106
rect 37826 31054 37828 31106
rect 37772 30996 37828 31054
rect 37772 30930 37828 30940
rect 39228 30996 39284 31006
rect 37548 30380 37828 30436
rect 37324 30270 37326 30322
rect 37378 30270 37380 30322
rect 37324 30258 37380 30270
rect 36316 30210 36932 30212
rect 36316 30158 36878 30210
rect 36930 30158 36932 30210
rect 36316 30156 36932 30158
rect 36876 30146 36932 30156
rect 37100 30156 37268 30212
rect 37548 30210 37604 30222
rect 37548 30158 37550 30210
rect 37602 30158 37604 30210
rect 36988 30100 37044 30110
rect 35756 29586 35812 29596
rect 36204 29986 36260 29998
rect 36204 29934 36206 29986
rect 36258 29934 36260 29986
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35532 27746 35588 27758
rect 35532 27694 35534 27746
rect 35586 27694 35588 27746
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 27188 35252 27198
rect 35084 27132 35196 27188
rect 35196 27094 35252 27132
rect 34748 27074 34804 27086
rect 34748 27022 34750 27074
rect 34802 27022 34804 27074
rect 34748 26964 34804 27022
rect 34748 26898 34804 26908
rect 35532 26852 35588 27694
rect 35980 27300 36036 27310
rect 36204 27300 36260 29934
rect 36428 29988 36484 29998
rect 36428 29540 36484 29932
rect 36428 29474 36484 29484
rect 36764 29764 36820 29774
rect 36764 29426 36820 29708
rect 36876 29652 36932 29662
rect 36876 29558 36932 29596
rect 36988 29650 37044 30044
rect 36988 29598 36990 29650
rect 37042 29598 37044 29650
rect 36988 29586 37044 29598
rect 36764 29374 36766 29426
rect 36818 29374 36820 29426
rect 36764 28644 36820 29374
rect 36764 28588 37044 28644
rect 36036 27244 36260 27300
rect 36316 28532 36372 28542
rect 35756 27188 35812 27198
rect 35308 26796 35532 26852
rect 34972 26516 35028 26526
rect 34692 26514 35028 26516
rect 34692 26462 34974 26514
rect 35026 26462 35028 26514
rect 34692 26460 35028 26462
rect 34636 26422 34692 26460
rect 34972 26450 35028 26460
rect 35308 26514 35364 26796
rect 35532 26786 35588 26796
rect 35644 27132 35756 27188
rect 35812 27132 35924 27188
rect 35308 26462 35310 26514
rect 35362 26462 35364 26514
rect 35308 26450 35364 26462
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34076 25442 34132 25452
rect 35644 24836 35700 27132
rect 35756 27122 35812 27132
rect 35868 27074 35924 27132
rect 35868 27022 35870 27074
rect 35922 27022 35924 27074
rect 35868 27010 35924 27022
rect 35980 27074 36036 27244
rect 35980 27022 35982 27074
rect 36034 27022 36036 27074
rect 35980 27010 36036 27022
rect 36092 27076 36148 27086
rect 36092 26982 36148 27020
rect 35756 26964 35812 26974
rect 35756 26516 35812 26908
rect 36204 26964 36260 26974
rect 36204 26870 36260 26908
rect 36316 26740 36372 28476
rect 36988 27188 37044 28588
rect 37100 27972 37156 30156
rect 37324 30100 37380 30110
rect 37100 27906 37156 27916
rect 37212 30044 37324 30100
rect 37212 27972 37268 30044
rect 37324 30034 37380 30044
rect 37436 29988 37492 29998
rect 37436 29426 37492 29932
rect 37436 29374 37438 29426
rect 37490 29374 37492 29426
rect 37436 29362 37492 29374
rect 37548 29316 37604 30158
rect 37660 30210 37716 30222
rect 37660 30158 37662 30210
rect 37714 30158 37716 30210
rect 37660 29764 37716 30158
rect 37660 29698 37716 29708
rect 37772 29538 37828 30380
rect 38668 30100 38724 30110
rect 38668 30006 38724 30044
rect 39228 30098 39284 30940
rect 39228 30046 39230 30098
rect 39282 30046 39284 30098
rect 39228 30034 39284 30046
rect 39340 30098 39396 30110
rect 39340 30046 39342 30098
rect 39394 30046 39396 30098
rect 39004 29988 39060 29998
rect 39004 29894 39060 29932
rect 37772 29486 37774 29538
rect 37826 29486 37828 29538
rect 37660 29316 37716 29326
rect 37548 29314 37716 29316
rect 37548 29262 37662 29314
rect 37714 29262 37716 29314
rect 37548 29260 37716 29262
rect 37660 29250 37716 29260
rect 37660 28532 37716 28542
rect 37772 28532 37828 29486
rect 37996 29540 38052 29550
rect 37996 29446 38052 29484
rect 37716 28476 37828 28532
rect 37660 28466 37716 28476
rect 39340 28196 39396 30046
rect 39116 28140 39396 28196
rect 38556 27972 38612 27982
rect 37212 27970 37492 27972
rect 37212 27918 37214 27970
rect 37266 27918 37492 27970
rect 37212 27916 37492 27918
rect 37212 27906 37268 27916
rect 37324 27188 37380 27198
rect 36988 27186 37380 27188
rect 36988 27134 37326 27186
rect 37378 27134 37380 27186
rect 36988 27132 37380 27134
rect 36428 26962 36484 26974
rect 36428 26910 36430 26962
rect 36482 26910 36484 26962
rect 36428 26908 36484 26910
rect 36988 26964 37044 26974
rect 36428 26852 36932 26908
rect 36988 26870 37044 26908
rect 36428 26786 36484 26796
rect 36204 26684 36372 26740
rect 35868 26516 35924 26526
rect 35756 26514 35924 26516
rect 35756 26462 35870 26514
rect 35922 26462 35924 26514
rect 35756 26460 35924 26462
rect 35868 26292 35924 26460
rect 35868 26226 35924 26236
rect 36204 26290 36260 26684
rect 36204 26238 36206 26290
rect 36258 26238 36260 26290
rect 36204 26226 36260 26238
rect 36316 26290 36372 26302
rect 36316 26238 36318 26290
rect 36370 26238 36372 26290
rect 35644 24770 35700 24780
rect 36092 24724 36148 24734
rect 36316 24724 36372 26238
rect 36764 26292 36820 26302
rect 36764 26198 36820 26236
rect 36148 24668 36372 24724
rect 36428 24836 36484 24846
rect 35868 24610 35924 24622
rect 35868 24558 35870 24610
rect 35922 24558 35924 24610
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 24052 35252 24062
rect 35196 23958 35252 23996
rect 35868 23940 35924 24558
rect 35980 24164 36036 24174
rect 35980 24050 36036 24108
rect 35980 23998 35982 24050
rect 36034 23998 36036 24050
rect 35980 23986 36036 23998
rect 36092 24052 36148 24668
rect 36092 23986 36148 23996
rect 36428 24050 36484 24780
rect 36428 23998 36430 24050
rect 36482 23998 36484 24050
rect 35420 23268 35476 23278
rect 35420 23266 35588 23268
rect 35420 23214 35422 23266
rect 35474 23214 35588 23266
rect 35420 23212 35588 23214
rect 35420 23202 35476 23212
rect 34076 23044 34132 23054
rect 34076 22950 34132 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 33628 22258 33684 22270
rect 33628 22206 33630 22258
rect 33682 22206 33684 22258
rect 33628 21476 33684 22206
rect 35532 22148 35588 23212
rect 35756 22484 35812 22494
rect 35756 22390 35812 22428
rect 35532 22082 35588 22092
rect 34300 21476 34356 21486
rect 33628 21474 34356 21476
rect 33628 21422 34302 21474
rect 34354 21422 34356 21474
rect 33628 21420 34356 21422
rect 34300 21410 34356 21420
rect 35868 21364 35924 23884
rect 36428 23828 36484 23998
rect 36428 23762 36484 23772
rect 36764 24610 36820 24622
rect 36764 24558 36766 24610
rect 36818 24558 36820 24610
rect 36428 23268 36484 23278
rect 36428 22484 36484 23212
rect 36764 23156 36820 24558
rect 36876 24052 36932 26852
rect 37100 24724 37156 24734
rect 37100 24630 37156 24668
rect 37100 24052 37156 24062
rect 36876 23996 37100 24052
rect 37100 23938 37156 23996
rect 37100 23886 37102 23938
rect 37154 23886 37156 23938
rect 37100 23874 37156 23886
rect 37212 23714 37268 23726
rect 37212 23662 37214 23714
rect 37266 23662 37268 23714
rect 37212 23604 37268 23662
rect 36764 23090 36820 23100
rect 36988 23548 37268 23604
rect 37324 23604 37380 27132
rect 37436 27074 37492 27916
rect 37436 27022 37438 27074
rect 37490 27022 37492 27074
rect 37436 27010 37492 27022
rect 37660 27858 37716 27870
rect 37660 27806 37662 27858
rect 37714 27806 37716 27858
rect 37436 26852 37492 26862
rect 37436 26402 37492 26796
rect 37436 26350 37438 26402
rect 37490 26350 37492 26402
rect 37436 26338 37492 26350
rect 37660 24612 37716 27806
rect 38108 27748 38164 27758
rect 38108 27654 38164 27692
rect 38332 27076 38388 27086
rect 38332 26982 38388 27020
rect 38556 26962 38612 27916
rect 38556 26910 38558 26962
rect 38610 26910 38612 26962
rect 38556 26898 38612 26910
rect 39004 27300 39060 27310
rect 39116 27300 39172 28140
rect 39060 27244 39172 27300
rect 39228 27748 39284 27758
rect 39004 26962 39060 27244
rect 39228 27076 39284 27692
rect 39228 27074 39620 27076
rect 39228 27022 39230 27074
rect 39282 27022 39620 27074
rect 39228 27020 39620 27022
rect 39228 27010 39284 27020
rect 39004 26910 39006 26962
rect 39058 26910 39060 26962
rect 39004 26898 39060 26910
rect 38332 26852 38388 26862
rect 38444 26852 38500 26862
rect 38388 26850 38500 26852
rect 38388 26798 38446 26850
rect 38498 26798 38500 26850
rect 38388 26796 38500 26798
rect 38332 26786 38388 26796
rect 38444 26786 38500 26796
rect 39564 26178 39620 27020
rect 39564 26126 39566 26178
rect 39618 26126 39620 26178
rect 39564 26114 39620 26126
rect 37660 24610 37828 24612
rect 37660 24558 37662 24610
rect 37714 24558 37828 24610
rect 37660 24556 37828 24558
rect 37660 24546 37716 24556
rect 37548 24052 37604 24062
rect 37548 24050 37716 24052
rect 37548 23998 37550 24050
rect 37602 23998 37716 24050
rect 37548 23996 37716 23998
rect 37548 23986 37604 23996
rect 37436 23940 37492 23950
rect 37436 23846 37492 23884
rect 37548 23828 37604 23838
rect 37548 23734 37604 23772
rect 37324 23548 37492 23604
rect 36092 22372 36148 22382
rect 36092 22258 36148 22316
rect 36428 22370 36484 22428
rect 36988 22482 37044 23548
rect 37100 23268 37156 23278
rect 37100 23174 37156 23212
rect 36988 22430 36990 22482
rect 37042 22430 37044 22482
rect 36988 22418 37044 22430
rect 37324 23156 37380 23166
rect 37324 22482 37380 23100
rect 37436 23042 37492 23548
rect 37436 22990 37438 23042
rect 37490 22990 37492 23042
rect 37436 22978 37492 22990
rect 37324 22430 37326 22482
rect 37378 22430 37380 22482
rect 37324 22418 37380 22430
rect 36428 22318 36430 22370
rect 36482 22318 36484 22370
rect 36428 22306 36484 22318
rect 37436 22372 37492 22382
rect 37436 22278 37492 22316
rect 36092 22206 36094 22258
rect 36146 22206 36148 22258
rect 36092 22036 36148 22206
rect 37660 22148 37716 23996
rect 37772 23492 37828 24556
rect 37772 22596 37828 23436
rect 38108 24052 38164 24062
rect 38108 22932 38164 23996
rect 38892 23828 38948 23838
rect 38220 23156 38276 23166
rect 38556 23156 38612 23166
rect 38220 23154 38612 23156
rect 38220 23102 38222 23154
rect 38274 23102 38558 23154
rect 38610 23102 38612 23154
rect 38220 23100 38612 23102
rect 38220 23090 38276 23100
rect 38556 23090 38612 23100
rect 38892 23154 38948 23772
rect 38892 23102 38894 23154
rect 38946 23102 38948 23154
rect 38108 22876 38500 22932
rect 37772 22530 37828 22540
rect 36092 21970 36148 21980
rect 37324 22092 37716 22148
rect 36652 21586 36708 21598
rect 36652 21534 36654 21586
rect 36706 21534 36708 21586
rect 36428 21476 36484 21486
rect 36652 21476 36708 21534
rect 36484 21420 36708 21476
rect 36428 21382 36484 21420
rect 35868 21298 35924 21308
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 37324 21028 37380 22092
rect 37436 21476 37492 21486
rect 37436 21474 37604 21476
rect 37436 21422 37438 21474
rect 37490 21422 37604 21474
rect 37436 21420 37604 21422
rect 37436 21410 37492 21420
rect 37436 21028 37492 21038
rect 37324 21026 37492 21028
rect 37324 20974 37438 21026
rect 37490 20974 37492 21026
rect 37324 20972 37492 20974
rect 37436 20962 37492 20972
rect 33068 20914 33460 20916
rect 33068 20862 33070 20914
rect 33122 20862 33460 20914
rect 33068 20860 33460 20862
rect 33068 20850 33124 20860
rect 33404 20802 33460 20860
rect 37548 20914 37604 21420
rect 37548 20862 37550 20914
rect 37602 20862 37604 20914
rect 37548 20850 37604 20862
rect 33404 20750 33406 20802
rect 33458 20750 33460 20802
rect 33404 20738 33460 20750
rect 37772 20802 37828 20814
rect 37772 20750 37774 20802
rect 37826 20750 37828 20802
rect 33740 20580 33796 20590
rect 33740 20486 33796 20524
rect 37100 20580 37156 20590
rect 37100 20486 37156 20524
rect 37772 20580 37828 20750
rect 37772 20514 37828 20524
rect 35756 20132 35812 20142
rect 35756 20018 35812 20076
rect 35756 19966 35758 20018
rect 35810 19966 35812 20018
rect 35756 19684 35812 19966
rect 35980 20130 36036 20142
rect 35980 20078 35982 20130
rect 36034 20078 36036 20130
rect 35980 19908 36036 20078
rect 35980 19842 36036 19852
rect 37548 19908 37604 19918
rect 35196 19628 35460 19638
rect 35756 19628 36372 19684
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 33404 19460 33460 19470
rect 33404 19366 33460 19404
rect 33404 19236 33460 19246
rect 33404 19142 33460 19180
rect 33740 19124 33796 19134
rect 33628 19122 33796 19124
rect 33628 19070 33742 19122
rect 33794 19070 33796 19122
rect 33628 19068 33796 19070
rect 33068 18674 33124 18686
rect 33068 18622 33070 18674
rect 33122 18622 33124 18674
rect 33068 18452 33124 18622
rect 33628 18452 33684 19068
rect 33740 19058 33796 19068
rect 36204 19124 36260 19134
rect 36204 19030 36260 19068
rect 36316 19122 36372 19628
rect 37548 19348 37604 19852
rect 37548 19254 37604 19292
rect 38332 19348 38388 19358
rect 36316 19070 36318 19122
rect 36370 19070 36372 19122
rect 36316 19058 36372 19070
rect 37324 19234 37380 19246
rect 37324 19182 37326 19234
rect 37378 19182 37380 19234
rect 37324 19124 37380 19182
rect 36540 19010 36596 19022
rect 36540 18958 36542 19010
rect 36594 18958 36596 19010
rect 35756 18562 35812 18574
rect 35756 18510 35758 18562
rect 35810 18510 35812 18562
rect 33068 18386 33124 18396
rect 33292 18396 33684 18452
rect 33740 18450 33796 18462
rect 33740 18398 33742 18450
rect 33794 18398 33796 18450
rect 33180 18228 33236 18238
rect 33292 18228 33348 18396
rect 33740 18340 33796 18398
rect 33628 18284 33796 18340
rect 33180 18226 33348 18228
rect 33180 18174 33182 18226
rect 33234 18174 33348 18226
rect 33180 18172 33348 18174
rect 33180 18162 33236 18172
rect 32956 17948 33236 18004
rect 31836 17612 32228 17668
rect 31612 17442 31780 17444
rect 31612 17390 31614 17442
rect 31666 17390 31780 17442
rect 31612 17388 31780 17390
rect 31612 17378 31668 17388
rect 31724 17108 31780 17388
rect 31724 17042 31780 17052
rect 31612 16994 31668 17006
rect 31612 16942 31614 16994
rect 31666 16942 31668 16994
rect 31612 16548 31668 16942
rect 31612 16482 31668 16492
rect 31836 16324 31892 17612
rect 32620 17556 32676 17566
rect 31948 17554 32676 17556
rect 31948 17502 32622 17554
rect 32674 17502 32676 17554
rect 31948 17500 32676 17502
rect 31948 16660 32004 17500
rect 32620 17490 32676 17500
rect 32060 17108 32116 17118
rect 32060 17014 32116 17052
rect 32172 16884 32228 16894
rect 32956 16884 33012 16894
rect 32172 16882 33012 16884
rect 32172 16830 32174 16882
rect 32226 16830 32958 16882
rect 33010 16830 33012 16882
rect 32172 16828 33012 16830
rect 32172 16818 32228 16828
rect 32956 16818 33012 16828
rect 32060 16660 32116 16670
rect 32284 16660 32340 16670
rect 31948 16658 32116 16660
rect 31948 16606 32062 16658
rect 32114 16606 32116 16658
rect 31948 16604 32116 16606
rect 32060 16594 32116 16604
rect 32172 16604 32284 16660
rect 31612 16212 31668 16222
rect 31836 16212 31892 16268
rect 31612 16210 31892 16212
rect 31612 16158 31614 16210
rect 31666 16158 31892 16210
rect 31612 16156 31892 16158
rect 31612 16146 31668 16156
rect 31948 15540 32004 15550
rect 31948 15314 32004 15484
rect 32060 15540 32116 15550
rect 32172 15540 32228 16604
rect 32284 16594 32340 16604
rect 32620 15988 32676 15998
rect 32060 15538 32228 15540
rect 32060 15486 32062 15538
rect 32114 15486 32228 15538
rect 32060 15484 32228 15486
rect 32508 15932 32620 15988
rect 32060 15474 32116 15484
rect 31948 15262 31950 15314
rect 32002 15262 32004 15314
rect 31948 15250 32004 15262
rect 32172 15316 32228 15326
rect 32508 15316 32564 15932
rect 32620 15922 32676 15932
rect 32172 15314 32564 15316
rect 32172 15262 32174 15314
rect 32226 15262 32564 15314
rect 32172 15260 32564 15262
rect 32172 15250 32228 15260
rect 32508 15148 32564 15260
rect 32620 15316 32676 15326
rect 32956 15316 33012 15326
rect 32620 15314 33012 15316
rect 32620 15262 32622 15314
rect 32674 15262 32958 15314
rect 33010 15262 33012 15314
rect 32620 15260 33012 15262
rect 32620 15250 32676 15260
rect 32956 15250 33012 15260
rect 31724 15092 31780 15102
rect 32508 15092 32676 15148
rect 31724 14642 31780 15036
rect 31724 14590 31726 14642
rect 31778 14590 31780 14642
rect 31724 14578 31780 14590
rect 32396 12964 32452 12974
rect 32284 12962 32452 12964
rect 32284 12910 32398 12962
rect 32450 12910 32452 12962
rect 32284 12908 32452 12910
rect 31500 12338 31556 12348
rect 31612 12850 31668 12862
rect 31612 12798 31614 12850
rect 31666 12798 31668 12850
rect 31612 12628 31668 12798
rect 31948 12852 32004 12862
rect 32172 12852 32228 12862
rect 31948 12850 32228 12852
rect 31948 12798 31950 12850
rect 32002 12798 32174 12850
rect 32226 12798 32228 12850
rect 31948 12796 32228 12798
rect 31948 12786 32004 12796
rect 32172 12786 32228 12796
rect 31612 12068 31668 12572
rect 31724 12738 31780 12750
rect 31724 12686 31726 12738
rect 31778 12686 31780 12738
rect 31724 12404 31780 12686
rect 32284 12628 32340 12908
rect 32396 12898 32452 12908
rect 32620 12964 32676 15092
rect 32620 12870 32676 12908
rect 32732 15092 32788 15102
rect 32396 12740 32452 12750
rect 32396 12646 32452 12684
rect 31724 12338 31780 12348
rect 32172 12572 32340 12628
rect 31612 12012 32004 12068
rect 31724 11282 31780 11294
rect 31724 11230 31726 11282
rect 31778 11230 31780 11282
rect 31724 10050 31780 11230
rect 31836 11170 31892 11182
rect 31836 11118 31838 11170
rect 31890 11118 31892 11170
rect 31836 10164 31892 11118
rect 31948 10610 32004 12012
rect 32060 11172 32116 11182
rect 32172 11172 32228 12572
rect 32732 12404 32788 15036
rect 33068 15092 33124 15102
rect 33068 13076 33124 15036
rect 33180 13970 33236 17948
rect 33292 17780 33348 18172
rect 33292 17714 33348 17724
rect 33404 18226 33460 18238
rect 33404 18174 33406 18226
rect 33458 18174 33460 18226
rect 33180 13918 33182 13970
rect 33234 13918 33236 13970
rect 33180 13524 33236 13918
rect 33292 16996 33348 17006
rect 33292 13860 33348 16940
rect 33404 15988 33460 18174
rect 33628 16548 33684 18284
rect 33740 18116 33796 18284
rect 33964 18340 34020 18350
rect 33964 18246 34020 18284
rect 34412 18338 34468 18350
rect 34412 18286 34414 18338
rect 34466 18286 34468 18338
rect 34412 18116 34468 18286
rect 33740 18060 34468 18116
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 34748 17780 34804 17790
rect 33628 16482 33684 16492
rect 33740 17778 34804 17780
rect 33740 17726 34750 17778
rect 34802 17726 34804 17778
rect 33740 17724 34804 17726
rect 33740 16210 33796 17724
rect 34748 17714 34804 17724
rect 35756 17444 35812 18510
rect 36092 18562 36148 18574
rect 36092 18510 36094 18562
rect 36146 18510 36148 18562
rect 35868 18450 35924 18462
rect 35868 18398 35870 18450
rect 35922 18398 35924 18450
rect 35868 17556 35924 18398
rect 35980 18340 36036 18350
rect 35980 18246 36036 18284
rect 36092 18116 36148 18510
rect 36316 18452 36372 18462
rect 36316 18358 36372 18396
rect 36092 18050 36148 18060
rect 36540 17892 36596 18958
rect 36540 17826 36596 17836
rect 36988 19010 37044 19022
rect 36988 18958 36990 19010
rect 37042 18958 37044 19010
rect 36988 17666 37044 18958
rect 37324 18564 37380 19068
rect 38332 18674 38388 19292
rect 38332 18622 38334 18674
rect 38386 18622 38388 18674
rect 38332 18610 38388 18622
rect 37100 18450 37156 18462
rect 37100 18398 37102 18450
rect 37154 18398 37156 18450
rect 37100 18340 37156 18398
rect 37100 18274 37156 18284
rect 37212 18226 37268 18238
rect 37212 18174 37214 18226
rect 37266 18174 37268 18226
rect 37212 18116 37268 18174
rect 37212 18050 37268 18060
rect 37212 17892 37268 17902
rect 37100 17780 37156 17790
rect 37100 17686 37156 17724
rect 36988 17614 36990 17666
rect 37042 17614 37044 17666
rect 36988 17602 37044 17614
rect 37212 17668 37268 17836
rect 37212 17574 37268 17612
rect 35868 17500 36708 17556
rect 35756 17378 35812 17388
rect 36652 17106 36708 17500
rect 37324 17444 37380 18508
rect 38108 18564 38164 18574
rect 38108 18470 38164 18508
rect 38220 18452 38276 18462
rect 38220 18358 38276 18396
rect 37548 18340 37604 18350
rect 37548 18338 37940 18340
rect 37548 18286 37550 18338
rect 37602 18286 37940 18338
rect 37548 18284 37940 18286
rect 37548 18274 37604 18284
rect 37436 18116 37492 18126
rect 37436 17668 37492 18060
rect 37884 17780 37940 18284
rect 37884 17724 38388 17780
rect 37436 17612 37940 17668
rect 37436 17554 37492 17612
rect 37436 17502 37438 17554
rect 37490 17502 37492 17554
rect 37436 17490 37492 17502
rect 37884 17554 37940 17612
rect 37884 17502 37886 17554
rect 37938 17502 37940 17554
rect 37884 17490 37940 17502
rect 37996 17556 38052 17566
rect 37996 17462 38052 17500
rect 36652 17054 36654 17106
rect 36706 17054 36708 17106
rect 36652 17042 36708 17054
rect 37100 17388 37380 17444
rect 37660 17444 37716 17454
rect 35308 16994 35364 17006
rect 35308 16942 35310 16994
rect 35362 16942 35364 16994
rect 35308 16884 35364 16942
rect 35308 16818 35364 16828
rect 35868 16772 35924 16782
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 33740 16158 33742 16210
rect 33794 16158 33796 16210
rect 33740 16146 33796 16158
rect 34636 16324 34692 16334
rect 34412 16100 34468 16110
rect 34412 16006 34468 16044
rect 33404 15922 33460 15932
rect 33292 13794 33348 13804
rect 34412 13860 34468 13870
rect 33740 13524 33796 13534
rect 33180 13458 33236 13468
rect 33292 13522 33796 13524
rect 33292 13470 33742 13522
rect 33794 13470 33796 13522
rect 33292 13468 33796 13470
rect 33180 13076 33236 13086
rect 33068 13074 33236 13076
rect 33068 13022 33182 13074
rect 33234 13022 33236 13074
rect 33068 13020 33236 13022
rect 33180 13010 33236 13020
rect 33292 12962 33348 13468
rect 33740 13458 33796 13468
rect 33628 13300 33684 13310
rect 33292 12910 33294 12962
rect 33346 12910 33348 12962
rect 33292 12898 33348 12910
rect 33404 12964 33460 12974
rect 33460 12908 33572 12964
rect 33404 12898 33460 12908
rect 33068 12740 33124 12750
rect 33068 12646 33124 12684
rect 33404 12740 33460 12750
rect 32732 12348 33348 12404
rect 33180 12178 33236 12190
rect 33180 12126 33182 12178
rect 33234 12126 33236 12178
rect 32620 11508 32676 11518
rect 32620 11506 33124 11508
rect 32620 11454 32622 11506
rect 32674 11454 33124 11506
rect 32620 11452 33124 11454
rect 32620 11442 32676 11452
rect 32116 11116 32228 11172
rect 32284 11282 32340 11294
rect 32284 11230 32286 11282
rect 32338 11230 32340 11282
rect 32060 11078 32116 11116
rect 32284 10612 32340 11230
rect 32508 11172 32564 11182
rect 31948 10558 31950 10610
rect 32002 10558 32004 10610
rect 31948 10546 32004 10558
rect 32060 10556 32340 10612
rect 32396 11170 32564 11172
rect 32396 11118 32510 11170
rect 32562 11118 32564 11170
rect 32396 11116 32564 11118
rect 31836 10098 31892 10108
rect 31724 9998 31726 10050
rect 31778 9998 31780 10050
rect 31724 9986 31780 9998
rect 32060 9940 32116 10556
rect 32396 10500 32452 11116
rect 32508 11106 32564 11116
rect 32508 10612 32564 10622
rect 32508 10518 32564 10556
rect 33068 10610 33124 11452
rect 33068 10558 33070 10610
rect 33122 10558 33124 10610
rect 33068 10546 33124 10558
rect 33180 11172 33236 12126
rect 33180 10612 33236 11116
rect 33292 10836 33348 12348
rect 33404 12402 33460 12684
rect 33404 12350 33406 12402
rect 33458 12350 33460 12402
rect 33404 12338 33460 12350
rect 33516 12404 33572 12908
rect 33628 12962 33684 13244
rect 34412 13074 34468 13804
rect 34412 13022 34414 13074
rect 34466 13022 34468 13074
rect 34412 13010 34468 13022
rect 33628 12910 33630 12962
rect 33682 12910 33684 12962
rect 33628 12898 33684 12910
rect 34188 12964 34244 12974
rect 34188 12870 34244 12908
rect 33964 12852 34020 12862
rect 33740 12850 34020 12852
rect 33740 12798 33966 12850
rect 34018 12798 34020 12850
rect 33740 12796 34020 12798
rect 33628 12404 33684 12414
rect 33516 12402 33684 12404
rect 33516 12350 33630 12402
rect 33682 12350 33684 12402
rect 33516 12348 33684 12350
rect 33628 12338 33684 12348
rect 33740 12402 33796 12796
rect 33964 12786 34020 12796
rect 34300 12852 34356 12862
rect 33740 12350 33742 12402
rect 33794 12350 33796 12402
rect 33740 12338 33796 12350
rect 33964 12404 34020 12414
rect 33964 12066 34020 12348
rect 33964 12014 33966 12066
rect 34018 12014 34020 12066
rect 33964 12002 34020 12014
rect 34076 12292 34132 12302
rect 34076 11844 34132 12236
rect 34300 11956 34356 12796
rect 34524 12850 34580 12862
rect 34524 12798 34526 12850
rect 34578 12798 34580 12850
rect 34524 12628 34580 12798
rect 34524 12562 34580 12572
rect 33852 11788 34132 11844
rect 34188 11954 34356 11956
rect 34188 11902 34302 11954
rect 34354 11902 34356 11954
rect 34188 11900 34356 11902
rect 33292 10780 33460 10836
rect 33292 10612 33348 10622
rect 33180 10610 33348 10612
rect 33180 10558 33294 10610
rect 33346 10558 33348 10610
rect 33180 10556 33348 10558
rect 33292 10546 33348 10556
rect 32284 10444 32452 10500
rect 31836 9884 32116 9940
rect 32172 10386 32228 10398
rect 32172 10334 32174 10386
rect 32226 10334 32228 10386
rect 32172 9940 32228 10334
rect 31836 9826 31892 9884
rect 32172 9874 32228 9884
rect 31836 9774 31838 9826
rect 31890 9774 31892 9826
rect 31724 9602 31780 9614
rect 31724 9550 31726 9602
rect 31778 9550 31780 9602
rect 31724 9492 31780 9550
rect 31724 9426 31780 9436
rect 31836 9156 31892 9774
rect 32172 9714 32228 9726
rect 32172 9662 32174 9714
rect 32226 9662 32228 9714
rect 32172 9604 32228 9662
rect 32284 9716 32340 10444
rect 32508 10276 32564 10286
rect 32396 10220 32508 10276
rect 32396 9826 32452 10220
rect 32508 10210 32564 10220
rect 33404 10052 33460 10780
rect 33516 10724 33572 10734
rect 33516 10388 33572 10668
rect 33740 10612 33796 10622
rect 33740 10518 33796 10556
rect 33516 10322 33572 10332
rect 33628 10498 33684 10510
rect 33628 10446 33630 10498
rect 33682 10446 33684 10498
rect 33628 10276 33684 10446
rect 33628 10210 33684 10220
rect 33516 10052 33572 10062
rect 33404 10050 33572 10052
rect 33404 9998 33518 10050
rect 33570 9998 33572 10050
rect 33404 9996 33572 9998
rect 33516 9986 33572 9996
rect 32732 9940 32788 9950
rect 33292 9940 33348 9950
rect 32732 9938 33236 9940
rect 32732 9886 32734 9938
rect 32786 9886 33236 9938
rect 32732 9884 33236 9886
rect 32732 9874 32788 9884
rect 32396 9774 32398 9826
rect 32450 9774 32452 9826
rect 32396 9762 32452 9774
rect 32508 9828 32564 9838
rect 32284 9650 32340 9660
rect 32172 9538 32228 9548
rect 31724 8930 31780 8942
rect 31724 8878 31726 8930
rect 31778 8878 31780 8930
rect 31612 8818 31668 8830
rect 31612 8766 31614 8818
rect 31666 8766 31668 8818
rect 31612 8260 31668 8766
rect 31500 8258 31668 8260
rect 31500 8206 31614 8258
rect 31666 8206 31668 8258
rect 31500 8204 31668 8206
rect 31500 7474 31556 8204
rect 31612 8194 31668 8204
rect 31724 7812 31780 8878
rect 31836 8370 31892 9100
rect 31836 8318 31838 8370
rect 31890 8318 31892 8370
rect 31836 8306 31892 8318
rect 31724 7746 31780 7756
rect 31948 8148 32004 8158
rect 32284 8148 32340 8158
rect 31948 8146 32340 8148
rect 31948 8094 31950 8146
rect 32002 8094 32286 8146
rect 32338 8094 32340 8146
rect 31948 8092 32340 8094
rect 31500 7422 31502 7474
rect 31554 7422 31556 7474
rect 31500 7410 31556 7422
rect 31948 6916 32004 8092
rect 32284 8082 32340 8092
rect 32396 8148 32452 8158
rect 32508 8148 32564 9772
rect 32620 9716 32676 9726
rect 32620 9622 32676 9660
rect 33068 9716 33124 9726
rect 32732 9602 32788 9614
rect 32732 9550 32734 9602
rect 32786 9550 32788 9602
rect 32732 9380 32788 9550
rect 32732 9314 32788 9324
rect 32844 9604 32900 9614
rect 32620 8372 32676 8382
rect 32620 8258 32676 8316
rect 32620 8206 32622 8258
rect 32674 8206 32676 8258
rect 32620 8194 32676 8206
rect 32396 8146 32564 8148
rect 32396 8094 32398 8146
rect 32450 8094 32564 8146
rect 32396 8092 32564 8094
rect 32732 8148 32788 8158
rect 32396 8082 32452 8092
rect 32732 7924 32788 8092
rect 32396 7868 32788 7924
rect 32172 7700 32228 7710
rect 32172 7606 32228 7644
rect 32396 7698 32452 7868
rect 32396 7646 32398 7698
rect 32450 7646 32452 7698
rect 32396 7634 32452 7646
rect 32508 7476 32564 7486
rect 32508 7382 32564 7420
rect 31948 6850 32004 6860
rect 31388 5182 31390 5234
rect 31442 5182 31444 5234
rect 31388 5170 31444 5182
rect 31612 6580 31668 6590
rect 29708 4562 29876 4564
rect 29708 4510 29710 4562
rect 29762 4510 29876 4562
rect 29708 4508 29876 4510
rect 31276 5124 31332 5134
rect 29708 4498 29764 4508
rect 29260 4286 29262 4338
rect 29314 4286 29316 4338
rect 29260 4274 29316 4286
rect 28700 3614 28702 3666
rect 28754 3614 28756 3666
rect 28700 3602 28756 3614
rect 31276 3554 31332 5068
rect 31276 3502 31278 3554
rect 31330 3502 31332 3554
rect 31276 3490 31332 3502
rect 31500 4226 31556 4238
rect 31500 4174 31502 4226
rect 31554 4174 31556 4226
rect 31500 3556 31556 4174
rect 31500 3490 31556 3500
rect 17948 3332 18228 3388
rect 18508 3444 18564 3482
rect 18508 3378 18564 3388
rect 31052 3444 31108 3482
rect 31052 3378 31108 3388
rect 31612 3442 31668 6524
rect 32284 6244 32340 6254
rect 32060 5908 32116 5918
rect 31948 5852 32060 5908
rect 31948 4900 32004 5852
rect 32060 5842 32116 5852
rect 32284 5794 32340 6188
rect 32284 5742 32286 5794
rect 32338 5742 32340 5794
rect 32060 5236 32116 5246
rect 32284 5236 32340 5742
rect 32732 5796 32788 5806
rect 32116 5180 32676 5236
rect 32060 5122 32116 5180
rect 32060 5070 32062 5122
rect 32114 5070 32116 5122
rect 32060 5058 32116 5070
rect 32620 5122 32676 5180
rect 32620 5070 32622 5122
rect 32674 5070 32676 5122
rect 32620 5058 32676 5070
rect 32732 4900 32788 5740
rect 31948 4844 32228 4900
rect 31948 4452 32004 4462
rect 31948 4358 32004 4396
rect 32172 4450 32228 4844
rect 32508 4844 32788 4900
rect 32508 4562 32564 4844
rect 32508 4510 32510 4562
rect 32562 4510 32564 4562
rect 32508 4498 32564 4510
rect 32620 4676 32676 4686
rect 32172 4398 32174 4450
rect 32226 4398 32228 4450
rect 32172 4386 32228 4398
rect 32620 3554 32676 4620
rect 32620 3502 32622 3554
rect 32674 3502 32676 3554
rect 32620 3490 32676 3502
rect 31612 3390 31614 3442
rect 31666 3390 31668 3442
rect 31612 3378 31668 3390
rect 32284 3442 32340 3454
rect 32284 3390 32286 3442
rect 32338 3390 32340 3442
rect 32284 3388 32340 3390
rect 32844 3388 32900 9548
rect 33068 9042 33124 9660
rect 33068 8990 33070 9042
rect 33122 8990 33124 9042
rect 33068 8978 33124 8990
rect 33180 8428 33236 9884
rect 33348 9884 33460 9940
rect 33292 9874 33348 9884
rect 33292 9604 33348 9614
rect 33292 9510 33348 9548
rect 33404 9380 33460 9884
rect 33404 9324 33572 9380
rect 33516 9268 33572 9324
rect 33628 9268 33684 9278
rect 33516 9266 33684 9268
rect 33516 9214 33630 9266
rect 33682 9214 33684 9266
rect 33516 9212 33684 9214
rect 33628 9202 33684 9212
rect 33516 9042 33572 9054
rect 33740 9044 33796 9054
rect 33516 8990 33518 9042
rect 33570 8990 33572 9042
rect 33180 8372 33348 8428
rect 33180 8258 33236 8270
rect 33180 8206 33182 8258
rect 33234 8206 33236 8258
rect 33180 7812 33236 8206
rect 33180 7746 33236 7756
rect 33292 6914 33348 8372
rect 33404 8260 33460 8270
rect 33404 8166 33460 8204
rect 33516 7812 33572 8990
rect 33516 7746 33572 7756
rect 33628 9042 33796 9044
rect 33628 8990 33742 9042
rect 33794 8990 33796 9042
rect 33628 8988 33796 8990
rect 33628 8258 33684 8988
rect 33740 8978 33796 8988
rect 33628 8206 33630 8258
rect 33682 8206 33684 8258
rect 33628 7476 33684 8206
rect 33852 7588 33908 11788
rect 33964 10500 34020 10510
rect 33964 8484 34020 10444
rect 34076 9156 34132 9166
rect 34076 9062 34132 9100
rect 34076 8484 34132 8494
rect 33964 8482 34132 8484
rect 33964 8430 34078 8482
rect 34130 8430 34132 8482
rect 33964 8428 34132 8430
rect 34076 8418 34132 8428
rect 33852 7522 33908 7532
rect 33628 7410 33684 7420
rect 33292 6862 33294 6914
rect 33346 6862 33348 6914
rect 33292 6850 33348 6862
rect 33852 7362 33908 7374
rect 33852 7310 33854 7362
rect 33906 7310 33908 7362
rect 33404 6466 33460 6478
rect 33404 6414 33406 6466
rect 33458 6414 33460 6466
rect 33404 6020 33460 6414
rect 33292 5964 33460 6020
rect 33516 6468 33572 6478
rect 33852 6468 33908 7310
rect 33516 6466 33852 6468
rect 33516 6414 33518 6466
rect 33570 6414 33852 6466
rect 33516 6412 33852 6414
rect 33292 5236 33348 5964
rect 33404 5796 33460 5806
rect 33516 5796 33572 6412
rect 33852 6374 33908 6412
rect 34188 6130 34244 11900
rect 34300 11890 34356 11900
rect 34300 9492 34356 9502
rect 34300 9266 34356 9436
rect 34300 9214 34302 9266
rect 34354 9214 34356 9266
rect 34300 8146 34356 9214
rect 34524 9268 34580 9278
rect 34636 9268 34692 16268
rect 35532 16324 35588 16334
rect 35532 16098 35588 16268
rect 35532 16046 35534 16098
rect 35586 16046 35588 16098
rect 35532 16034 35588 16046
rect 34860 15988 34916 15998
rect 34860 15894 34916 15932
rect 35196 15988 35252 15998
rect 35196 15894 35252 15932
rect 35868 15988 35924 16716
rect 36988 16658 37044 16670
rect 36988 16606 36990 16658
rect 37042 16606 37044 16658
rect 36988 16210 37044 16606
rect 36988 16158 36990 16210
rect 37042 16158 37044 16210
rect 36988 16146 37044 16158
rect 35308 15426 35364 15438
rect 35308 15374 35310 15426
rect 35362 15374 35364 15426
rect 35308 15092 35364 15374
rect 35868 15148 35924 15932
rect 36316 16100 36372 16110
rect 36316 15540 36372 16044
rect 36316 15538 36708 15540
rect 36316 15486 36318 15538
rect 36370 15486 36708 15538
rect 36316 15484 36708 15486
rect 36316 15474 36372 15484
rect 36652 15314 36708 15484
rect 36652 15262 36654 15314
rect 36706 15262 36708 15314
rect 36652 15250 36708 15262
rect 37100 15148 37156 17388
rect 37660 17350 37716 17388
rect 37212 16772 37268 16782
rect 37212 16678 37268 16716
rect 38332 16324 38388 17724
rect 35868 15092 36260 15148
rect 35308 15026 35364 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35532 14420 35588 14430
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34860 12962 34916 12974
rect 34860 12910 34862 12962
rect 34914 12910 34916 12962
rect 34748 12852 34804 12862
rect 34860 12852 34916 12910
rect 34804 12796 34916 12852
rect 34972 12964 35028 12974
rect 34748 12786 34804 12796
rect 34972 12738 35028 12908
rect 34972 12686 34974 12738
rect 35026 12686 35028 12738
rect 34860 12628 34916 12638
rect 34860 12402 34916 12572
rect 34860 12350 34862 12402
rect 34914 12350 34916 12402
rect 34860 12338 34916 12350
rect 34860 10610 34916 10622
rect 34860 10558 34862 10610
rect 34914 10558 34916 10610
rect 34860 9828 34916 10558
rect 34860 9762 34916 9772
rect 34524 9266 34804 9268
rect 34524 9214 34526 9266
rect 34578 9214 34804 9266
rect 34524 9212 34804 9214
rect 34524 9202 34580 9212
rect 34636 9044 34692 9054
rect 34636 8950 34692 8988
rect 34524 8260 34580 8270
rect 34524 8166 34580 8204
rect 34300 8094 34302 8146
rect 34354 8094 34356 8146
rect 34300 8082 34356 8094
rect 34412 6916 34468 6926
rect 34412 6690 34468 6860
rect 34412 6638 34414 6690
rect 34466 6638 34468 6690
rect 34412 6626 34468 6638
rect 34748 6690 34804 9212
rect 34972 8148 35028 12686
rect 35196 12740 35252 12750
rect 35196 12646 35252 12684
rect 35084 12178 35140 12190
rect 35084 12126 35086 12178
rect 35138 12126 35140 12178
rect 35084 10500 35140 12126
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35532 11620 35588 14364
rect 35868 13860 35924 13870
rect 35868 13766 35924 13804
rect 35644 12964 35700 12974
rect 35644 11788 35700 12908
rect 35868 12628 35924 12638
rect 35868 12290 35924 12572
rect 35868 12238 35870 12290
rect 35922 12238 35924 12290
rect 35868 12226 35924 12238
rect 36204 12180 36260 15092
rect 36988 15092 37156 15148
rect 37212 16268 38388 16324
rect 36428 13972 36484 13982
rect 36428 13074 36484 13916
rect 36428 13022 36430 13074
rect 36482 13022 36484 13074
rect 36204 12178 36372 12180
rect 36204 12126 36206 12178
rect 36258 12126 36372 12178
rect 36204 12124 36372 12126
rect 36204 12114 36260 12124
rect 36204 11954 36260 11966
rect 36204 11902 36206 11954
rect 36258 11902 36260 11954
rect 35644 11732 35812 11788
rect 35532 11282 35588 11564
rect 35532 11230 35534 11282
rect 35586 11230 35588 11282
rect 35532 11218 35588 11230
rect 35420 11172 35476 11182
rect 35420 10834 35476 11116
rect 35420 10782 35422 10834
rect 35474 10782 35476 10834
rect 35420 10770 35476 10782
rect 35308 10612 35364 10622
rect 35308 10518 35364 10556
rect 35532 10610 35588 10622
rect 35532 10558 35534 10610
rect 35586 10558 35588 10610
rect 35084 10434 35140 10444
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35532 9044 35588 10558
rect 35756 10612 35812 11732
rect 35644 9714 35700 9726
rect 35644 9662 35646 9714
rect 35698 9662 35700 9714
rect 35644 9604 35700 9662
rect 35644 9538 35700 9548
rect 35756 9266 35812 10556
rect 35756 9214 35758 9266
rect 35810 9214 35812 9266
rect 35756 9202 35812 9214
rect 35868 11170 35924 11182
rect 35868 11118 35870 11170
rect 35922 11118 35924 11170
rect 35868 9268 35924 11118
rect 36204 10836 36260 11902
rect 36204 10770 36260 10780
rect 36316 10610 36372 12124
rect 36428 11508 36484 13022
rect 36764 13524 36820 13534
rect 36428 11506 36708 11508
rect 36428 11454 36430 11506
rect 36482 11454 36708 11506
rect 36428 11452 36708 11454
rect 36428 11442 36484 11452
rect 36316 10558 36318 10610
rect 36370 10558 36372 10610
rect 36316 10546 36372 10558
rect 36540 10948 36596 10958
rect 36540 10610 36596 10892
rect 36540 10558 36542 10610
rect 36594 10558 36596 10610
rect 36540 10546 36596 10558
rect 35980 10500 36036 10510
rect 35980 10406 36036 10444
rect 36428 10164 36484 10174
rect 36316 9828 36372 9838
rect 36316 9492 36372 9772
rect 35868 9212 36036 9268
rect 35532 8978 35588 8988
rect 35868 9042 35924 9054
rect 35868 8990 35870 9042
rect 35922 8990 35924 9042
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35868 8372 35924 8990
rect 35980 8820 36036 9212
rect 36316 9266 36372 9436
rect 36316 9214 36318 9266
rect 36370 9214 36372 9266
rect 36316 9202 36372 9214
rect 36204 9044 36260 9054
rect 36204 8950 36260 8988
rect 35980 8754 36036 8764
rect 36316 8820 36372 8830
rect 36428 8820 36484 10108
rect 36316 8818 36484 8820
rect 36316 8766 36318 8818
rect 36370 8766 36484 8818
rect 36316 8764 36484 8766
rect 36540 9940 36596 9950
rect 36540 9156 36596 9884
rect 36652 9828 36708 11452
rect 36652 9762 36708 9772
rect 36316 8754 36372 8764
rect 34972 8082 35028 8092
rect 35756 8260 35812 8270
rect 35644 7588 35700 7598
rect 35644 7494 35700 7532
rect 35308 7364 35364 7374
rect 35308 7362 35588 7364
rect 35308 7310 35310 7362
rect 35362 7310 35588 7362
rect 35308 7308 35588 7310
rect 35308 7298 35364 7308
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34748 6638 34750 6690
rect 34802 6638 34804 6690
rect 34748 6626 34804 6638
rect 34860 6692 34916 6702
rect 34300 6580 34356 6590
rect 34300 6486 34356 6524
rect 34860 6578 34916 6636
rect 34860 6526 34862 6578
rect 34914 6526 34916 6578
rect 34860 6514 34916 6526
rect 35532 6244 35588 7308
rect 35756 6692 35812 8204
rect 35532 6178 35588 6188
rect 35644 6690 35812 6692
rect 35644 6638 35758 6690
rect 35810 6638 35812 6690
rect 35644 6636 35812 6638
rect 34188 6078 34190 6130
rect 34242 6078 34244 6130
rect 34188 6066 34244 6078
rect 35644 6020 35700 6636
rect 35756 6626 35812 6636
rect 35868 6692 35924 8316
rect 36428 8484 36484 8494
rect 36316 8260 36372 8270
rect 36204 8146 36260 8158
rect 36204 8094 36206 8146
rect 36258 8094 36260 8146
rect 35980 7588 36036 7598
rect 35980 7494 36036 7532
rect 36204 6804 36260 8094
rect 36316 8146 36372 8204
rect 36316 8094 36318 8146
rect 36370 8094 36372 8146
rect 36316 8082 36372 8094
rect 36204 6738 36260 6748
rect 36316 7924 36372 7934
rect 35924 6636 36036 6692
rect 35868 6626 35924 6636
rect 35868 6466 35924 6478
rect 35868 6414 35870 6466
rect 35922 6414 35924 6466
rect 35532 5964 35700 6020
rect 35756 6018 35812 6030
rect 35756 5966 35758 6018
rect 35810 5966 35812 6018
rect 33404 5794 33572 5796
rect 33404 5742 33406 5794
rect 33458 5742 33572 5794
rect 33404 5740 33572 5742
rect 33628 5796 33684 5806
rect 33404 5730 33460 5740
rect 33628 5702 33684 5740
rect 34524 5794 34580 5806
rect 34524 5742 34526 5794
rect 34578 5742 34580 5794
rect 33852 5684 33908 5694
rect 33852 5590 33908 5628
rect 33404 5236 33460 5246
rect 33292 5234 33460 5236
rect 33292 5182 33406 5234
rect 33458 5182 33460 5234
rect 33292 5180 33460 5182
rect 33404 5170 33460 5180
rect 34524 5124 34580 5742
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35532 5234 35588 5964
rect 35532 5182 35534 5234
rect 35586 5182 35588 5234
rect 35532 5170 35588 5182
rect 35644 5348 35700 5358
rect 35308 5124 35364 5134
rect 34524 5058 34580 5068
rect 35196 5068 35308 5124
rect 34076 5012 34132 5022
rect 33516 4452 33572 4462
rect 33516 4358 33572 4396
rect 19852 3332 19908 3342
rect 20860 3332 20916 3342
rect 22204 3332 22260 3342
rect 32284 3332 32900 3388
rect 33404 3556 33460 3566
rect 33404 3442 33460 3500
rect 33404 3390 33406 3442
rect 33458 3390 33460 3442
rect 33404 3378 33460 3390
rect 17948 800 18004 3332
rect 19292 3330 19908 3332
rect 19292 3278 19854 3330
rect 19906 3278 19908 3330
rect 19292 3276 19908 3278
rect 19292 800 19348 3276
rect 19852 3266 19908 3276
rect 20636 3330 20916 3332
rect 20636 3278 20862 3330
rect 20914 3278 20916 3330
rect 20636 3276 20916 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20636 800 20692 3276
rect 20860 3266 20916 3276
rect 21980 3330 22260 3332
rect 21980 3278 22206 3330
rect 22258 3278 22260 3330
rect 21980 3276 22260 3278
rect 21980 800 22036 3276
rect 22204 3266 22260 3276
rect 34076 800 34132 4956
rect 34524 4788 34580 4798
rect 34524 4226 34580 4732
rect 35196 4450 35252 5068
rect 35308 5058 35364 5068
rect 35196 4398 35198 4450
rect 35250 4398 35252 4450
rect 35196 4386 35252 4398
rect 34524 4174 34526 4226
rect 34578 4174 34580 4226
rect 34524 4162 34580 4174
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35532 3780 35588 3790
rect 35644 3780 35700 5292
rect 35532 3778 35700 3780
rect 35532 3726 35534 3778
rect 35586 3726 35700 3778
rect 35532 3724 35700 3726
rect 35756 3780 35812 5966
rect 35868 5684 35924 6414
rect 35980 6356 36036 6636
rect 36316 6578 36372 7868
rect 36316 6526 36318 6578
rect 36370 6526 36372 6578
rect 36316 6514 36372 6526
rect 35980 6290 36036 6300
rect 35868 5346 35924 5628
rect 35868 5294 35870 5346
rect 35922 5294 35924 5346
rect 35868 5282 35924 5294
rect 35980 5796 36036 5806
rect 35980 5124 36036 5740
rect 36204 5682 36260 5694
rect 36204 5630 36206 5682
rect 36258 5630 36260 5682
rect 36204 5124 36260 5630
rect 35980 5068 36148 5124
rect 36092 5010 36148 5068
rect 36204 5058 36260 5068
rect 36092 4958 36094 5010
rect 36146 4958 36148 5010
rect 36092 4946 36148 4958
rect 35980 4900 36036 4910
rect 35980 4806 36036 4844
rect 36316 4228 36372 4238
rect 36428 4228 36484 8428
rect 36540 8258 36596 9100
rect 36540 8206 36542 8258
rect 36594 8206 36596 8258
rect 36540 8194 36596 8206
rect 36652 8260 36708 8270
rect 36652 8036 36708 8204
rect 36652 7970 36708 7980
rect 36540 7362 36596 7374
rect 36540 7310 36542 7362
rect 36594 7310 36596 7362
rect 36540 5908 36596 7310
rect 36764 6468 36820 13468
rect 36988 12964 37044 15092
rect 37212 14644 37268 16268
rect 37436 16100 37492 16110
rect 37436 16006 37492 16044
rect 37884 16100 37940 16110
rect 37884 16098 38164 16100
rect 37884 16046 37886 16098
rect 37938 16046 38164 16098
rect 37884 16044 38164 16046
rect 37884 16034 37940 16044
rect 37436 15202 37492 15214
rect 37436 15150 37438 15202
rect 37490 15150 37492 15202
rect 37436 14756 37492 15150
rect 38108 15148 38164 16044
rect 38332 15986 38388 16268
rect 38332 15934 38334 15986
rect 38386 15934 38388 15986
rect 38332 15922 38388 15934
rect 38108 15092 38276 15148
rect 37436 14700 38052 14756
rect 37212 14588 37828 14644
rect 37100 14308 37156 14318
rect 37100 13970 37156 14252
rect 37100 13918 37102 13970
rect 37154 13918 37156 13970
rect 37100 13412 37156 13918
rect 37212 13970 37268 14588
rect 37212 13918 37214 13970
rect 37266 13918 37268 13970
rect 37212 13906 37268 13918
rect 37324 14418 37380 14430
rect 37324 14366 37326 14418
rect 37378 14366 37380 14418
rect 37324 13970 37380 14366
rect 37324 13918 37326 13970
rect 37378 13918 37380 13970
rect 37324 13906 37380 13918
rect 37660 13972 37716 13982
rect 37436 13860 37492 13870
rect 37436 13766 37492 13804
rect 37660 13858 37716 13916
rect 37660 13806 37662 13858
rect 37714 13806 37716 13858
rect 37660 13794 37716 13806
rect 37324 13748 37380 13758
rect 37100 13356 37268 13412
rect 36988 12898 37044 12908
rect 37212 12962 37268 13356
rect 37212 12910 37214 12962
rect 37266 12910 37268 12962
rect 37212 12898 37268 12910
rect 36988 12738 37044 12750
rect 37324 12740 37380 13692
rect 37660 13076 37716 13086
rect 36988 12686 36990 12738
rect 37042 12686 37044 12738
rect 36988 12404 37044 12686
rect 36876 12348 37044 12404
rect 37100 12684 37380 12740
rect 37436 13074 37716 13076
rect 37436 13022 37662 13074
rect 37714 13022 37716 13074
rect 37436 13020 37716 13022
rect 37100 12402 37156 12684
rect 37100 12350 37102 12402
rect 37154 12350 37156 12402
rect 36876 10164 36932 12348
rect 37100 12338 37156 12350
rect 37212 12292 37268 12302
rect 37212 12198 37268 12236
rect 36988 12178 37044 12190
rect 36988 12126 36990 12178
rect 37042 12126 37044 12178
rect 36988 11170 37044 12126
rect 37436 12178 37492 13020
rect 37660 13010 37716 13020
rect 37772 12852 37828 14588
rect 37772 12758 37828 12796
rect 37884 14532 37940 14542
rect 37436 12126 37438 12178
rect 37490 12126 37492 12178
rect 37436 12114 37492 12126
rect 37548 12290 37604 12302
rect 37548 12238 37550 12290
rect 37602 12238 37604 12290
rect 37324 12068 37380 12078
rect 37100 12012 37324 12068
rect 37100 11506 37156 12012
rect 37324 12002 37380 12012
rect 37548 11732 37604 12238
rect 37884 11788 37940 14476
rect 37996 13634 38052 14700
rect 37996 13582 37998 13634
rect 38050 13582 38052 13634
rect 37996 13570 38052 13582
rect 38108 14196 38164 14206
rect 38108 13858 38164 14140
rect 38108 13806 38110 13858
rect 38162 13806 38164 13858
rect 38108 13524 38164 13806
rect 38108 13458 38164 13468
rect 37100 11454 37102 11506
rect 37154 11454 37156 11506
rect 37100 11442 37156 11454
rect 37436 11676 37604 11732
rect 37660 11732 37940 11788
rect 37996 12850 38052 12862
rect 37996 12798 37998 12850
rect 38050 12798 38052 12850
rect 36988 11118 36990 11170
rect 37042 11118 37044 11170
rect 36988 10386 37044 11118
rect 36988 10334 36990 10386
rect 37042 10334 37044 10386
rect 36988 10322 37044 10334
rect 37212 11170 37268 11182
rect 37212 11118 37214 11170
rect 37266 11118 37268 11170
rect 36876 10108 37044 10164
rect 36988 9828 37044 10108
rect 37212 9940 37268 11118
rect 37436 11172 37492 11676
rect 37660 11396 37716 11732
rect 37884 11620 37940 11630
rect 37996 11620 38052 12798
rect 37884 11618 37996 11620
rect 37884 11566 37886 11618
rect 37938 11566 37996 11618
rect 37884 11564 37996 11566
rect 37884 11554 37940 11564
rect 37996 11526 38052 11564
rect 37436 11078 37492 11116
rect 37548 11340 37716 11396
rect 38108 11508 38164 11518
rect 37436 10836 37492 10846
rect 37436 10742 37492 10780
rect 37548 10164 37604 11340
rect 38108 11282 38164 11452
rect 38108 11230 38110 11282
rect 38162 11230 38164 11282
rect 37660 11172 37716 11182
rect 37660 10834 37716 11116
rect 37996 11170 38052 11182
rect 37996 11118 37998 11170
rect 38050 11118 38052 11170
rect 37884 10948 37940 10958
rect 37660 10782 37662 10834
rect 37714 10782 37716 10834
rect 37660 10770 37716 10782
rect 37772 10892 37884 10948
rect 37772 10388 37828 10892
rect 37884 10882 37940 10892
rect 37884 10612 37940 10622
rect 37996 10612 38052 11118
rect 38108 10948 38164 11230
rect 38108 10882 38164 10892
rect 38220 10724 38276 15092
rect 38332 14308 38388 14318
rect 38332 13858 38388 14252
rect 38444 13972 38500 22876
rect 38892 21476 38948 23102
rect 39116 23042 39172 23054
rect 39116 22990 39118 23042
rect 39170 22990 39172 23042
rect 39116 22596 39172 22990
rect 39116 22530 39172 22540
rect 38892 21410 38948 21420
rect 39564 21476 39620 21486
rect 39564 21382 39620 21420
rect 38556 20580 38612 20590
rect 38556 16324 38612 20524
rect 38556 16268 38724 16324
rect 38556 16098 38612 16110
rect 38556 16046 38558 16098
rect 38610 16046 38612 16098
rect 38556 15204 38612 16046
rect 38556 15138 38612 15148
rect 38556 14196 38612 14206
rect 38668 14196 38724 16268
rect 39564 15204 39620 15214
rect 39564 15110 39620 15148
rect 39676 14308 39732 14318
rect 39676 14214 39732 14252
rect 38612 14140 38724 14196
rect 38556 14130 38612 14140
rect 38444 13906 38500 13916
rect 38332 13806 38334 13858
rect 38386 13806 38388 13858
rect 38332 13794 38388 13806
rect 38556 13860 38612 13870
rect 38780 13860 38836 13870
rect 38556 13766 38612 13804
rect 38668 13858 38836 13860
rect 38668 13806 38782 13858
rect 38834 13806 38836 13858
rect 38668 13804 38836 13806
rect 38668 13412 38724 13804
rect 38780 13794 38836 13804
rect 38892 13748 38948 13758
rect 38892 13654 38948 13692
rect 39340 13634 39396 13646
rect 39340 13582 39342 13634
rect 39394 13582 39396 13634
rect 39340 13524 39396 13582
rect 39340 13458 39396 13468
rect 38444 13356 38724 13412
rect 38444 13186 38500 13356
rect 38444 13134 38446 13186
rect 38498 13134 38500 13186
rect 38444 13122 38500 13134
rect 38332 12850 38388 12862
rect 38332 12798 38334 12850
rect 38386 12798 38388 12850
rect 38332 12068 38388 12798
rect 38444 12852 38500 12862
rect 38444 12758 38500 12796
rect 38332 12002 38388 12012
rect 38556 11508 38612 11518
rect 38612 11452 38724 11508
rect 38556 11442 38612 11452
rect 38556 11282 38612 11294
rect 38556 11230 38558 11282
rect 38610 11230 38612 11282
rect 38444 10836 38500 10846
rect 38556 10836 38612 11230
rect 38668 11282 38724 11452
rect 38668 11230 38670 11282
rect 38722 11230 38724 11282
rect 38668 11218 38724 11230
rect 38892 11172 38948 11182
rect 38892 11170 39060 11172
rect 38892 11118 38894 11170
rect 38946 11118 39060 11170
rect 38892 11116 39060 11118
rect 38892 11106 38948 11116
rect 38668 10836 38724 10846
rect 38556 10834 38724 10836
rect 38556 10782 38670 10834
rect 38722 10782 38724 10834
rect 38556 10780 38724 10782
rect 38220 10668 38388 10724
rect 37884 10610 38052 10612
rect 37884 10558 37886 10610
rect 37938 10558 38052 10610
rect 37884 10556 38052 10558
rect 38108 10610 38164 10622
rect 38108 10558 38110 10610
rect 38162 10558 38164 10610
rect 37884 10546 37940 10556
rect 37772 10332 38052 10388
rect 37548 10108 37940 10164
rect 37212 9874 37268 9884
rect 37548 9828 37604 9838
rect 36988 9826 37156 9828
rect 36988 9774 36990 9826
rect 37042 9774 37156 9826
rect 36988 9772 37156 9774
rect 36988 9762 37044 9772
rect 37100 9380 37156 9772
rect 37548 9734 37604 9772
rect 37212 9604 37268 9614
rect 37212 9510 37268 9548
rect 37324 9602 37380 9614
rect 37324 9550 37326 9602
rect 37378 9550 37380 9602
rect 37324 9380 37380 9550
rect 37436 9604 37492 9614
rect 37436 9510 37492 9548
rect 37100 9314 37156 9324
rect 37212 9324 37380 9380
rect 37772 9380 37828 9390
rect 36988 9156 37044 9166
rect 36988 9062 37044 9100
rect 36876 8820 36932 8830
rect 36876 7924 36932 8764
rect 36988 8148 37044 8158
rect 36988 8054 37044 8092
rect 37100 8034 37156 8046
rect 37100 7982 37102 8034
rect 37154 7982 37156 8034
rect 37100 7924 37156 7982
rect 37212 8036 37268 9324
rect 37324 9156 37380 9166
rect 37324 9062 37380 9100
rect 37660 9154 37716 9166
rect 37660 9102 37662 9154
rect 37714 9102 37716 9154
rect 37324 8260 37380 8270
rect 37324 8166 37380 8204
rect 37548 8146 37604 8158
rect 37548 8094 37550 8146
rect 37602 8094 37604 8146
rect 37212 7980 37492 8036
rect 36876 7868 37044 7924
rect 37100 7868 37380 7924
rect 36988 7812 37044 7868
rect 36988 7756 37156 7812
rect 36764 6402 36820 6412
rect 36876 6804 36932 6814
rect 36988 6804 37044 6814
rect 36932 6802 37044 6804
rect 36932 6750 36990 6802
rect 37042 6750 37044 6802
rect 36932 6748 37044 6750
rect 36540 5842 36596 5852
rect 36652 6244 36708 6254
rect 36876 6244 36932 6748
rect 36988 6738 37044 6748
rect 37100 6802 37156 7756
rect 37100 6750 37102 6802
rect 37154 6750 37156 6802
rect 37100 6738 37156 6750
rect 37212 7588 37268 7598
rect 37212 6578 37268 7532
rect 37212 6526 37214 6578
rect 37266 6526 37268 6578
rect 37212 6514 37268 6526
rect 36652 4338 36708 6188
rect 36764 6188 36932 6244
rect 36764 4900 36820 6188
rect 37324 6132 37380 7868
rect 37324 6066 37380 6076
rect 37100 5012 37156 5022
rect 37100 4918 37156 4956
rect 36764 4834 36820 4844
rect 37436 4900 37492 7980
rect 37548 6580 37604 8094
rect 37660 7924 37716 9102
rect 37772 8372 37828 9324
rect 37884 8708 37940 10108
rect 37996 9716 38052 10332
rect 38108 10164 38164 10558
rect 38108 10098 38164 10108
rect 38220 10498 38276 10510
rect 38220 10446 38222 10498
rect 38274 10446 38276 10498
rect 38220 9828 38276 10446
rect 38332 10500 38388 10668
rect 38444 10612 38500 10780
rect 38668 10770 38724 10780
rect 38780 10724 38836 10734
rect 38780 10630 38836 10668
rect 38556 10612 38612 10622
rect 38444 10610 38612 10612
rect 38444 10558 38558 10610
rect 38610 10558 38612 10610
rect 38444 10556 38612 10558
rect 38556 10546 38612 10556
rect 38332 10444 38500 10500
rect 38220 9762 38276 9772
rect 37996 9622 38052 9660
rect 38332 9604 38388 9614
rect 38220 9602 38388 9604
rect 38220 9550 38334 9602
rect 38386 9550 38388 9602
rect 38220 9548 38388 9550
rect 38108 9380 38164 9390
rect 38220 9380 38276 9548
rect 38332 9538 38388 9548
rect 38164 9324 38276 9380
rect 38108 9314 38164 9324
rect 38444 9268 38500 10444
rect 39004 9716 39060 11116
rect 39116 10610 39172 10622
rect 39116 10558 39118 10610
rect 39170 10558 39172 10610
rect 39116 10164 39172 10558
rect 39116 10098 39172 10108
rect 39228 9828 39284 9838
rect 39228 9734 39284 9772
rect 39116 9716 39172 9726
rect 39004 9714 39172 9716
rect 39004 9662 39118 9714
rect 39170 9662 39172 9714
rect 39004 9660 39172 9662
rect 39116 9650 39172 9660
rect 38892 9604 38948 9614
rect 38892 9510 38948 9548
rect 39004 9492 39060 9502
rect 38444 9212 38724 9268
rect 37996 9154 38052 9166
rect 37996 9102 37998 9154
rect 38050 9102 38052 9154
rect 37996 9044 38052 9102
rect 38332 9156 38388 9194
rect 38332 9090 38388 9100
rect 38556 9044 38612 9054
rect 37996 8988 38276 9044
rect 37884 8652 38164 8708
rect 37772 8258 37828 8316
rect 37772 8206 37774 8258
rect 37826 8206 37828 8258
rect 37772 8194 37828 8206
rect 37996 8372 38052 8382
rect 37660 7868 37940 7924
rect 37548 6514 37604 6524
rect 37660 7586 37716 7598
rect 37660 7534 37662 7586
rect 37714 7534 37716 7586
rect 37660 5236 37716 7534
rect 37660 5170 37716 5180
rect 37772 6466 37828 6478
rect 37772 6414 37774 6466
rect 37826 6414 37828 6466
rect 37772 5012 37828 6414
rect 37884 6244 37940 7868
rect 37996 7588 38052 8316
rect 38108 8258 38164 8652
rect 38108 8206 38110 8258
rect 38162 8206 38164 8258
rect 38108 8148 38164 8206
rect 38108 8082 38164 8092
rect 37996 7522 38052 7532
rect 37884 6178 37940 6188
rect 38108 7362 38164 7374
rect 38108 7310 38110 7362
rect 38162 7310 38164 7362
rect 37772 4946 37828 4956
rect 37436 4834 37492 4844
rect 38108 4676 38164 7310
rect 38220 6802 38276 8988
rect 38444 9042 38612 9044
rect 38444 8990 38558 9042
rect 38610 8990 38612 9042
rect 38444 8988 38612 8990
rect 38332 8484 38388 8494
rect 38444 8484 38500 8988
rect 38556 8978 38612 8988
rect 38668 8820 38724 9212
rect 39004 9266 39060 9436
rect 39004 9214 39006 9266
rect 39058 9214 39060 9266
rect 39004 9202 39060 9214
rect 38388 8428 38500 8484
rect 38556 8764 38724 8820
rect 39228 9042 39284 9054
rect 39228 8990 39230 9042
rect 39282 8990 39284 9042
rect 38556 8428 38612 8764
rect 38332 8418 38388 8428
rect 38556 8372 38948 8428
rect 38556 8260 38612 8372
rect 38556 8194 38612 8204
rect 38892 8258 38948 8372
rect 39228 8372 39284 8990
rect 39228 8306 39284 8316
rect 38892 8206 38894 8258
rect 38946 8206 38948 8258
rect 38892 8194 38948 8206
rect 39004 8146 39060 8158
rect 39004 8094 39006 8146
rect 39058 8094 39060 8146
rect 38220 6750 38222 6802
rect 38274 6750 38276 6802
rect 38220 6738 38276 6750
rect 38556 8034 38612 8046
rect 38556 7982 38558 8034
rect 38610 7982 38612 8034
rect 38108 4610 38164 4620
rect 38332 6020 38388 6030
rect 38556 6020 38612 7982
rect 39004 6916 39060 8094
rect 39228 8036 39284 8046
rect 39228 7942 39284 7980
rect 39004 6850 39060 6860
rect 39228 7586 39284 7598
rect 39228 7534 39230 7586
rect 39282 7534 39284 7586
rect 38332 6018 38612 6020
rect 38332 5966 38334 6018
rect 38386 5966 38612 6018
rect 38332 5964 38612 5966
rect 38892 6692 38948 6702
rect 36652 4286 36654 4338
rect 36706 4286 36708 4338
rect 36652 4274 36708 4286
rect 36764 4452 36820 4462
rect 36316 4226 36484 4228
rect 36316 4174 36318 4226
rect 36370 4174 36484 4226
rect 36316 4172 36484 4174
rect 36316 4162 36372 4172
rect 35868 3780 35924 3790
rect 35756 3778 35924 3780
rect 35756 3726 35870 3778
rect 35922 3726 35924 3778
rect 35756 3724 35924 3726
rect 35532 3714 35588 3724
rect 35868 3714 35924 3724
rect 35420 3444 35476 3454
rect 35420 800 35476 3388
rect 36764 800 36820 4396
rect 37436 4228 37492 4238
rect 37436 4134 37492 4172
rect 37996 3444 38052 3482
rect 38332 3388 38388 5964
rect 38892 5124 38948 6636
rect 39116 6580 39172 6590
rect 39004 6578 39172 6580
rect 39004 6526 39118 6578
rect 39170 6526 39172 6578
rect 39004 6524 39172 6526
rect 39004 5348 39060 6524
rect 39116 6514 39172 6524
rect 39116 6356 39172 6366
rect 39116 6130 39172 6300
rect 39116 6078 39118 6130
rect 39170 6078 39172 6130
rect 39116 6066 39172 6078
rect 39228 5460 39284 7534
rect 39340 6132 39396 6142
rect 39340 5908 39396 6076
rect 39340 5906 39620 5908
rect 39340 5854 39342 5906
rect 39394 5854 39620 5906
rect 39340 5852 39620 5854
rect 39340 5842 39396 5852
rect 39004 5282 39060 5292
rect 39116 5404 39284 5460
rect 38892 5068 39060 5124
rect 38780 5012 38836 5022
rect 38780 3778 38836 4956
rect 38780 3726 38782 3778
rect 38834 3726 38836 3778
rect 38780 3714 38836 3726
rect 38892 4228 38948 4238
rect 38892 3666 38948 4172
rect 38892 3614 38894 3666
rect 38946 3614 38948 3666
rect 38892 3602 38948 3614
rect 37996 3378 38052 3388
rect 38108 3332 38388 3388
rect 39004 3442 39060 5068
rect 39116 4788 39172 5404
rect 39228 5236 39284 5246
rect 39228 5142 39284 5180
rect 39116 4722 39172 4732
rect 39564 4226 39620 5852
rect 39564 4174 39566 4226
rect 39618 4174 39620 4226
rect 39564 4162 39620 4174
rect 39004 3390 39006 3442
rect 39058 3390 39060 3442
rect 39004 3378 39060 3390
rect 39452 3444 39508 3454
rect 38108 800 38164 3332
rect 39452 800 39508 3388
rect 1792 0 1904 800
rect 3136 0 3248 800
rect 4480 0 4592 800
rect 5824 0 5936 800
rect 7168 0 7280 800
rect 8512 0 8624 800
rect 9856 0 9968 800
rect 11200 0 11312 800
rect 12544 0 12656 800
rect 13888 0 14000 800
rect 15232 0 15344 800
rect 16576 0 16688 800
rect 17920 0 18032 800
rect 19264 0 19376 800
rect 20608 0 20720 800
rect 21952 0 22064 800
rect 23296 0 23408 800
rect 24640 0 24752 800
rect 25984 0 26096 800
rect 27328 0 27440 800
rect 28672 0 28784 800
rect 30016 0 30128 800
rect 31360 0 31472 800
rect 32704 0 32816 800
rect 34048 0 34160 800
rect 35392 0 35504 800
rect 36736 0 36848 800
rect 38080 0 38192 800
rect 39424 0 39536 800
<< via2 >>
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 17724 39676 17780 39732
rect 11788 39004 11844 39060
rect 9996 38780 10052 38836
rect 11340 38780 11396 38836
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 9660 38220 9716 38276
rect 10556 38220 10612 38276
rect 9996 38162 10052 38164
rect 9996 38110 9998 38162
rect 9998 38110 10050 38162
rect 10050 38110 10052 38162
rect 9996 38108 10052 38110
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 5628 35196 5684 35252
rect 6188 35196 6244 35252
rect 6412 35026 6468 35028
rect 6412 34974 6414 35026
rect 6414 34974 6466 35026
rect 6466 34974 6468 35026
rect 6412 34972 6468 34974
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 1932 29426 1988 29428
rect 1932 29374 1934 29426
rect 1934 29374 1986 29426
rect 1986 29374 1988 29426
rect 1932 29372 1988 29374
rect 8988 35084 9044 35140
rect 9660 35196 9716 35252
rect 6860 33404 6916 33460
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 3612 30380 3668 30436
rect 2828 29372 2884 29428
rect 5180 29372 5236 29428
rect 4732 29314 4788 29316
rect 4732 29262 4734 29314
rect 4734 29262 4786 29314
rect 4786 29262 4788 29314
rect 4732 29260 4788 29262
rect 6748 29484 6804 29540
rect 6636 29260 6692 29316
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 1820 26908 1876 26964
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3836 26908 3892 26964
rect 4620 26236 4676 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 3276 23884 3332 23940
rect 3500 24722 3556 24724
rect 3500 24670 3502 24722
rect 3502 24670 3554 24722
rect 3554 24670 3556 24722
rect 3500 24668 3556 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 6748 27746 6804 27748
rect 6748 27694 6750 27746
rect 6750 27694 6802 27746
rect 6802 27694 6804 27746
rect 6748 27692 6804 27694
rect 5068 26962 5124 26964
rect 5068 26910 5070 26962
rect 5070 26910 5122 26962
rect 5122 26910 5124 26962
rect 5068 26908 5124 26910
rect 6860 26572 6916 26628
rect 6412 26290 6468 26292
rect 6412 26238 6414 26290
rect 6414 26238 6466 26290
rect 6466 26238 6468 26290
rect 6412 26236 6468 26238
rect 6412 25452 6468 25508
rect 8204 33234 8260 33236
rect 8204 33182 8206 33234
rect 8206 33182 8258 33234
rect 8258 33182 8260 33234
rect 8204 33180 8260 33182
rect 7196 31106 7252 31108
rect 7196 31054 7198 31106
rect 7198 31054 7250 31106
rect 7250 31054 7252 31106
rect 7196 31052 7252 31054
rect 9324 33346 9380 33348
rect 9324 33294 9326 33346
rect 9326 33294 9378 33346
rect 9378 33294 9380 33346
rect 9324 33292 9380 33294
rect 9548 33964 9604 34020
rect 8428 31052 8484 31108
rect 8764 31164 8820 31220
rect 8540 30994 8596 30996
rect 8540 30942 8542 30994
rect 8542 30942 8594 30994
rect 8594 30942 8596 30994
rect 8540 30940 8596 30942
rect 7980 28812 8036 28868
rect 5740 24892 5796 24948
rect 4956 24780 5012 24836
rect 5964 24834 6020 24836
rect 5964 24782 5966 24834
rect 5966 24782 6018 24834
rect 6018 24782 6020 24834
rect 5964 24780 6020 24782
rect 4396 23938 4452 23940
rect 4396 23886 4398 23938
rect 4398 23886 4450 23938
rect 4450 23886 4452 23938
rect 4396 23884 4452 23886
rect 4844 23938 4900 23940
rect 4844 23886 4846 23938
rect 4846 23886 4898 23938
rect 4898 23886 4900 23938
rect 4844 23884 4900 23886
rect 5628 23884 5684 23940
rect 3500 22876 3556 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 6076 23100 6132 23156
rect 5852 22428 5908 22484
rect 5964 22316 6020 22372
rect 5068 22092 5124 22148
rect 5852 22092 5908 22148
rect 6524 24668 6580 24724
rect 6972 24668 7028 24724
rect 7196 26962 7252 26964
rect 7196 26910 7198 26962
rect 7198 26910 7250 26962
rect 7250 26910 7252 26962
rect 7196 26908 7252 26910
rect 8764 30268 8820 30324
rect 8652 29372 8708 29428
rect 8428 29260 8484 29316
rect 8540 28754 8596 28756
rect 8540 28702 8542 28754
rect 8542 28702 8594 28754
rect 8594 28702 8596 28754
rect 8540 28700 8596 28702
rect 8876 28812 8932 28868
rect 8764 28588 8820 28644
rect 8428 28028 8484 28084
rect 9660 33180 9716 33236
rect 11676 38722 11732 38724
rect 11676 38670 11678 38722
rect 11678 38670 11730 38722
rect 11730 38670 11732 38722
rect 11676 38668 11732 38670
rect 10444 34018 10500 34020
rect 10444 33966 10446 34018
rect 10446 33966 10498 34018
rect 10498 33966 10500 34018
rect 10444 33964 10500 33966
rect 11564 37996 11620 38052
rect 11564 36316 11620 36372
rect 12908 39004 12964 39060
rect 13580 39004 13636 39060
rect 15372 39004 15428 39060
rect 12684 38834 12740 38836
rect 12684 38782 12686 38834
rect 12686 38782 12738 38834
rect 12738 38782 12740 38834
rect 12684 38780 12740 38782
rect 12012 38668 12068 38724
rect 11788 35196 11844 35252
rect 11564 34300 11620 34356
rect 11340 33964 11396 34020
rect 11340 33516 11396 33572
rect 9996 33180 10052 33236
rect 9660 31106 9716 31108
rect 9660 31054 9662 31106
rect 9662 31054 9714 31106
rect 9714 31054 9716 31106
rect 9660 31052 9716 31054
rect 9324 30156 9380 30212
rect 11228 31836 11284 31892
rect 9996 30940 10052 30996
rect 10108 30268 10164 30324
rect 10220 30210 10276 30212
rect 10220 30158 10222 30210
rect 10222 30158 10274 30210
rect 10274 30158 10276 30210
rect 10220 30156 10276 30158
rect 9884 29372 9940 29428
rect 10108 29932 10164 29988
rect 11228 31164 11284 31220
rect 9100 29260 9156 29316
rect 10108 29260 10164 29316
rect 10556 29708 10612 29764
rect 10668 29596 10724 29652
rect 10332 29426 10388 29428
rect 10332 29374 10334 29426
rect 10334 29374 10386 29426
rect 10386 29374 10388 29426
rect 10332 29372 10388 29374
rect 9436 28754 9492 28756
rect 9436 28702 9438 28754
rect 9438 28702 9490 28754
rect 9490 28702 9492 28754
rect 9436 28700 9492 28702
rect 8988 28082 9044 28084
rect 8988 28030 8990 28082
rect 8990 28030 9042 28082
rect 9042 28030 9044 28082
rect 8988 28028 9044 28030
rect 9548 28642 9604 28644
rect 9548 28590 9550 28642
rect 9550 28590 9602 28642
rect 9602 28590 9604 28642
rect 9548 28588 9604 28590
rect 10220 28642 10276 28644
rect 10220 28590 10222 28642
rect 10222 28590 10274 28642
rect 10274 28590 10276 28642
rect 10220 28588 10276 28590
rect 9212 27804 9268 27860
rect 7532 26572 7588 26628
rect 7308 25506 7364 25508
rect 7308 25454 7310 25506
rect 7310 25454 7362 25506
rect 7362 25454 7364 25506
rect 7308 25452 7364 25454
rect 7868 24892 7924 24948
rect 7196 24556 7252 24612
rect 7644 24668 7700 24724
rect 6300 22428 6356 22484
rect 6748 22370 6804 22372
rect 6748 22318 6750 22370
rect 6750 22318 6802 22370
rect 6802 22318 6804 22370
rect 6748 22316 6804 22318
rect 3724 21586 3780 21588
rect 3724 21534 3726 21586
rect 3726 21534 3778 21586
rect 3778 21534 3780 21586
rect 3724 21532 3780 21534
rect 5068 21586 5124 21588
rect 5068 21534 5070 21586
rect 5070 21534 5122 21586
rect 5122 21534 5124 21586
rect 5068 21532 5124 21534
rect 4956 21308 5012 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5404 21308 5460 21364
rect 5516 20636 5572 20692
rect 2492 19068 2548 19124
rect 1820 17666 1876 17668
rect 1820 17614 1822 17666
rect 1822 17614 1874 17666
rect 1874 17614 1876 17666
rect 1820 17612 1876 17614
rect 1932 16828 1988 16884
rect 2828 15314 2884 15316
rect 2828 15262 2830 15314
rect 2830 15262 2882 15314
rect 2882 15262 2884 15314
rect 2828 15260 2884 15262
rect 1932 13580 1988 13636
rect 1932 6412 1988 6468
rect 2268 13580 2324 13636
rect 3948 20076 4004 20132
rect 5068 19964 5124 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 3500 19122 3556 19124
rect 3500 19070 3502 19122
rect 3502 19070 3554 19122
rect 3554 19070 3556 19122
rect 3500 19068 3556 19070
rect 3612 18844 3668 18900
rect 3052 16716 3108 16772
rect 4732 19180 4788 19236
rect 4396 18844 4452 18900
rect 5068 18508 5124 18564
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4620 17778 4676 17780
rect 4620 17726 4622 17778
rect 4622 17726 4674 17778
rect 4674 17726 4676 17778
rect 4620 17724 4676 17726
rect 5068 17612 5124 17668
rect 4172 16716 4228 16772
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 3276 15820 3332 15876
rect 3500 15260 3556 15316
rect 3500 14754 3556 14756
rect 3500 14702 3502 14754
rect 3502 14702 3554 14754
rect 3554 14702 3556 14754
rect 3500 14700 3556 14702
rect 4060 15874 4116 15876
rect 4060 15822 4062 15874
rect 4062 15822 4114 15874
rect 4114 15822 4116 15874
rect 4060 15820 4116 15822
rect 4284 15820 4340 15876
rect 4956 15820 5012 15876
rect 4956 15484 5012 15540
rect 4060 15148 4116 15204
rect 4396 15314 4452 15316
rect 4396 15262 4398 15314
rect 4398 15262 4450 15314
rect 4450 15262 4452 15314
rect 4396 15260 4452 15262
rect 5068 15426 5124 15428
rect 5068 15374 5070 15426
rect 5070 15374 5122 15426
rect 5122 15374 5124 15426
rect 5068 15372 5124 15374
rect 3164 9660 3220 9716
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4508 14700 4564 14756
rect 4956 14530 5012 14532
rect 4956 14478 4958 14530
rect 4958 14478 5010 14530
rect 5010 14478 5012 14530
rect 4956 14476 5012 14478
rect 5292 15148 5348 15204
rect 5180 13634 5236 13636
rect 5180 13582 5182 13634
rect 5182 13582 5234 13634
rect 5234 13582 5236 13634
rect 5180 13580 5236 13582
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4060 9714 4116 9716
rect 4060 9662 4062 9714
rect 4062 9662 4114 9714
rect 4114 9662 4116 9714
rect 4060 9660 4116 9662
rect 4620 8764 4676 8820
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 5068 8146 5124 8148
rect 5068 8094 5070 8146
rect 5070 8094 5122 8146
rect 5122 8094 5124 8146
rect 5068 8092 5124 8094
rect 3724 7644 3780 7700
rect 4956 7644 5012 7700
rect 6860 21868 6916 21924
rect 7084 23436 7140 23492
rect 7196 22540 7252 22596
rect 7980 23436 8036 23492
rect 7980 23154 8036 23156
rect 7980 23102 7982 23154
rect 7982 23102 8034 23154
rect 8034 23102 8036 23154
rect 7980 23100 8036 23102
rect 7756 22988 7812 23044
rect 7756 22540 7812 22596
rect 7084 22204 7140 22260
rect 7084 21532 7140 21588
rect 7308 22146 7364 22148
rect 7308 22094 7310 22146
rect 7310 22094 7362 22146
rect 7362 22094 7364 22146
rect 7308 22092 7364 22094
rect 7420 20914 7476 20916
rect 7420 20862 7422 20914
rect 7422 20862 7474 20914
rect 7474 20862 7476 20914
rect 7420 20860 7476 20862
rect 6412 20524 6468 20580
rect 5628 20076 5684 20132
rect 6524 20018 6580 20020
rect 6524 19966 6526 20018
rect 6526 19966 6578 20018
rect 6578 19966 6580 20018
rect 6524 19964 6580 19966
rect 5740 17666 5796 17668
rect 5740 17614 5742 17666
rect 5742 17614 5794 17666
rect 5794 17614 5796 17666
rect 5740 17612 5796 17614
rect 6188 19234 6244 19236
rect 6188 19182 6190 19234
rect 6190 19182 6242 19234
rect 6242 19182 6244 19234
rect 6188 19180 6244 19182
rect 5964 18508 6020 18564
rect 5852 16716 5908 16772
rect 6076 16322 6132 16324
rect 6076 16270 6078 16322
rect 6078 16270 6130 16322
rect 6130 16270 6132 16322
rect 6076 16268 6132 16270
rect 5628 15426 5684 15428
rect 5628 15374 5630 15426
rect 5630 15374 5682 15426
rect 5682 15374 5684 15426
rect 5628 15372 5684 15374
rect 6076 15538 6132 15540
rect 6076 15486 6078 15538
rect 6078 15486 6130 15538
rect 6130 15486 6132 15538
rect 6076 15484 6132 15486
rect 6188 15820 6244 15876
rect 5852 15148 5908 15204
rect 7644 21308 7700 21364
rect 7084 20578 7140 20580
rect 7084 20526 7086 20578
rect 7086 20526 7138 20578
rect 7138 20526 7140 20578
rect 7084 20524 7140 20526
rect 8316 24556 8372 24612
rect 8428 23938 8484 23940
rect 8428 23886 8430 23938
rect 8430 23886 8482 23938
rect 8482 23886 8484 23938
rect 8428 23884 8484 23886
rect 8316 22930 8372 22932
rect 8316 22878 8318 22930
rect 8318 22878 8370 22930
rect 8370 22878 8372 22930
rect 8316 22876 8372 22878
rect 8204 22652 8260 22708
rect 8204 22482 8260 22484
rect 8204 22430 8206 22482
rect 8206 22430 8258 22482
rect 8258 22430 8260 22482
rect 8204 22428 8260 22430
rect 9436 28476 9492 28532
rect 10668 28754 10724 28756
rect 10668 28702 10670 28754
rect 10670 28702 10722 28754
rect 10722 28702 10724 28754
rect 10668 28700 10724 28702
rect 10332 28476 10388 28532
rect 10444 27858 10500 27860
rect 10444 27806 10446 27858
rect 10446 27806 10498 27858
rect 10498 27806 10500 27858
rect 10444 27804 10500 27806
rect 9436 27692 9492 27748
rect 7980 21644 8036 21700
rect 7756 20748 7812 20804
rect 9212 21980 9268 22036
rect 8764 21644 8820 21700
rect 8540 21308 8596 21364
rect 8652 20802 8708 20804
rect 8652 20750 8654 20802
rect 8654 20750 8706 20802
rect 8706 20750 8708 20802
rect 8652 20748 8708 20750
rect 8316 20690 8372 20692
rect 8316 20638 8318 20690
rect 8318 20638 8370 20690
rect 8370 20638 8372 20690
rect 8316 20636 8372 20638
rect 8876 20972 8932 21028
rect 8764 20188 8820 20244
rect 8204 20076 8260 20132
rect 7756 19180 7812 19236
rect 12012 38220 12068 38276
rect 12236 38610 12292 38612
rect 12236 38558 12238 38610
rect 12238 38558 12290 38610
rect 12290 38558 12292 38610
rect 12236 38556 12292 38558
rect 13132 38444 13188 38500
rect 12348 37938 12404 37940
rect 12348 37886 12350 37938
rect 12350 37886 12402 37938
rect 12402 37886 12404 37938
rect 12348 37884 12404 37886
rect 12236 37436 12292 37492
rect 13468 37938 13524 37940
rect 13468 37886 13470 37938
rect 13470 37886 13522 37938
rect 13522 37886 13524 37938
rect 13468 37884 13524 37886
rect 13020 37826 13076 37828
rect 13020 37774 13022 37826
rect 13022 37774 13074 37826
rect 13074 37774 13076 37826
rect 13020 37772 13076 37774
rect 12796 37660 12852 37716
rect 13804 38556 13860 38612
rect 14700 38108 14756 38164
rect 13916 38050 13972 38052
rect 13916 37998 13918 38050
rect 13918 37998 13970 38050
rect 13970 37998 13972 38050
rect 13916 37996 13972 37998
rect 13692 37826 13748 37828
rect 13692 37774 13694 37826
rect 13694 37774 13746 37826
rect 13746 37774 13748 37826
rect 13692 37772 13748 37774
rect 13580 37660 13636 37716
rect 13468 37490 13524 37492
rect 13468 37438 13470 37490
rect 13470 37438 13522 37490
rect 13522 37438 13524 37490
rect 13468 37436 13524 37438
rect 13356 36428 13412 36484
rect 13916 37266 13972 37268
rect 13916 37214 13918 37266
rect 13918 37214 13970 37266
rect 13970 37214 13972 37266
rect 13916 37212 13972 37214
rect 14140 38050 14196 38052
rect 14140 37998 14142 38050
rect 14142 37998 14194 38050
rect 14194 37998 14196 38050
rect 14140 37996 14196 37998
rect 16156 38108 16212 38164
rect 15932 38050 15988 38052
rect 15932 37998 15934 38050
rect 15934 37998 15986 38050
rect 15986 37998 15988 38050
rect 15932 37996 15988 37998
rect 16604 38780 16660 38836
rect 16492 38444 16548 38500
rect 16492 38108 16548 38164
rect 16268 37826 16324 37828
rect 16268 37774 16270 37826
rect 16270 37774 16322 37826
rect 16322 37774 16324 37826
rect 16268 37772 16324 37774
rect 15036 37548 15092 37604
rect 14364 37266 14420 37268
rect 14364 37214 14366 37266
rect 14366 37214 14418 37266
rect 14418 37214 14420 37266
rect 14364 37212 14420 37214
rect 13468 36370 13524 36372
rect 13468 36318 13470 36370
rect 13470 36318 13522 36370
rect 13522 36318 13524 36370
rect 13468 36316 13524 36318
rect 12012 34972 12068 35028
rect 12124 35084 12180 35140
rect 11788 31836 11844 31892
rect 11564 31778 11620 31780
rect 11564 31726 11566 31778
rect 11566 31726 11618 31778
rect 11618 31726 11620 31778
rect 11564 31724 11620 31726
rect 11228 29932 11284 29988
rect 12012 31836 12068 31892
rect 13804 35756 13860 35812
rect 12348 35586 12404 35588
rect 12348 35534 12350 35586
rect 12350 35534 12402 35586
rect 12402 35534 12404 35586
rect 12348 35532 12404 35534
rect 12908 34802 12964 34804
rect 12908 34750 12910 34802
rect 12910 34750 12962 34802
rect 12962 34750 12964 34802
rect 12908 34748 12964 34750
rect 12460 34412 12516 34468
rect 12796 34354 12852 34356
rect 12796 34302 12798 34354
rect 12798 34302 12850 34354
rect 12850 34302 12852 34354
rect 12796 34300 12852 34302
rect 13468 34300 13524 34356
rect 12124 31778 12180 31780
rect 12124 31726 12126 31778
rect 12126 31726 12178 31778
rect 12178 31726 12180 31778
rect 12124 31724 12180 31726
rect 11676 30044 11732 30100
rect 11564 29708 11620 29764
rect 10892 28812 10948 28868
rect 11116 29260 11172 29316
rect 11340 29650 11396 29652
rect 11340 29598 11342 29650
rect 11342 29598 11394 29650
rect 11394 29598 11396 29650
rect 11340 29596 11396 29598
rect 11676 29202 11732 29204
rect 11676 29150 11678 29202
rect 11678 29150 11730 29202
rect 11730 29150 11732 29202
rect 11676 29148 11732 29150
rect 10892 28364 10948 28420
rect 11228 28700 11284 28756
rect 9772 27186 9828 27188
rect 9772 27134 9774 27186
rect 9774 27134 9826 27186
rect 9826 27134 9828 27186
rect 9772 27132 9828 27134
rect 10444 27186 10500 27188
rect 10444 27134 10446 27186
rect 10446 27134 10498 27186
rect 10498 27134 10500 27186
rect 10444 27132 10500 27134
rect 11452 28812 11508 28868
rect 11900 28924 11956 28980
rect 12124 28700 12180 28756
rect 12012 28642 12068 28644
rect 12012 28590 12014 28642
rect 12014 28590 12066 28642
rect 12066 28590 12068 28642
rect 12012 28588 12068 28590
rect 12348 28530 12404 28532
rect 12348 28478 12350 28530
rect 12350 28478 12402 28530
rect 12402 28478 12404 28530
rect 12348 28476 12404 28478
rect 12236 27132 12292 27188
rect 13580 34188 13636 34244
rect 12796 33516 12852 33572
rect 12572 33234 12628 33236
rect 12572 33182 12574 33234
rect 12574 33182 12626 33234
rect 12626 33182 12628 33234
rect 12572 33180 12628 33182
rect 12572 31890 12628 31892
rect 12572 31838 12574 31890
rect 12574 31838 12626 31890
rect 12626 31838 12628 31890
rect 12572 31836 12628 31838
rect 12684 31724 12740 31780
rect 13916 33516 13972 33572
rect 14028 36428 14084 36484
rect 14476 35810 14532 35812
rect 14476 35758 14478 35810
rect 14478 35758 14530 35810
rect 14530 35758 14532 35810
rect 14476 35756 14532 35758
rect 14700 35810 14756 35812
rect 14700 35758 14702 35810
rect 14702 35758 14754 35810
rect 14754 35758 14756 35810
rect 14700 35756 14756 35758
rect 14140 35698 14196 35700
rect 14140 35646 14142 35698
rect 14142 35646 14194 35698
rect 14194 35646 14196 35698
rect 14140 35644 14196 35646
rect 14364 35586 14420 35588
rect 14364 35534 14366 35586
rect 14366 35534 14418 35586
rect 14418 35534 14420 35586
rect 14364 35532 14420 35534
rect 14140 34412 14196 34468
rect 14140 34130 14196 34132
rect 14140 34078 14142 34130
rect 14142 34078 14194 34130
rect 14194 34078 14196 34130
rect 14140 34076 14196 34078
rect 14924 34914 14980 34916
rect 14924 34862 14926 34914
rect 14926 34862 14978 34914
rect 14978 34862 14980 34914
rect 14924 34860 14980 34862
rect 14812 34802 14868 34804
rect 14812 34750 14814 34802
rect 14814 34750 14866 34802
rect 14866 34750 14868 34802
rect 14812 34748 14868 34750
rect 14924 34636 14980 34692
rect 14700 34242 14756 34244
rect 14700 34190 14702 34242
rect 14702 34190 14754 34242
rect 14754 34190 14756 34242
rect 14700 34188 14756 34190
rect 14588 34130 14644 34132
rect 14588 34078 14590 34130
rect 14590 34078 14642 34130
rect 14642 34078 14644 34130
rect 14588 34076 14644 34078
rect 14140 33180 14196 33236
rect 14252 33346 14308 33348
rect 14252 33294 14254 33346
rect 14254 33294 14306 33346
rect 14306 33294 14308 33346
rect 14252 33292 14308 33294
rect 14028 31836 14084 31892
rect 13580 31500 13636 31556
rect 13468 28642 13524 28644
rect 13468 28590 13470 28642
rect 13470 28590 13522 28642
rect 13522 28590 13524 28642
rect 13468 28588 13524 28590
rect 12460 26908 12516 26964
rect 13468 28364 13524 28420
rect 10332 22988 10388 23044
rect 9884 22370 9940 22372
rect 9884 22318 9886 22370
rect 9886 22318 9938 22370
rect 9938 22318 9940 22370
rect 9884 22316 9940 22318
rect 9996 22258 10052 22260
rect 9996 22206 9998 22258
rect 9998 22206 10050 22258
rect 10050 22206 10052 22258
rect 9996 22204 10052 22206
rect 9548 21980 9604 22036
rect 9548 21698 9604 21700
rect 9548 21646 9550 21698
rect 9550 21646 9602 21698
rect 9602 21646 9604 21698
rect 9548 21644 9604 21646
rect 9548 21026 9604 21028
rect 9548 20974 9550 21026
rect 9550 20974 9602 21026
rect 9602 20974 9604 21026
rect 9548 20972 9604 20974
rect 10780 22258 10836 22260
rect 10780 22206 10782 22258
rect 10782 22206 10834 22258
rect 10834 22206 10836 22258
rect 10780 22204 10836 22206
rect 10444 21756 10500 21812
rect 9772 20972 9828 21028
rect 10444 20802 10500 20804
rect 10444 20750 10446 20802
rect 10446 20750 10498 20802
rect 10498 20750 10500 20802
rect 10444 20748 10500 20750
rect 10332 20524 10388 20580
rect 9772 20188 9828 20244
rect 9436 19516 9492 19572
rect 8428 19180 8484 19236
rect 8540 17612 8596 17668
rect 7644 17500 7700 17556
rect 8428 17554 8484 17556
rect 8428 17502 8430 17554
rect 8430 17502 8482 17554
rect 8482 17502 8484 17554
rect 8428 17500 8484 17502
rect 9212 19122 9268 19124
rect 9212 19070 9214 19122
rect 9214 19070 9266 19122
rect 9266 19070 9268 19122
rect 9212 19068 9268 19070
rect 10220 19068 10276 19124
rect 7308 16716 7364 16772
rect 7756 16716 7812 16772
rect 6972 16268 7028 16324
rect 7644 16268 7700 16324
rect 7420 15874 7476 15876
rect 7420 15822 7422 15874
rect 7422 15822 7474 15874
rect 7474 15822 7476 15874
rect 7420 15820 7476 15822
rect 7308 15484 7364 15540
rect 6860 15314 6916 15316
rect 6860 15262 6862 15314
rect 6862 15262 6914 15314
rect 6914 15262 6916 15314
rect 6860 15260 6916 15262
rect 6524 15148 6580 15204
rect 6748 15036 6804 15092
rect 5628 13580 5684 13636
rect 5964 11564 6020 11620
rect 6748 11564 6804 11620
rect 6188 11170 6244 11172
rect 6188 11118 6190 11170
rect 6190 11118 6242 11170
rect 6242 11118 6244 11170
rect 6188 11116 6244 11118
rect 5516 8428 5572 8484
rect 5964 8988 6020 9044
rect 5628 8146 5684 8148
rect 5628 8094 5630 8146
rect 5630 8094 5682 8146
rect 5682 8094 5684 8146
rect 5628 8092 5684 8094
rect 6524 10780 6580 10836
rect 6300 8988 6356 9044
rect 7196 15148 7252 15204
rect 13020 26124 13076 26180
rect 16156 34636 16212 34692
rect 15036 34076 15092 34132
rect 15596 34130 15652 34132
rect 15596 34078 15598 34130
rect 15598 34078 15650 34130
rect 15650 34078 15652 34130
rect 15596 34076 15652 34078
rect 15708 33346 15764 33348
rect 15708 33294 15710 33346
rect 15710 33294 15762 33346
rect 15762 33294 15764 33346
rect 15708 33292 15764 33294
rect 14588 33068 14644 33124
rect 13804 31164 13860 31220
rect 13692 30940 13748 30996
rect 14028 30268 14084 30324
rect 13804 29986 13860 29988
rect 13804 29934 13806 29986
rect 13806 29934 13858 29986
rect 13858 29934 13860 29986
rect 13804 29932 13860 29934
rect 14364 30210 14420 30212
rect 14364 30158 14366 30210
rect 14366 30158 14418 30210
rect 14418 30158 14420 30210
rect 14364 30156 14420 30158
rect 14476 30098 14532 30100
rect 14476 30046 14478 30098
rect 14478 30046 14530 30098
rect 14530 30046 14532 30098
rect 14476 30044 14532 30046
rect 14252 29986 14308 29988
rect 14252 29934 14254 29986
rect 14254 29934 14306 29986
rect 14306 29934 14308 29986
rect 14252 29932 14308 29934
rect 14364 29372 14420 29428
rect 13804 29260 13860 29316
rect 13692 29148 13748 29204
rect 13916 28642 13972 28644
rect 13916 28590 13918 28642
rect 13918 28590 13970 28642
rect 13970 28590 13972 28642
rect 13916 28588 13972 28590
rect 14364 29036 14420 29092
rect 15596 33122 15652 33124
rect 15596 33070 15598 33122
rect 15598 33070 15650 33122
rect 15650 33070 15652 33122
rect 15596 33068 15652 33070
rect 14924 31778 14980 31780
rect 14924 31726 14926 31778
rect 14926 31726 14978 31778
rect 14978 31726 14980 31778
rect 14924 31724 14980 31726
rect 14812 31666 14868 31668
rect 14812 31614 14814 31666
rect 14814 31614 14866 31666
rect 14866 31614 14868 31666
rect 14812 31612 14868 31614
rect 14700 31554 14756 31556
rect 14700 31502 14702 31554
rect 14702 31502 14754 31554
rect 14754 31502 14756 31554
rect 14700 31500 14756 31502
rect 18620 39730 18676 39732
rect 18620 39678 18622 39730
rect 18622 39678 18674 39730
rect 18674 39678 18676 39730
rect 18620 39676 18676 39678
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 16716 37436 16772 37492
rect 16828 38332 16884 38388
rect 17164 38220 17220 38276
rect 17388 38108 17444 38164
rect 18172 38834 18228 38836
rect 18172 38782 18174 38834
rect 18174 38782 18226 38834
rect 18226 38782 18228 38834
rect 18172 38780 18228 38782
rect 21308 38892 21364 38948
rect 18396 38780 18452 38836
rect 17836 38220 17892 38276
rect 16828 37548 16884 37604
rect 16604 35868 16660 35924
rect 16604 33852 16660 33908
rect 17388 37772 17444 37828
rect 18172 37884 18228 37940
rect 17500 37490 17556 37492
rect 17500 37438 17502 37490
rect 17502 37438 17554 37490
rect 17554 37438 17556 37490
rect 17500 37436 17556 37438
rect 17612 37378 17668 37380
rect 17612 37326 17614 37378
rect 17614 37326 17666 37378
rect 17666 37326 17668 37378
rect 17612 37324 17668 37326
rect 18060 37212 18116 37268
rect 17500 35308 17556 35364
rect 17276 34914 17332 34916
rect 17276 34862 17278 34914
rect 17278 34862 17330 34914
rect 17330 34862 17332 34914
rect 17276 34860 17332 34862
rect 17948 34914 18004 34916
rect 17948 34862 17950 34914
rect 17950 34862 18002 34914
rect 18002 34862 18004 34914
rect 17948 34860 18004 34862
rect 17612 34636 17668 34692
rect 15372 31164 15428 31220
rect 14924 30268 14980 30324
rect 14588 28924 14644 28980
rect 14700 28588 14756 28644
rect 13804 28476 13860 28532
rect 12796 24050 12852 24052
rect 12796 23998 12798 24050
rect 12798 23998 12850 24050
rect 12850 23998 12852 24050
rect 12796 23996 12852 23998
rect 11900 23938 11956 23940
rect 11900 23886 11902 23938
rect 11902 23886 11954 23938
rect 11954 23886 11956 23938
rect 11900 23884 11956 23886
rect 14028 25564 14084 25620
rect 14252 26908 14308 26964
rect 13804 23996 13860 24052
rect 12908 23714 12964 23716
rect 12908 23662 12910 23714
rect 12910 23662 12962 23714
rect 12962 23662 12964 23714
rect 12908 23660 12964 23662
rect 11564 22876 11620 22932
rect 11340 21756 11396 21812
rect 11452 21980 11508 22036
rect 10780 20130 10836 20132
rect 10780 20078 10782 20130
rect 10782 20078 10834 20130
rect 10834 20078 10836 20130
rect 10780 20076 10836 20078
rect 11116 19234 11172 19236
rect 11116 19182 11118 19234
rect 11118 19182 11170 19234
rect 11170 19182 11172 19234
rect 11116 19180 11172 19182
rect 9884 16604 9940 16660
rect 9772 16156 9828 16212
rect 8988 15426 9044 15428
rect 8988 15374 8990 15426
rect 8990 15374 9042 15426
rect 9042 15374 9044 15426
rect 8988 15372 9044 15374
rect 9212 15260 9268 15316
rect 10332 16828 10388 16884
rect 10444 17052 10500 17108
rect 11340 20076 11396 20132
rect 10892 16658 10948 16660
rect 10892 16606 10894 16658
rect 10894 16606 10946 16658
rect 10946 16606 10948 16658
rect 10892 16604 10948 16606
rect 10444 16210 10500 16212
rect 10444 16158 10446 16210
rect 10446 16158 10498 16210
rect 10498 16158 10500 16210
rect 10444 16156 10500 16158
rect 10220 15484 10276 15540
rect 7308 14476 7364 14532
rect 7196 13468 7252 13524
rect 10108 15202 10164 15204
rect 10108 15150 10110 15202
rect 10110 15150 10162 15202
rect 10162 15150 10164 15202
rect 10108 15148 10164 15150
rect 8204 13916 8260 13972
rect 8092 13468 8148 13524
rect 9660 13970 9716 13972
rect 9660 13918 9662 13970
rect 9662 13918 9714 13970
rect 9714 13918 9716 13970
rect 9660 13916 9716 13918
rect 9548 13468 9604 13524
rect 8204 12124 8260 12180
rect 7084 11116 7140 11172
rect 7308 10834 7364 10836
rect 7308 10782 7310 10834
rect 7310 10782 7362 10834
rect 7362 10782 7364 10834
rect 7308 10780 7364 10782
rect 7420 10498 7476 10500
rect 7420 10446 7422 10498
rect 7422 10446 7474 10498
rect 7474 10446 7476 10498
rect 7420 10444 7476 10446
rect 8092 11116 8148 11172
rect 7532 9996 7588 10052
rect 8316 10444 8372 10500
rect 6972 8764 7028 8820
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4956 6412 5012 6468
rect 5292 6412 5348 6468
rect 5404 6748 5460 6804
rect 6300 6636 6356 6692
rect 5628 6524 5684 6580
rect 4956 5852 5012 5908
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4732 5234 4788 5236
rect 4732 5182 4734 5234
rect 4734 5182 4786 5234
rect 4786 5182 4788 5234
rect 4732 5180 4788 5182
rect 2604 5010 2660 5012
rect 2604 4958 2606 5010
rect 2606 4958 2658 5010
rect 2658 4958 2660 5010
rect 2604 4956 2660 4958
rect 3948 4562 4004 4564
rect 3948 4510 3950 4562
rect 3950 4510 4002 4562
rect 4002 4510 4004 4562
rect 3948 4508 4004 4510
rect 5740 6018 5796 6020
rect 5740 5966 5742 6018
rect 5742 5966 5794 6018
rect 5794 5966 5796 6018
rect 5740 5964 5796 5966
rect 6076 5906 6132 5908
rect 6076 5854 6078 5906
rect 6078 5854 6130 5906
rect 6130 5854 6132 5906
rect 6076 5852 6132 5854
rect 5852 5740 5908 5796
rect 5516 5180 5572 5236
rect 5628 5516 5684 5572
rect 6076 5628 6132 5684
rect 5964 4956 6020 5012
rect 4732 4338 4788 4340
rect 4732 4286 4734 4338
rect 4734 4286 4786 4338
rect 4786 4286 4788 4338
rect 4732 4284 4788 4286
rect 5516 4284 5572 4340
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 5068 3554 5124 3556
rect 5068 3502 5070 3554
rect 5070 3502 5122 3554
rect 5122 3502 5124 3554
rect 5068 3500 5124 3502
rect 5740 3554 5796 3556
rect 5740 3502 5742 3554
rect 5742 3502 5794 3554
rect 5794 3502 5796 3554
rect 5740 3500 5796 3502
rect 7196 6860 7252 6916
rect 6860 6802 6916 6804
rect 6860 6750 6862 6802
rect 6862 6750 6914 6802
rect 6914 6750 6916 6802
rect 6860 6748 6916 6750
rect 6748 6524 6804 6580
rect 7756 6578 7812 6580
rect 7756 6526 7758 6578
rect 7758 6526 7810 6578
rect 7810 6526 7812 6578
rect 7756 6524 7812 6526
rect 8876 12178 8932 12180
rect 8876 12126 8878 12178
rect 8878 12126 8930 12178
rect 8930 12126 8932 12178
rect 8876 12124 8932 12126
rect 8652 9996 8708 10052
rect 8652 9212 8708 9268
rect 9212 9436 9268 9492
rect 8876 8764 8932 8820
rect 8428 8316 8484 8372
rect 8092 7586 8148 7588
rect 8092 7534 8094 7586
rect 8094 7534 8146 7586
rect 8146 7534 8148 7586
rect 8092 7532 8148 7534
rect 7980 6748 8036 6804
rect 8092 6636 8148 6692
rect 8876 7980 8932 8036
rect 8428 6860 8484 6916
rect 8652 7532 8708 7588
rect 8652 6860 8708 6916
rect 10332 15426 10388 15428
rect 10332 15374 10334 15426
rect 10334 15374 10386 15426
rect 10386 15374 10388 15426
rect 10332 15372 10388 15374
rect 12460 22316 12516 22372
rect 12796 22204 12852 22260
rect 12684 21532 12740 21588
rect 11564 19964 11620 20020
rect 11676 20076 11732 20132
rect 11788 17948 11844 18004
rect 11676 17836 11732 17892
rect 11676 17106 11732 17108
rect 11676 17054 11678 17106
rect 11678 17054 11730 17106
rect 11730 17054 11732 17106
rect 11676 17052 11732 17054
rect 11788 16156 11844 16212
rect 10668 13468 10724 13524
rect 11116 12850 11172 12852
rect 11116 12798 11118 12850
rect 11118 12798 11170 12850
rect 11170 12798 11172 12850
rect 11116 12796 11172 12798
rect 9996 11228 10052 11284
rect 9996 9548 10052 9604
rect 9660 9266 9716 9268
rect 9660 9214 9662 9266
rect 9662 9214 9714 9266
rect 9714 9214 9716 9266
rect 9660 9212 9716 9214
rect 9436 9042 9492 9044
rect 9436 8990 9438 9042
rect 9438 8990 9490 9042
rect 9490 8990 9492 9042
rect 9436 8988 9492 8990
rect 9324 8316 9380 8372
rect 9884 8092 9940 8148
rect 9660 7698 9716 7700
rect 9660 7646 9662 7698
rect 9662 7646 9714 7698
rect 9714 7646 9716 7698
rect 9660 7644 9716 7646
rect 11788 15148 11844 15204
rect 11676 14306 11732 14308
rect 11676 14254 11678 14306
rect 11678 14254 11730 14306
rect 11730 14254 11732 14306
rect 11676 14252 11732 14254
rect 11452 13468 11508 13524
rect 13916 23714 13972 23716
rect 13916 23662 13918 23714
rect 13918 23662 13970 23714
rect 13970 23662 13972 23714
rect 13916 23660 13972 23662
rect 14028 23212 14084 23268
rect 14028 22594 14084 22596
rect 14028 22542 14030 22594
rect 14030 22542 14082 22594
rect 14082 22542 14084 22594
rect 14028 22540 14084 22542
rect 13356 22204 13412 22260
rect 13468 21586 13524 21588
rect 13468 21534 13470 21586
rect 13470 21534 13522 21586
rect 13522 21534 13524 21586
rect 13468 21532 13524 21534
rect 14140 22092 14196 22148
rect 15372 28476 15428 28532
rect 14812 26962 14868 26964
rect 14812 26910 14814 26962
rect 14814 26910 14866 26962
rect 14866 26910 14868 26962
rect 14812 26908 14868 26910
rect 14812 22876 14868 22932
rect 14588 22258 14644 22260
rect 14588 22206 14590 22258
rect 14590 22206 14642 22258
rect 14642 22206 14644 22258
rect 14588 22204 14644 22206
rect 14700 22092 14756 22148
rect 14364 21756 14420 21812
rect 14476 21644 14532 21700
rect 14588 21586 14644 21588
rect 14588 21534 14590 21586
rect 14590 21534 14642 21586
rect 14642 21534 14644 21586
rect 14588 21532 14644 21534
rect 12908 20748 12964 20804
rect 12460 19906 12516 19908
rect 12460 19854 12462 19906
rect 12462 19854 12514 19906
rect 12514 19854 12516 19906
rect 12460 19852 12516 19854
rect 13804 20076 13860 20132
rect 13356 20018 13412 20020
rect 13356 19966 13358 20018
rect 13358 19966 13410 20018
rect 13410 19966 13412 20018
rect 13356 19964 13412 19966
rect 13692 19852 13748 19908
rect 13580 19292 13636 19348
rect 12796 18396 12852 18452
rect 12236 16716 12292 16772
rect 12572 16604 12628 16660
rect 12684 15820 12740 15876
rect 11900 14924 11956 14980
rect 13580 14812 13636 14868
rect 12348 13916 12404 13972
rect 12012 13746 12068 13748
rect 12012 13694 12014 13746
rect 12014 13694 12066 13746
rect 12066 13694 12068 13746
rect 12012 13692 12068 13694
rect 13468 14306 13524 14308
rect 13468 14254 13470 14306
rect 13470 14254 13522 14306
rect 13522 14254 13524 14306
rect 13468 14252 13524 14254
rect 11452 11564 11508 11620
rect 12236 11564 12292 11620
rect 11564 11282 11620 11284
rect 11564 11230 11566 11282
rect 11566 11230 11618 11282
rect 11618 11230 11620 11282
rect 11564 11228 11620 11230
rect 12460 11452 12516 11508
rect 13580 12796 13636 12852
rect 14028 21420 14084 21476
rect 14924 21196 14980 21252
rect 15372 27356 15428 27412
rect 15148 23884 15204 23940
rect 15260 22428 15316 22484
rect 15148 21084 15204 21140
rect 14924 20076 14980 20132
rect 15148 20130 15204 20132
rect 15148 20078 15150 20130
rect 15150 20078 15202 20130
rect 15202 20078 15204 20130
rect 15148 20076 15204 20078
rect 16156 31666 16212 31668
rect 16156 31614 16158 31666
rect 16158 31614 16210 31666
rect 16210 31614 16212 31666
rect 16156 31612 16212 31614
rect 16268 31554 16324 31556
rect 16268 31502 16270 31554
rect 16270 31502 16322 31554
rect 16322 31502 16324 31554
rect 16268 31500 16324 31502
rect 16604 31052 16660 31108
rect 17388 33458 17444 33460
rect 17388 33406 17390 33458
rect 17390 33406 17442 33458
rect 17442 33406 17444 33458
rect 17388 33404 17444 33406
rect 17276 33180 17332 33236
rect 18284 37100 18340 37156
rect 19292 38108 19348 38164
rect 18396 36876 18452 36932
rect 18956 37938 19012 37940
rect 18956 37886 18958 37938
rect 18958 37886 19010 37938
rect 19010 37886 19012 37938
rect 18956 37884 19012 37886
rect 20300 38780 20356 38836
rect 20076 38332 20132 38388
rect 18732 37772 18788 37828
rect 19628 37826 19684 37828
rect 19628 37774 19630 37826
rect 19630 37774 19682 37826
rect 19682 37774 19684 37826
rect 19628 37772 19684 37774
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19068 37154 19124 37156
rect 19068 37102 19070 37154
rect 19070 37102 19122 37154
rect 19122 37102 19124 37154
rect 19068 37100 19124 37102
rect 20972 38834 21028 38836
rect 20972 38782 20974 38834
rect 20974 38782 21026 38834
rect 21026 38782 21028 38834
rect 20972 38780 21028 38782
rect 20860 38444 20916 38500
rect 21644 38444 21700 38500
rect 20524 37826 20580 37828
rect 20524 37774 20526 37826
rect 20526 37774 20578 37826
rect 20578 37774 20580 37826
rect 20524 37772 20580 37774
rect 20412 37154 20468 37156
rect 20412 37102 20414 37154
rect 20414 37102 20466 37154
rect 20466 37102 20468 37154
rect 20412 37100 20468 37102
rect 20524 36876 20580 36932
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 18396 35308 18452 35364
rect 17836 33852 17892 33908
rect 17388 31836 17444 31892
rect 17724 32172 17780 32228
rect 17276 31554 17332 31556
rect 17276 31502 17278 31554
rect 17278 31502 17330 31554
rect 17330 31502 17332 31554
rect 17276 31500 17332 31502
rect 17500 31554 17556 31556
rect 17500 31502 17502 31554
rect 17502 31502 17554 31554
rect 17554 31502 17556 31554
rect 17500 31500 17556 31502
rect 17388 31106 17444 31108
rect 17388 31054 17390 31106
rect 17390 31054 17442 31106
rect 17442 31054 17444 31106
rect 17388 31052 17444 31054
rect 17164 29986 17220 29988
rect 17164 29934 17166 29986
rect 17166 29934 17218 29986
rect 17218 29934 17220 29986
rect 17164 29932 17220 29934
rect 16716 29820 16772 29876
rect 17948 31836 18004 31892
rect 18060 31666 18116 31668
rect 18060 31614 18062 31666
rect 18062 31614 18114 31666
rect 18114 31614 18116 31666
rect 18060 31612 18116 31614
rect 18284 33964 18340 34020
rect 18284 33180 18340 33236
rect 18620 34412 18676 34468
rect 19852 35644 19908 35700
rect 21196 35532 21252 35588
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 18732 33292 18788 33348
rect 17612 30268 17668 30324
rect 16716 27356 16772 27412
rect 15484 26124 15540 26180
rect 15596 25618 15652 25620
rect 15596 25566 15598 25618
rect 15598 25566 15650 25618
rect 15650 25566 15652 25618
rect 15596 25564 15652 25566
rect 16268 25228 16324 25284
rect 16828 25282 16884 25284
rect 16828 25230 16830 25282
rect 16830 25230 16882 25282
rect 16882 25230 16884 25282
rect 16828 25228 16884 25230
rect 17052 23324 17108 23380
rect 15596 23212 15652 23268
rect 15932 22764 15988 22820
rect 16828 22876 16884 22932
rect 16156 22428 16212 22484
rect 16940 22482 16996 22484
rect 16940 22430 16942 22482
rect 16942 22430 16994 22482
rect 16994 22430 16996 22482
rect 16940 22428 16996 22430
rect 15708 22370 15764 22372
rect 15708 22318 15710 22370
rect 15710 22318 15762 22370
rect 15762 22318 15764 22370
rect 15708 22316 15764 22318
rect 16044 22370 16100 22372
rect 16044 22318 16046 22370
rect 16046 22318 16098 22370
rect 16098 22318 16100 22370
rect 16044 22316 16100 22318
rect 15596 22258 15652 22260
rect 15596 22206 15598 22258
rect 15598 22206 15650 22258
rect 15650 22206 15652 22258
rect 15596 22204 15652 22206
rect 15596 21474 15652 21476
rect 15596 21422 15598 21474
rect 15598 21422 15650 21474
rect 15650 21422 15652 21474
rect 15596 21420 15652 21422
rect 13804 12124 13860 12180
rect 13692 11506 13748 11508
rect 13692 11454 13694 11506
rect 13694 11454 13746 11506
rect 13746 11454 13748 11506
rect 13692 11452 13748 11454
rect 12348 11170 12404 11172
rect 12348 11118 12350 11170
rect 12350 11118 12402 11170
rect 12402 11118 12404 11170
rect 12348 11116 12404 11118
rect 11788 8930 11844 8932
rect 11788 8878 11790 8930
rect 11790 8878 11842 8930
rect 11842 8878 11844 8930
rect 11788 8876 11844 8878
rect 11340 8540 11396 8596
rect 12124 8428 12180 8484
rect 11676 8204 11732 8260
rect 10556 8092 10612 8148
rect 11228 7868 11284 7924
rect 9772 7586 9828 7588
rect 9772 7534 9774 7586
rect 9774 7534 9826 7586
rect 9826 7534 9828 7586
rect 9772 7532 9828 7534
rect 10668 7586 10724 7588
rect 10668 7534 10670 7586
rect 10670 7534 10722 7586
rect 10722 7534 10724 7586
rect 10668 7532 10724 7534
rect 10220 7474 10276 7476
rect 10220 7422 10222 7474
rect 10222 7422 10274 7474
rect 10274 7422 10276 7474
rect 10220 7420 10276 7422
rect 10668 6748 10724 6804
rect 8764 6524 8820 6580
rect 7644 5964 7700 6020
rect 7308 5740 7364 5796
rect 7084 5682 7140 5684
rect 7084 5630 7086 5682
rect 7086 5630 7138 5682
rect 7138 5630 7140 5682
rect 7084 5628 7140 5630
rect 8092 5516 8148 5572
rect 8652 5292 8708 5348
rect 8876 6466 8932 6468
rect 8876 6414 8878 6466
rect 8878 6414 8930 6466
rect 8930 6414 8932 6466
rect 8876 6412 8932 6414
rect 7756 5234 7812 5236
rect 7756 5182 7758 5234
rect 7758 5182 7810 5234
rect 7810 5182 7812 5234
rect 7756 5180 7812 5182
rect 8540 5122 8596 5124
rect 8540 5070 8542 5122
rect 8542 5070 8594 5122
rect 8594 5070 8596 5122
rect 8540 5068 8596 5070
rect 7756 3666 7812 3668
rect 7756 3614 7758 3666
rect 7758 3614 7810 3666
rect 7810 3614 7812 3666
rect 7756 3612 7812 3614
rect 8540 3612 8596 3668
rect 8988 5234 9044 5236
rect 8988 5182 8990 5234
rect 8990 5182 9042 5234
rect 9042 5182 9044 5234
rect 8988 5180 9044 5182
rect 9548 6412 9604 6468
rect 9212 5180 9268 5236
rect 9660 5964 9716 6020
rect 11004 6860 11060 6916
rect 10892 6076 10948 6132
rect 10332 5906 10388 5908
rect 10332 5854 10334 5906
rect 10334 5854 10386 5906
rect 10386 5854 10388 5906
rect 10332 5852 10388 5854
rect 11676 6860 11732 6916
rect 11452 6748 11508 6804
rect 12012 6076 12068 6132
rect 11788 6018 11844 6020
rect 11788 5966 11790 6018
rect 11790 5966 11842 6018
rect 11842 5966 11844 6018
rect 11788 5964 11844 5966
rect 10556 5740 10612 5796
rect 9548 5122 9604 5124
rect 9548 5070 9550 5122
rect 9550 5070 9602 5122
rect 9602 5070 9604 5122
rect 9548 5068 9604 5070
rect 9660 5180 9716 5236
rect 10556 4508 10612 4564
rect 13244 10108 13300 10164
rect 13244 9548 13300 9604
rect 12460 8540 12516 8596
rect 12236 8092 12292 8148
rect 12684 8316 12740 8372
rect 13692 8204 13748 8260
rect 13804 9660 13860 9716
rect 13580 7980 13636 8036
rect 13692 7420 13748 7476
rect 12908 6748 12964 6804
rect 13468 6636 13524 6692
rect 12684 6466 12740 6468
rect 12684 6414 12686 6466
rect 12686 6414 12738 6466
rect 12738 6414 12740 6466
rect 12684 6412 12740 6414
rect 12460 5964 12516 6020
rect 13132 6076 13188 6132
rect 12908 5794 12964 5796
rect 12908 5742 12910 5794
rect 12910 5742 12962 5794
rect 12962 5742 12964 5794
rect 12908 5740 12964 5742
rect 12796 5346 12852 5348
rect 12796 5294 12798 5346
rect 12798 5294 12850 5346
rect 12850 5294 12852 5346
rect 12796 5292 12852 5294
rect 13916 8258 13972 8260
rect 13916 8206 13918 8258
rect 13918 8206 13970 8258
rect 13970 8206 13972 8258
rect 13916 8204 13972 8206
rect 13692 6860 13748 6916
rect 13916 6130 13972 6132
rect 13916 6078 13918 6130
rect 13918 6078 13970 6130
rect 13970 6078 13972 6130
rect 13916 6076 13972 6078
rect 13804 4284 13860 4340
rect 12124 3612 12180 3668
rect 13132 3612 13188 3668
rect 14812 19404 14868 19460
rect 14588 19346 14644 19348
rect 14588 19294 14590 19346
rect 14590 19294 14642 19346
rect 14642 19294 14644 19346
rect 14588 19292 14644 19294
rect 14812 18172 14868 18228
rect 14364 16156 14420 16212
rect 14588 15986 14644 15988
rect 14588 15934 14590 15986
rect 14590 15934 14642 15986
rect 14642 15934 14644 15986
rect 14588 15932 14644 15934
rect 14924 15874 14980 15876
rect 14924 15822 14926 15874
rect 14926 15822 14978 15874
rect 14978 15822 14980 15874
rect 14924 15820 14980 15822
rect 14140 8876 14196 8932
rect 14140 6524 14196 6580
rect 14140 6300 14196 6356
rect 15260 16044 15316 16100
rect 15260 14812 15316 14868
rect 14588 14306 14644 14308
rect 14588 14254 14590 14306
rect 14590 14254 14642 14306
rect 14642 14254 14644 14306
rect 14588 14252 14644 14254
rect 15148 13916 15204 13972
rect 15036 13634 15092 13636
rect 15036 13582 15038 13634
rect 15038 13582 15090 13634
rect 15090 13582 15092 13634
rect 15036 13580 15092 13582
rect 14700 11452 14756 11508
rect 15036 11116 15092 11172
rect 15484 19740 15540 19796
rect 15484 19010 15540 19012
rect 15484 18958 15486 19010
rect 15486 18958 15538 19010
rect 15538 18958 15540 19010
rect 15484 18956 15540 18958
rect 15932 20076 15988 20132
rect 16380 20130 16436 20132
rect 16380 20078 16382 20130
rect 16382 20078 16434 20130
rect 16434 20078 16436 20130
rect 16380 20076 16436 20078
rect 15932 19404 15988 19460
rect 17500 29820 17556 29876
rect 17724 30156 17780 30212
rect 17724 29932 17780 29988
rect 17276 29260 17332 29316
rect 16716 19964 16772 20020
rect 16716 18844 16772 18900
rect 16604 18060 16660 18116
rect 15708 16210 15764 16212
rect 15708 16158 15710 16210
rect 15710 16158 15762 16210
rect 15762 16158 15764 16210
rect 15708 16156 15764 16158
rect 15596 13580 15652 13636
rect 16156 15148 16212 15204
rect 15820 12348 15876 12404
rect 15372 9436 15428 9492
rect 15932 8316 15988 8372
rect 15260 8258 15316 8260
rect 15260 8206 15262 8258
rect 15262 8206 15314 8258
rect 15314 8206 15316 8258
rect 15260 8204 15316 8206
rect 16044 8204 16100 8260
rect 14700 8146 14756 8148
rect 14700 8094 14702 8146
rect 14702 8094 14754 8146
rect 14754 8094 14756 8146
rect 14700 8092 14756 8094
rect 15372 8146 15428 8148
rect 15372 8094 15374 8146
rect 15374 8094 15426 8146
rect 15426 8094 15428 8146
rect 15372 8092 15428 8094
rect 17052 20076 17108 20132
rect 17724 29538 17780 29540
rect 17724 29486 17726 29538
rect 17726 29486 17778 29538
rect 17778 29486 17780 29538
rect 17724 29484 17780 29486
rect 17612 29036 17668 29092
rect 18620 31612 18676 31668
rect 19180 33964 19236 34020
rect 19628 34130 19684 34132
rect 19628 34078 19630 34130
rect 19630 34078 19682 34130
rect 19682 34078 19684 34130
rect 19628 34076 19684 34078
rect 19628 33458 19684 33460
rect 19628 33406 19630 33458
rect 19630 33406 19682 33458
rect 19682 33406 19684 33458
rect 19628 33404 19684 33406
rect 19068 33346 19124 33348
rect 19068 33294 19070 33346
rect 19070 33294 19122 33346
rect 19122 33294 19124 33346
rect 19068 33292 19124 33294
rect 20972 34018 21028 34020
rect 20972 33966 20974 34018
rect 20974 33966 21026 34018
rect 21026 33966 21028 34018
rect 20972 33964 21028 33966
rect 20300 33404 20356 33460
rect 20188 33292 20244 33348
rect 19852 33180 19908 33236
rect 19516 33068 19572 33124
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19628 32786 19684 32788
rect 19628 32734 19630 32786
rect 19630 32734 19682 32786
rect 19682 32734 19684 32786
rect 19628 32732 19684 32734
rect 19516 32338 19572 32340
rect 19516 32286 19518 32338
rect 19518 32286 19570 32338
rect 19570 32286 19572 32338
rect 19516 32284 19572 32286
rect 20524 33346 20580 33348
rect 20524 33294 20526 33346
rect 20526 33294 20578 33346
rect 20578 33294 20580 33346
rect 20524 33292 20580 33294
rect 20636 33234 20692 33236
rect 20636 33182 20638 33234
rect 20638 33182 20690 33234
rect 20690 33182 20692 33234
rect 20636 33180 20692 33182
rect 18956 31554 19012 31556
rect 18956 31502 18958 31554
rect 18958 31502 19010 31554
rect 19010 31502 19012 31554
rect 18956 31500 19012 31502
rect 18620 30940 18676 30996
rect 18396 30268 18452 30324
rect 18060 29932 18116 29988
rect 18396 29986 18452 29988
rect 18396 29934 18398 29986
rect 18398 29934 18450 29986
rect 18450 29934 18452 29986
rect 18396 29932 18452 29934
rect 18620 30156 18676 30212
rect 18732 30098 18788 30100
rect 18732 30046 18734 30098
rect 18734 30046 18786 30098
rect 18786 30046 18788 30098
rect 18732 30044 18788 30046
rect 18172 29538 18228 29540
rect 18172 29486 18174 29538
rect 18174 29486 18226 29538
rect 18226 29486 18228 29538
rect 18172 29484 18228 29486
rect 17948 28028 18004 28084
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19180 31052 19236 31108
rect 20412 30156 20468 30212
rect 19068 29932 19124 29988
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19180 29538 19236 29540
rect 19180 29486 19182 29538
rect 19182 29486 19234 29538
rect 19234 29486 19236 29538
rect 19180 29484 19236 29486
rect 20188 28642 20244 28644
rect 20188 28590 20190 28642
rect 20190 28590 20242 28642
rect 20242 28590 20244 28642
rect 20188 28588 20244 28590
rect 20636 29426 20692 29428
rect 20636 29374 20638 29426
rect 20638 29374 20690 29426
rect 20690 29374 20692 29426
rect 20636 29372 20692 29374
rect 21868 37938 21924 37940
rect 21868 37886 21870 37938
rect 21870 37886 21922 37938
rect 21922 37886 21924 37938
rect 21868 37884 21924 37886
rect 21756 37826 21812 37828
rect 21756 37774 21758 37826
rect 21758 37774 21810 37826
rect 21810 37774 21812 37826
rect 21756 37772 21812 37774
rect 22876 38946 22932 38948
rect 22876 38894 22878 38946
rect 22878 38894 22930 38946
rect 22930 38894 22932 38946
rect 22876 38892 22932 38894
rect 22428 37772 22484 37828
rect 24108 37884 24164 37940
rect 23100 37826 23156 37828
rect 23100 37774 23102 37826
rect 23102 37774 23154 37826
rect 23154 37774 23156 37826
rect 23100 37772 23156 37774
rect 22652 37324 22708 37380
rect 21756 37100 21812 37156
rect 22204 36988 22260 37044
rect 22428 36876 22484 36932
rect 21420 35644 21476 35700
rect 22764 36428 22820 36484
rect 23436 36482 23492 36484
rect 23436 36430 23438 36482
rect 23438 36430 23490 36482
rect 23490 36430 23492 36482
rect 23436 36428 23492 36430
rect 22204 35698 22260 35700
rect 22204 35646 22206 35698
rect 22206 35646 22258 35698
rect 22258 35646 22260 35698
rect 22204 35644 22260 35646
rect 21868 35586 21924 35588
rect 21868 35534 21870 35586
rect 21870 35534 21922 35586
rect 21922 35534 21924 35586
rect 21868 35532 21924 35534
rect 23212 35586 23268 35588
rect 23212 35534 23214 35586
rect 23214 35534 23266 35586
rect 23266 35534 23268 35586
rect 23212 35532 23268 35534
rect 22876 35026 22932 35028
rect 22876 34974 22878 35026
rect 22878 34974 22930 35026
rect 22930 34974 22932 35026
rect 22876 34972 22932 34974
rect 21308 33852 21364 33908
rect 21644 33964 21700 34020
rect 21308 33292 21364 33348
rect 21756 33852 21812 33908
rect 21420 33122 21476 33124
rect 21420 33070 21422 33122
rect 21422 33070 21474 33122
rect 21474 33070 21476 33122
rect 21420 33068 21476 33070
rect 21308 32732 21364 32788
rect 21196 29260 21252 29316
rect 21308 28700 21364 28756
rect 20748 28642 20804 28644
rect 20748 28590 20750 28642
rect 20750 28590 20802 28642
rect 20802 28590 20804 28642
rect 20748 28588 20804 28590
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 22316 33068 22372 33124
rect 21644 32284 21700 32340
rect 22652 30268 22708 30324
rect 21756 28476 21812 28532
rect 22764 28754 22820 28756
rect 22764 28702 22766 28754
rect 22766 28702 22818 28754
rect 22818 28702 22820 28754
rect 22764 28700 22820 28702
rect 22652 28082 22708 28084
rect 22652 28030 22654 28082
rect 22654 28030 22706 28082
rect 22706 28030 22708 28082
rect 22652 28028 22708 28030
rect 21644 27970 21700 27972
rect 21644 27918 21646 27970
rect 21646 27918 21698 27970
rect 21698 27918 21700 27970
rect 21644 27916 21700 27918
rect 18284 26460 18340 26516
rect 17500 26178 17556 26180
rect 17500 26126 17502 26178
rect 17502 26126 17554 26178
rect 17554 26126 17556 26178
rect 17500 26124 17556 26126
rect 17500 25788 17556 25844
rect 17500 25282 17556 25284
rect 17500 25230 17502 25282
rect 17502 25230 17554 25282
rect 17554 25230 17556 25282
rect 17500 25228 17556 25230
rect 17948 25228 18004 25284
rect 18844 26124 18900 26180
rect 17500 23378 17556 23380
rect 17500 23326 17502 23378
rect 17502 23326 17554 23378
rect 17554 23326 17556 23378
rect 17500 23324 17556 23326
rect 18172 23324 18228 23380
rect 17612 23212 17668 23268
rect 17388 22764 17444 22820
rect 17388 20130 17444 20132
rect 17388 20078 17390 20130
rect 17390 20078 17442 20130
rect 17442 20078 17444 20130
rect 17388 20076 17444 20078
rect 17948 22930 18004 22932
rect 17948 22878 17950 22930
rect 17950 22878 18002 22930
rect 18002 22878 18004 22930
rect 17948 22876 18004 22878
rect 18508 23154 18564 23156
rect 18508 23102 18510 23154
rect 18510 23102 18562 23154
rect 18562 23102 18564 23154
rect 18508 23100 18564 23102
rect 18172 22428 18228 22484
rect 18396 22876 18452 22932
rect 18284 22370 18340 22372
rect 18284 22318 18286 22370
rect 18286 22318 18338 22370
rect 18338 22318 18340 22370
rect 18284 22316 18340 22318
rect 17276 17836 17332 17892
rect 17388 18508 17444 18564
rect 17388 16828 17444 16884
rect 17836 17052 17892 17108
rect 17836 16882 17892 16884
rect 17836 16830 17838 16882
rect 17838 16830 17890 16882
rect 17890 16830 17892 16882
rect 17836 16828 17892 16830
rect 17948 18396 18004 18452
rect 18396 19852 18452 19908
rect 18844 24722 18900 24724
rect 18844 24670 18846 24722
rect 18846 24670 18898 24722
rect 18898 24670 18900 24722
rect 18844 24668 18900 24670
rect 19292 24722 19348 24724
rect 19292 24670 19294 24722
rect 19294 24670 19346 24722
rect 19346 24670 19348 24722
rect 19292 24668 19348 24670
rect 18732 21980 18788 22036
rect 19516 23548 19572 23604
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 23884 20356 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19180 23100 19236 23156
rect 18956 22370 19012 22372
rect 18956 22318 18958 22370
rect 18958 22318 19010 22370
rect 19010 22318 19012 22370
rect 18956 22316 19012 22318
rect 19516 22988 19572 23044
rect 19068 22258 19124 22260
rect 19068 22206 19070 22258
rect 19070 22206 19122 22258
rect 19122 22206 19124 22258
rect 19068 22204 19124 22206
rect 18956 22146 19012 22148
rect 18956 22094 18958 22146
rect 18958 22094 19010 22146
rect 19010 22094 19012 22146
rect 18956 22092 19012 22094
rect 18284 18674 18340 18676
rect 18284 18622 18286 18674
rect 18286 18622 18338 18674
rect 18338 18622 18340 18674
rect 18284 18620 18340 18622
rect 19068 21586 19124 21588
rect 19068 21534 19070 21586
rect 19070 21534 19122 21586
rect 19122 21534 19124 21586
rect 19068 21532 19124 21534
rect 18732 21420 18788 21476
rect 18844 20524 18900 20580
rect 19068 20188 19124 20244
rect 18844 19292 18900 19348
rect 19292 19964 19348 20020
rect 19628 22204 19684 22260
rect 19964 22988 20020 23044
rect 20412 23042 20468 23044
rect 20412 22990 20414 23042
rect 20414 22990 20466 23042
rect 20466 22990 20468 23042
rect 20412 22988 20468 22990
rect 20412 22258 20468 22260
rect 20412 22206 20414 22258
rect 20414 22206 20466 22258
rect 20466 22206 20468 22258
rect 20412 22204 20468 22206
rect 19628 21980 19684 22036
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 21532 20132 21588
rect 19964 21420 20020 21476
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19628 19964 19684 20020
rect 19740 20188 19796 20244
rect 20524 20130 20580 20132
rect 20524 20078 20526 20130
rect 20526 20078 20578 20130
rect 20578 20078 20580 20130
rect 20524 20076 20580 20078
rect 19516 19180 19572 19236
rect 18956 18956 19012 19012
rect 18844 18620 18900 18676
rect 18508 18396 18564 18452
rect 20748 26178 20804 26180
rect 20748 26126 20750 26178
rect 20750 26126 20802 26178
rect 20802 26126 20804 26178
rect 20748 26124 20804 26126
rect 20748 25618 20804 25620
rect 20748 25566 20750 25618
rect 20750 25566 20802 25618
rect 20802 25566 20804 25618
rect 20748 25564 20804 25566
rect 21756 23938 21812 23940
rect 21756 23886 21758 23938
rect 21758 23886 21810 23938
rect 21810 23886 21812 23938
rect 21756 23884 21812 23886
rect 21644 23772 21700 23828
rect 20636 19628 20692 19684
rect 21196 19906 21252 19908
rect 21196 19854 21198 19906
rect 21198 19854 21250 19906
rect 21250 19854 21252 19906
rect 21196 19852 21252 19854
rect 19628 19122 19684 19124
rect 19628 19070 19630 19122
rect 19630 19070 19682 19122
rect 19682 19070 19684 19122
rect 19628 19068 19684 19070
rect 20076 19068 20132 19124
rect 20188 19010 20244 19012
rect 20188 18958 20190 19010
rect 20190 18958 20242 19010
rect 20242 18958 20244 19010
rect 20188 18956 20244 18958
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19852 18620 19908 18676
rect 19292 18396 19348 18452
rect 19628 18284 19684 18340
rect 18396 17724 18452 17780
rect 19068 18172 19124 18228
rect 18172 16882 18228 16884
rect 18172 16830 18174 16882
rect 18174 16830 18226 16882
rect 18226 16830 18228 16882
rect 18172 16828 18228 16830
rect 18732 17724 18788 17780
rect 18172 16380 18228 16436
rect 17836 15932 17892 15988
rect 17724 15820 17780 15876
rect 16268 14252 16324 14308
rect 16268 13692 16324 13748
rect 16156 7868 16212 7924
rect 14364 6636 14420 6692
rect 15820 6860 15876 6916
rect 15484 6748 15540 6804
rect 15372 6690 15428 6692
rect 15372 6638 15374 6690
rect 15374 6638 15426 6690
rect 15426 6638 15428 6690
rect 15372 6636 15428 6638
rect 15596 6690 15652 6692
rect 15596 6638 15598 6690
rect 15598 6638 15650 6690
rect 15650 6638 15652 6690
rect 15596 6636 15652 6638
rect 15372 6188 15428 6244
rect 15036 5964 15092 6020
rect 16940 9996 16996 10052
rect 16940 8988 16996 9044
rect 16492 8370 16548 8372
rect 16492 8318 16494 8370
rect 16494 8318 16546 8370
rect 16546 8318 16548 8370
rect 16492 8316 16548 8318
rect 17052 7644 17108 7700
rect 16156 6524 16212 6580
rect 16716 6860 16772 6916
rect 16940 6578 16996 6580
rect 16940 6526 16942 6578
rect 16942 6526 16994 6578
rect 16994 6526 16996 6578
rect 16940 6524 16996 6526
rect 16380 6412 16436 6468
rect 17612 14924 17668 14980
rect 17612 13970 17668 13972
rect 17612 13918 17614 13970
rect 17614 13918 17666 13970
rect 17666 13918 17668 13970
rect 17612 13916 17668 13918
rect 17948 14700 18004 14756
rect 17836 14140 17892 14196
rect 17948 13746 18004 13748
rect 17948 13694 17950 13746
rect 17950 13694 18002 13746
rect 18002 13694 18004 13746
rect 17948 13692 18004 13694
rect 17948 12908 18004 12964
rect 18172 16210 18228 16212
rect 18172 16158 18174 16210
rect 18174 16158 18226 16210
rect 18226 16158 18228 16210
rect 18172 16156 18228 16158
rect 18396 15708 18452 15764
rect 18508 16268 18564 16324
rect 18620 16156 18676 16212
rect 19740 18226 19796 18228
rect 19740 18174 19742 18226
rect 19742 18174 19794 18226
rect 19794 18174 19796 18226
rect 19740 18172 19796 18174
rect 19628 17666 19684 17668
rect 19628 17614 19630 17666
rect 19630 17614 19682 17666
rect 19682 17614 19684 17666
rect 19628 17612 19684 17614
rect 19740 17724 19796 17780
rect 18844 17106 18900 17108
rect 18844 17054 18846 17106
rect 18846 17054 18898 17106
rect 18898 17054 18900 17106
rect 18844 17052 18900 17054
rect 19292 16828 19348 16884
rect 19292 16268 19348 16324
rect 18508 15372 18564 15428
rect 18620 15596 18676 15652
rect 18396 15202 18452 15204
rect 18396 15150 18398 15202
rect 18398 15150 18450 15202
rect 18450 15150 18452 15202
rect 18396 15148 18452 15150
rect 18956 15932 19012 15988
rect 18284 14140 18340 14196
rect 18396 13970 18452 13972
rect 18396 13918 18398 13970
rect 18398 13918 18450 13970
rect 18450 13918 18452 13970
rect 18396 13916 18452 13918
rect 18620 14754 18676 14756
rect 18620 14702 18622 14754
rect 18622 14702 18674 14754
rect 18674 14702 18676 14754
rect 18620 14700 18676 14702
rect 18844 15090 18900 15092
rect 18844 15038 18846 15090
rect 18846 15038 18898 15090
rect 18898 15038 18900 15090
rect 18844 15036 18900 15038
rect 18732 14140 18788 14196
rect 18620 13580 18676 13636
rect 19068 15484 19124 15540
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19404 15820 19460 15876
rect 19404 15260 19460 15316
rect 19516 15202 19572 15204
rect 19516 15150 19518 15202
rect 19518 15150 19570 15202
rect 19570 15150 19572 15202
rect 19516 15148 19572 15150
rect 20748 16492 20804 16548
rect 19852 16268 19908 16324
rect 20188 16156 20244 16212
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20076 15538 20132 15540
rect 20076 15486 20078 15538
rect 20078 15486 20130 15538
rect 20130 15486 20132 15538
rect 20076 15484 20132 15486
rect 19740 15372 19796 15428
rect 20300 15314 20356 15316
rect 20300 15262 20302 15314
rect 20302 15262 20354 15314
rect 20354 15262 20356 15314
rect 20300 15260 20356 15262
rect 20748 15148 20804 15204
rect 24220 36204 24276 36260
rect 24444 37378 24500 37380
rect 24444 37326 24446 37378
rect 24446 37326 24498 37378
rect 24498 37326 24500 37378
rect 24444 37324 24500 37326
rect 24332 35756 24388 35812
rect 23996 34972 24052 35028
rect 23100 32732 23156 32788
rect 23212 31106 23268 31108
rect 23212 31054 23214 31106
rect 23214 31054 23266 31106
rect 23266 31054 23268 31106
rect 23212 31052 23268 31054
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 24668 37324 24724 37380
rect 28252 37324 28308 37380
rect 28812 37378 28868 37380
rect 28812 37326 28814 37378
rect 28814 37326 28866 37378
rect 28866 37326 28868 37378
rect 28812 37324 28868 37326
rect 24556 37154 24612 37156
rect 24556 37102 24558 37154
rect 24558 37102 24610 37154
rect 24610 37102 24612 37154
rect 24556 37100 24612 37102
rect 27580 37154 27636 37156
rect 27580 37102 27582 37154
rect 27582 37102 27634 37154
rect 27634 37102 27636 37154
rect 27580 37100 27636 37102
rect 25340 36988 25396 37044
rect 26236 36988 26292 37044
rect 24780 36370 24836 36372
rect 24780 36318 24782 36370
rect 24782 36318 24834 36370
rect 24834 36318 24836 36370
rect 24780 36316 24836 36318
rect 25564 36370 25620 36372
rect 25564 36318 25566 36370
rect 25566 36318 25618 36370
rect 25618 36318 25620 36370
rect 25564 36316 25620 36318
rect 24892 36204 24948 36260
rect 25004 35756 25060 35812
rect 24444 33068 24500 33124
rect 23548 32786 23604 32788
rect 23548 32734 23550 32786
rect 23550 32734 23602 32786
rect 23602 32734 23604 32786
rect 23548 32732 23604 32734
rect 25788 35756 25844 35812
rect 26684 35756 26740 35812
rect 25340 34972 25396 35028
rect 23660 32620 23716 32676
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 33068 36258 33124 36260
rect 33068 36206 33070 36258
rect 33070 36206 33122 36258
rect 33122 36206 33124 36258
rect 33068 36204 33124 36206
rect 33404 35756 33460 35812
rect 33740 36258 33796 36260
rect 33740 36206 33742 36258
rect 33742 36206 33794 36258
rect 33794 36206 33796 36258
rect 33740 36204 33796 36206
rect 28364 35026 28420 35028
rect 28364 34974 28366 35026
rect 28366 34974 28418 35026
rect 28418 34974 28420 35026
rect 28364 34972 28420 34974
rect 29148 34354 29204 34356
rect 29148 34302 29150 34354
rect 29150 34302 29202 34354
rect 29202 34302 29204 34354
rect 29148 34300 29204 34302
rect 25340 32732 25396 32788
rect 25452 33122 25508 33124
rect 25452 33070 25454 33122
rect 25454 33070 25506 33122
rect 25506 33070 25508 33122
rect 25452 33068 25508 33070
rect 25116 32620 25172 32676
rect 24108 30882 24164 30884
rect 24108 30830 24110 30882
rect 24110 30830 24162 30882
rect 24162 30830 24164 30882
rect 24108 30828 24164 30830
rect 23996 30322 24052 30324
rect 23996 30270 23998 30322
rect 23998 30270 24050 30322
rect 24050 30270 24052 30322
rect 23996 30268 24052 30270
rect 26012 31388 26068 31444
rect 26460 32562 26516 32564
rect 26460 32510 26462 32562
rect 26462 32510 26514 32562
rect 26514 32510 26516 32562
rect 26460 32508 26516 32510
rect 25004 30156 25060 30212
rect 25788 30604 25844 30660
rect 23548 29372 23604 29428
rect 22876 28140 22932 28196
rect 23100 27970 23156 27972
rect 23100 27918 23102 27970
rect 23102 27918 23154 27970
rect 23154 27918 23156 27970
rect 23100 27916 23156 27918
rect 22876 26178 22932 26180
rect 22876 26126 22878 26178
rect 22878 26126 22930 26178
rect 22930 26126 22932 26178
rect 22876 26124 22932 26126
rect 23996 29426 24052 29428
rect 23996 29374 23998 29426
rect 23998 29374 24050 29426
rect 24050 29374 24052 29426
rect 23996 29372 24052 29374
rect 23772 28530 23828 28532
rect 23772 28478 23774 28530
rect 23774 28478 23826 28530
rect 23826 28478 23828 28530
rect 23772 28476 23828 28478
rect 22428 24722 22484 24724
rect 22428 24670 22430 24722
rect 22430 24670 22482 24722
rect 22482 24670 22484 24722
rect 22428 24668 22484 24670
rect 22428 23826 22484 23828
rect 22428 23774 22430 23826
rect 22430 23774 22482 23826
rect 22482 23774 22484 23826
rect 22428 23772 22484 23774
rect 21980 23100 22036 23156
rect 21644 20300 21700 20356
rect 21644 19906 21700 19908
rect 21644 19854 21646 19906
rect 21646 19854 21698 19906
rect 21698 19854 21700 19906
rect 21644 19852 21700 19854
rect 21868 19906 21924 19908
rect 21868 19854 21870 19906
rect 21870 19854 21922 19906
rect 21922 19854 21924 19906
rect 21868 19852 21924 19854
rect 21308 19234 21364 19236
rect 21308 19182 21310 19234
rect 21310 19182 21362 19234
rect 21362 19182 21364 19234
rect 21308 19180 21364 19182
rect 21868 19404 21924 19460
rect 21644 19122 21700 19124
rect 21644 19070 21646 19122
rect 21646 19070 21698 19122
rect 21698 19070 21700 19122
rect 21644 19068 21700 19070
rect 21868 18732 21924 18788
rect 21532 18620 21588 18676
rect 22092 23042 22148 23044
rect 22092 22990 22094 23042
rect 22094 22990 22146 23042
rect 22146 22990 22148 23042
rect 22092 22988 22148 22990
rect 22540 22876 22596 22932
rect 23100 25788 23156 25844
rect 22764 23154 22820 23156
rect 22764 23102 22766 23154
rect 22766 23102 22818 23154
rect 22818 23102 22820 23154
rect 22764 23100 22820 23102
rect 22988 23154 23044 23156
rect 22988 23102 22990 23154
rect 22990 23102 23042 23154
rect 23042 23102 23044 23154
rect 22988 23100 23044 23102
rect 24668 24722 24724 24724
rect 24668 24670 24670 24722
rect 24670 24670 24722 24722
rect 24722 24670 24724 24722
rect 24668 24668 24724 24670
rect 24556 24108 24612 24164
rect 23548 23884 23604 23940
rect 23660 23324 23716 23380
rect 23436 23100 23492 23156
rect 23436 21980 23492 22036
rect 22876 20802 22932 20804
rect 22876 20750 22878 20802
rect 22878 20750 22930 20802
rect 22930 20750 22932 20802
rect 22876 20748 22932 20750
rect 22652 20076 22708 20132
rect 21868 17948 21924 18004
rect 22540 17666 22596 17668
rect 22540 17614 22542 17666
rect 22542 17614 22594 17666
rect 22594 17614 22596 17666
rect 22540 17612 22596 17614
rect 22540 16716 22596 16772
rect 22092 16380 22148 16436
rect 19516 14530 19572 14532
rect 19516 14478 19518 14530
rect 19518 14478 19570 14530
rect 19570 14478 19572 14530
rect 19516 14476 19572 14478
rect 19404 14140 19460 14196
rect 19180 13692 19236 13748
rect 18284 12402 18340 12404
rect 18284 12350 18286 12402
rect 18286 12350 18338 12402
rect 18338 12350 18340 12402
rect 18284 12348 18340 12350
rect 17612 11340 17668 11396
rect 17724 11788 17780 11844
rect 17836 11564 17892 11620
rect 18060 11340 18116 11396
rect 19068 12962 19124 12964
rect 19068 12910 19070 12962
rect 19070 12910 19122 12962
rect 19122 12910 19124 12962
rect 19068 12908 19124 12910
rect 18844 12348 18900 12404
rect 18956 12460 19012 12516
rect 19836 14138 19892 14140
rect 19628 14028 19684 14084
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19964 13970 20020 13972
rect 19964 13918 19966 13970
rect 19966 13918 20018 13970
rect 20018 13918 20020 13970
rect 19964 13916 20020 13918
rect 20300 13916 20356 13972
rect 20188 13580 20244 13636
rect 19516 12796 19572 12852
rect 19404 12402 19460 12404
rect 19404 12350 19406 12402
rect 19406 12350 19458 12402
rect 19458 12350 19460 12402
rect 19404 12348 19460 12350
rect 18620 11788 18676 11844
rect 19068 11900 19124 11956
rect 18844 11618 18900 11620
rect 18844 11566 18846 11618
rect 18846 11566 18898 11618
rect 18898 11566 18900 11618
rect 18844 11564 18900 11566
rect 19740 12738 19796 12740
rect 19740 12686 19742 12738
rect 19742 12686 19794 12738
rect 19794 12686 19796 12738
rect 19740 12684 19796 12686
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19516 11900 19572 11956
rect 18732 11452 18788 11508
rect 17948 11282 18004 11284
rect 17948 11230 17950 11282
rect 17950 11230 18002 11282
rect 18002 11230 18004 11282
rect 17948 11228 18004 11230
rect 18172 11004 18228 11060
rect 19068 11394 19124 11396
rect 19068 11342 19070 11394
rect 19070 11342 19122 11394
rect 19122 11342 19124 11394
rect 19068 11340 19124 11342
rect 17388 9436 17444 9492
rect 18396 9714 18452 9716
rect 18396 9662 18398 9714
rect 18398 9662 18450 9714
rect 18450 9662 18452 9714
rect 18396 9660 18452 9662
rect 18732 8316 18788 8372
rect 17724 7698 17780 7700
rect 17724 7646 17726 7698
rect 17726 7646 17778 7698
rect 17778 7646 17780 7698
rect 17724 7644 17780 7646
rect 19404 11452 19460 11508
rect 19964 11394 20020 11396
rect 19964 11342 19966 11394
rect 19966 11342 20018 11394
rect 20018 11342 20020 11394
rect 19964 11340 20020 11342
rect 20748 11394 20804 11396
rect 20748 11342 20750 11394
rect 20750 11342 20802 11394
rect 20802 11342 20804 11394
rect 20748 11340 20804 11342
rect 19404 10780 19460 10836
rect 19516 11004 19572 11060
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19740 10834 19796 10836
rect 19740 10782 19742 10834
rect 19742 10782 19794 10834
rect 19794 10782 19796 10834
rect 19740 10780 19796 10782
rect 20188 10834 20244 10836
rect 20188 10782 20190 10834
rect 20190 10782 20242 10834
rect 20242 10782 20244 10834
rect 20188 10780 20244 10782
rect 19628 10556 19684 10612
rect 20076 9660 20132 9716
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 21196 10610 21252 10612
rect 21196 10558 21198 10610
rect 21198 10558 21250 10610
rect 21250 10558 21252 10610
rect 21196 10556 21252 10558
rect 20748 8204 20804 8260
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 17948 7532 18004 7588
rect 17388 5906 17444 5908
rect 17388 5854 17390 5906
rect 17390 5854 17442 5906
rect 17442 5854 17444 5906
rect 17388 5852 17444 5854
rect 17836 6412 17892 6468
rect 16268 5794 16324 5796
rect 16268 5742 16270 5794
rect 16270 5742 16322 5794
rect 16322 5742 16324 5794
rect 16268 5740 16324 5742
rect 17612 5794 17668 5796
rect 17612 5742 17614 5794
rect 17614 5742 17666 5794
rect 17666 5742 17668 5794
rect 17612 5740 17668 5742
rect 16268 5234 16324 5236
rect 16268 5182 16270 5234
rect 16270 5182 16322 5234
rect 16322 5182 16324 5234
rect 16268 5180 16324 5182
rect 21420 13580 21476 13636
rect 21420 12402 21476 12404
rect 21420 12350 21422 12402
rect 21422 12350 21474 12402
rect 21474 12350 21476 12402
rect 21420 12348 21476 12350
rect 21980 12908 22036 12964
rect 21644 11282 21700 11284
rect 21644 11230 21646 11282
rect 21646 11230 21698 11282
rect 21698 11230 21700 11282
rect 21644 11228 21700 11230
rect 20972 7474 21028 7476
rect 20972 7422 20974 7474
rect 20974 7422 21026 7474
rect 21026 7422 21028 7474
rect 20972 7420 21028 7422
rect 21868 11394 21924 11396
rect 21868 11342 21870 11394
rect 21870 11342 21922 11394
rect 21922 11342 21924 11394
rect 21868 11340 21924 11342
rect 22540 16044 22596 16100
rect 22204 15932 22260 15988
rect 22428 15986 22484 15988
rect 22428 15934 22430 15986
rect 22430 15934 22482 15986
rect 22482 15934 22484 15986
rect 22428 15932 22484 15934
rect 22204 15484 22260 15540
rect 22876 17836 22932 17892
rect 22876 17106 22932 17108
rect 22876 17054 22878 17106
rect 22878 17054 22930 17106
rect 22930 17054 22932 17106
rect 22876 17052 22932 17054
rect 22876 15820 22932 15876
rect 23100 20018 23156 20020
rect 23100 19966 23102 20018
rect 23102 19966 23154 20018
rect 23154 19966 23156 20018
rect 23100 19964 23156 19966
rect 23884 23042 23940 23044
rect 23884 22990 23886 23042
rect 23886 22990 23938 23042
rect 23938 22990 23940 23042
rect 23884 22988 23940 22990
rect 23772 20076 23828 20132
rect 23996 19906 24052 19908
rect 23996 19854 23998 19906
rect 23998 19854 24050 19906
rect 24050 19854 24052 19906
rect 23996 19852 24052 19854
rect 24444 20018 24500 20020
rect 24444 19966 24446 20018
rect 24446 19966 24498 20018
rect 24498 19966 24500 20018
rect 24444 19964 24500 19966
rect 24220 19852 24276 19908
rect 23660 19404 23716 19460
rect 23212 18732 23268 18788
rect 23100 17612 23156 17668
rect 23212 17164 23268 17220
rect 23548 18508 23604 18564
rect 24556 18508 24612 18564
rect 23772 17836 23828 17892
rect 23436 17500 23492 17556
rect 23548 16994 23604 16996
rect 23548 16942 23550 16994
rect 23550 16942 23602 16994
rect 23602 16942 23604 16994
rect 23548 16940 23604 16942
rect 24332 17554 24388 17556
rect 24332 17502 24334 17554
rect 24334 17502 24386 17554
rect 24386 17502 24388 17554
rect 24332 17500 24388 17502
rect 24444 17442 24500 17444
rect 24444 17390 24446 17442
rect 24446 17390 24498 17442
rect 24498 17390 24500 17442
rect 24444 17388 24500 17390
rect 24108 16882 24164 16884
rect 24108 16830 24110 16882
rect 24110 16830 24162 16882
rect 24162 16830 24164 16882
rect 24108 16828 24164 16830
rect 23772 16044 23828 16100
rect 23324 15986 23380 15988
rect 23324 15934 23326 15986
rect 23326 15934 23378 15986
rect 23378 15934 23380 15986
rect 23324 15932 23380 15934
rect 23100 15820 23156 15876
rect 23436 15820 23492 15876
rect 23100 15538 23156 15540
rect 23100 15486 23102 15538
rect 23102 15486 23154 15538
rect 23154 15486 23156 15538
rect 23100 15484 23156 15486
rect 23996 15874 24052 15876
rect 23996 15822 23998 15874
rect 23998 15822 24050 15874
rect 24050 15822 24052 15874
rect 23996 15820 24052 15822
rect 23772 15484 23828 15540
rect 24556 16828 24612 16884
rect 25676 27020 25732 27076
rect 25228 26124 25284 26180
rect 25004 23938 25060 23940
rect 25004 23886 25006 23938
rect 25006 23886 25058 23938
rect 25058 23886 25060 23938
rect 25004 23884 25060 23886
rect 25452 25564 25508 25620
rect 25228 21308 25284 21364
rect 25228 20524 25284 20580
rect 25340 20188 25396 20244
rect 25564 24722 25620 24724
rect 25564 24670 25566 24722
rect 25566 24670 25618 24722
rect 25618 24670 25620 24722
rect 25564 24668 25620 24670
rect 25452 20300 25508 20356
rect 25564 24108 25620 24164
rect 25900 28588 25956 28644
rect 28252 33122 28308 33124
rect 28252 33070 28254 33122
rect 28254 33070 28306 33122
rect 28306 33070 28308 33122
rect 28252 33068 28308 33070
rect 28140 32562 28196 32564
rect 28140 32510 28142 32562
rect 28142 32510 28194 32562
rect 28194 32510 28196 32562
rect 28140 32508 28196 32510
rect 27468 30716 27524 30772
rect 27580 32396 27636 32452
rect 26236 29932 26292 29988
rect 26348 30156 26404 30212
rect 27468 30210 27524 30212
rect 27468 30158 27470 30210
rect 27470 30158 27522 30210
rect 27522 30158 27524 30210
rect 27468 30156 27524 30158
rect 26460 29932 26516 29988
rect 26796 29650 26852 29652
rect 26796 29598 26798 29650
rect 26798 29598 26850 29650
rect 26850 29598 26852 29650
rect 26796 29596 26852 29598
rect 26684 29538 26740 29540
rect 26684 29486 26686 29538
rect 26686 29486 26738 29538
rect 26738 29486 26740 29538
rect 26684 29484 26740 29486
rect 27356 30098 27412 30100
rect 27356 30046 27358 30098
rect 27358 30046 27410 30098
rect 27410 30046 27412 30098
rect 27356 30044 27412 30046
rect 27132 29932 27188 29988
rect 27020 29484 27076 29540
rect 26572 29372 26628 29428
rect 27132 29426 27188 29428
rect 27132 29374 27134 29426
rect 27134 29374 27186 29426
rect 27186 29374 27188 29426
rect 27132 29372 27188 29374
rect 26572 28588 26628 28644
rect 27356 29596 27412 29652
rect 25788 25506 25844 25508
rect 25788 25454 25790 25506
rect 25790 25454 25842 25506
rect 25842 25454 25844 25506
rect 25788 25452 25844 25454
rect 26908 28418 26964 28420
rect 26908 28366 26910 28418
rect 26910 28366 26962 28418
rect 26962 28366 26964 28418
rect 26908 28364 26964 28366
rect 26908 27858 26964 27860
rect 26908 27806 26910 27858
rect 26910 27806 26962 27858
rect 26962 27806 26964 27858
rect 26908 27804 26964 27806
rect 26236 27020 26292 27076
rect 26796 27074 26852 27076
rect 26796 27022 26798 27074
rect 26798 27022 26850 27074
rect 26850 27022 26852 27074
rect 26796 27020 26852 27022
rect 26572 26572 26628 26628
rect 26236 26236 26292 26292
rect 26012 24108 26068 24164
rect 26684 25900 26740 25956
rect 28588 31948 28644 32004
rect 28700 31164 28756 31220
rect 28476 31052 28532 31108
rect 27804 30940 27860 30996
rect 28252 30156 28308 30212
rect 27692 29932 27748 29988
rect 27580 29372 27636 29428
rect 28028 28588 28084 28644
rect 27468 28476 27524 28532
rect 27468 26572 27524 26628
rect 27020 26290 27076 26292
rect 27020 26238 27022 26290
rect 27022 26238 27074 26290
rect 27074 26238 27076 26290
rect 27020 26236 27076 26238
rect 26908 25788 26964 25844
rect 26236 24722 26292 24724
rect 26236 24670 26238 24722
rect 26238 24670 26290 24722
rect 26290 24670 26292 24722
rect 26236 24668 26292 24670
rect 27804 26572 27860 26628
rect 26908 23826 26964 23828
rect 26908 23774 26910 23826
rect 26910 23774 26962 23826
rect 26962 23774 26964 23826
rect 26908 23772 26964 23774
rect 27356 25116 27412 25172
rect 28140 28476 28196 28532
rect 28476 30044 28532 30100
rect 28476 29484 28532 29540
rect 28364 28642 28420 28644
rect 28364 28590 28366 28642
rect 28366 28590 28418 28642
rect 28418 28590 28420 28642
rect 28364 28588 28420 28590
rect 28700 28530 28756 28532
rect 28700 28478 28702 28530
rect 28702 28478 28754 28530
rect 28754 28478 28756 28530
rect 28700 28476 28756 28478
rect 28588 28418 28644 28420
rect 28588 28366 28590 28418
rect 28590 28366 28642 28418
rect 28642 28366 28644 28418
rect 28588 28364 28644 28366
rect 28252 27858 28308 27860
rect 28252 27806 28254 27858
rect 28254 27806 28306 27858
rect 28306 27806 28308 27858
rect 28252 27804 28308 27806
rect 28140 27132 28196 27188
rect 28252 26066 28308 26068
rect 28252 26014 28254 26066
rect 28254 26014 28306 26066
rect 28306 26014 28308 26066
rect 28252 26012 28308 26014
rect 28140 25004 28196 25060
rect 28252 25788 28308 25844
rect 29260 32732 29316 32788
rect 29484 32562 29540 32564
rect 29484 32510 29486 32562
rect 29486 32510 29538 32562
rect 29538 32510 29540 32562
rect 29484 32508 29540 32510
rect 29932 33964 29988 34020
rect 29820 33068 29876 33124
rect 30828 34242 30884 34244
rect 30828 34190 30830 34242
rect 30830 34190 30882 34242
rect 30882 34190 30884 34242
rect 30828 34188 30884 34190
rect 30380 32786 30436 32788
rect 30380 32734 30382 32786
rect 30382 32734 30434 32786
rect 30434 32734 30436 32786
rect 30380 32732 30436 32734
rect 30604 32732 30660 32788
rect 29596 32396 29652 32452
rect 30268 32396 30324 32452
rect 30492 32562 30548 32564
rect 30492 32510 30494 32562
rect 30494 32510 30546 32562
rect 30546 32510 30548 32562
rect 30492 32508 30548 32510
rect 29708 31218 29764 31220
rect 29708 31166 29710 31218
rect 29710 31166 29762 31218
rect 29762 31166 29764 31218
rect 29708 31164 29764 31166
rect 30268 30770 30324 30772
rect 30268 30718 30270 30770
rect 30270 30718 30322 30770
rect 30322 30718 30324 30770
rect 30268 30716 30324 30718
rect 30156 30268 30212 30324
rect 29148 27804 29204 27860
rect 29708 28530 29764 28532
rect 29708 28478 29710 28530
rect 29710 28478 29762 28530
rect 29762 28478 29764 28530
rect 29708 28476 29764 28478
rect 30380 30156 30436 30212
rect 30604 31724 30660 31780
rect 31052 33964 31108 34020
rect 31164 34972 31220 35028
rect 35084 35756 35140 35812
rect 31164 34076 31220 34132
rect 31724 34860 31780 34916
rect 32172 34242 32228 34244
rect 32172 34190 32174 34242
rect 32174 34190 32226 34242
rect 32226 34190 32228 34242
rect 32172 34188 32228 34190
rect 31276 34018 31332 34020
rect 31276 33966 31278 34018
rect 31278 33966 31330 34018
rect 31330 33966 31332 34018
rect 31276 33964 31332 33966
rect 31836 32562 31892 32564
rect 31836 32510 31838 32562
rect 31838 32510 31890 32562
rect 31890 32510 31892 32562
rect 31836 32508 31892 32510
rect 33180 33292 33236 33348
rect 32956 32786 33012 32788
rect 32956 32734 32958 32786
rect 32958 32734 33010 32786
rect 33010 32734 33012 32786
rect 32956 32732 33012 32734
rect 30828 32002 30884 32004
rect 30828 31950 30830 32002
rect 30830 31950 30882 32002
rect 30882 31950 30884 32002
rect 30828 31948 30884 31950
rect 31388 32060 31444 32116
rect 32284 32396 32340 32452
rect 30940 31724 30996 31780
rect 31276 31724 31332 31780
rect 31724 31724 31780 31780
rect 30940 31276 30996 31332
rect 31948 31778 32004 31780
rect 31948 31726 31950 31778
rect 31950 31726 32002 31778
rect 32002 31726 32004 31778
rect 31948 31724 32004 31726
rect 31836 31164 31892 31220
rect 31836 30994 31892 30996
rect 31836 30942 31838 30994
rect 31838 30942 31890 30994
rect 31890 30942 31892 30994
rect 31836 30940 31892 30942
rect 33292 32562 33348 32564
rect 33292 32510 33294 32562
rect 33294 32510 33346 32562
rect 33346 32510 33348 32562
rect 33292 32508 33348 32510
rect 34076 34130 34132 34132
rect 34076 34078 34078 34130
rect 34078 34078 34130 34130
rect 34130 34078 34132 34130
rect 34076 34076 34132 34078
rect 34076 33516 34132 33572
rect 34076 32508 34132 32564
rect 33180 32396 33236 32452
rect 32060 30994 32116 30996
rect 32060 30942 32062 30994
rect 32062 30942 32114 30994
rect 32114 30942 32116 30994
rect 32060 30940 32116 30942
rect 34076 31612 34132 31668
rect 33180 31218 33236 31220
rect 33180 31166 33182 31218
rect 33182 31166 33234 31218
rect 33234 31166 33236 31218
rect 33180 31164 33236 31166
rect 33404 30994 33460 30996
rect 33404 30942 33406 30994
rect 33406 30942 33458 30994
rect 33458 30942 33460 30994
rect 33404 30940 33460 30942
rect 31948 30604 32004 30660
rect 31164 30268 31220 30324
rect 31388 30210 31444 30212
rect 31388 30158 31390 30210
rect 31390 30158 31442 30210
rect 31442 30158 31444 30210
rect 31388 30156 31444 30158
rect 30044 28364 30100 28420
rect 31164 29538 31220 29540
rect 31164 29486 31166 29538
rect 31166 29486 31218 29538
rect 31218 29486 31220 29538
rect 31164 29484 31220 29486
rect 30492 28418 30548 28420
rect 30492 28366 30494 28418
rect 30494 28366 30546 28418
rect 30546 28366 30548 28418
rect 30492 28364 30548 28366
rect 30268 27916 30324 27972
rect 30044 27244 30100 27300
rect 29372 27186 29428 27188
rect 29372 27134 29374 27186
rect 29374 27134 29426 27186
rect 29426 27134 29428 27186
rect 29372 27132 29428 27134
rect 28924 25004 28980 25060
rect 28364 24834 28420 24836
rect 28364 24782 28366 24834
rect 28366 24782 28418 24834
rect 28418 24782 28420 24834
rect 28364 24780 28420 24782
rect 28588 24722 28644 24724
rect 28588 24670 28590 24722
rect 28590 24670 28642 24722
rect 28642 24670 28644 24722
rect 28588 24668 28644 24670
rect 29484 25788 29540 25844
rect 29148 25116 29204 25172
rect 29372 24834 29428 24836
rect 29372 24782 29374 24834
rect 29374 24782 29426 24834
rect 29426 24782 29428 24834
rect 29372 24780 29428 24782
rect 29708 24722 29764 24724
rect 29708 24670 29710 24722
rect 29710 24670 29762 24722
rect 29762 24670 29764 24722
rect 29708 24668 29764 24670
rect 27132 23772 27188 23828
rect 26908 23266 26964 23268
rect 26908 23214 26910 23266
rect 26910 23214 26962 23266
rect 26962 23214 26964 23266
rect 26908 23212 26964 23214
rect 25900 21586 25956 21588
rect 25900 21534 25902 21586
rect 25902 21534 25954 21586
rect 25954 21534 25956 21586
rect 25900 21532 25956 21534
rect 25676 21308 25732 21364
rect 26124 21084 26180 21140
rect 26012 20690 26068 20692
rect 26012 20638 26014 20690
rect 26014 20638 26066 20690
rect 26066 20638 26068 20690
rect 26012 20636 26068 20638
rect 25900 20300 25956 20356
rect 25228 19292 25284 19348
rect 24892 17052 24948 17108
rect 25228 16994 25284 16996
rect 25228 16942 25230 16994
rect 25230 16942 25282 16994
rect 25282 16942 25284 16994
rect 25228 16940 25284 16942
rect 24668 16268 24724 16324
rect 23884 15260 23940 15316
rect 23884 14476 23940 14532
rect 23772 14418 23828 14420
rect 23772 14366 23774 14418
rect 23774 14366 23826 14418
rect 23826 14366 23828 14418
rect 23772 14364 23828 14366
rect 22988 14252 23044 14308
rect 22316 12962 22372 12964
rect 22316 12910 22318 12962
rect 22318 12910 22370 12962
rect 22370 12910 22372 12962
rect 22316 12908 22372 12910
rect 22652 13634 22708 13636
rect 22652 13582 22654 13634
rect 22654 13582 22706 13634
rect 22706 13582 22708 13634
rect 22652 13580 22708 13582
rect 22876 13580 22932 13636
rect 22764 13522 22820 13524
rect 22764 13470 22766 13522
rect 22766 13470 22818 13522
rect 22818 13470 22820 13522
rect 22764 13468 22820 13470
rect 22764 12962 22820 12964
rect 22764 12910 22766 12962
rect 22766 12910 22818 12962
rect 22818 12910 22820 12962
rect 22764 12908 22820 12910
rect 22204 12178 22260 12180
rect 22204 12126 22206 12178
rect 22206 12126 22258 12178
rect 22258 12126 22260 12178
rect 22204 12124 22260 12126
rect 22204 11900 22260 11956
rect 22988 12850 23044 12852
rect 22988 12798 22990 12850
rect 22990 12798 23042 12850
rect 23042 12798 23044 12850
rect 22988 12796 23044 12798
rect 23884 13468 23940 13524
rect 23100 12460 23156 12516
rect 23436 12684 23492 12740
rect 22764 12124 22820 12180
rect 22092 11340 22148 11396
rect 21756 11116 21812 11172
rect 22092 11170 22148 11172
rect 22092 11118 22094 11170
rect 22094 11118 22146 11170
rect 22146 11118 22148 11170
rect 22092 11116 22148 11118
rect 22540 9660 22596 9716
rect 21084 6636 21140 6692
rect 19628 6524 19684 6580
rect 22092 7474 22148 7476
rect 22092 7422 22094 7474
rect 22094 7422 22146 7474
rect 22146 7422 22148 7474
rect 22092 7420 22148 7422
rect 23212 11452 23268 11508
rect 22988 11340 23044 11396
rect 24668 15260 24724 15316
rect 25228 14364 25284 14420
rect 24780 13692 24836 13748
rect 24780 12066 24836 12068
rect 24780 12014 24782 12066
rect 24782 12014 24834 12066
rect 24834 12014 24836 12066
rect 24780 12012 24836 12014
rect 24444 11900 24500 11956
rect 23436 11340 23492 11396
rect 23660 11282 23716 11284
rect 23660 11230 23662 11282
rect 23662 11230 23714 11282
rect 23714 11230 23716 11282
rect 23660 11228 23716 11230
rect 24108 11228 24164 11284
rect 22652 7644 22708 7700
rect 22876 10556 22932 10612
rect 23100 10444 23156 10500
rect 23996 10498 24052 10500
rect 23996 10446 23998 10498
rect 23998 10446 24050 10498
rect 24050 10446 24052 10498
rect 23996 10444 24052 10446
rect 24556 10610 24612 10612
rect 24556 10558 24558 10610
rect 24558 10558 24610 10610
rect 24610 10558 24612 10610
rect 24556 10556 24612 10558
rect 25452 19180 25508 19236
rect 26124 20076 26180 20132
rect 25564 16716 25620 16772
rect 26460 18284 26516 18340
rect 27020 21420 27076 21476
rect 26796 20802 26852 20804
rect 26796 20750 26798 20802
rect 26798 20750 26850 20802
rect 26850 20750 26852 20802
rect 26796 20748 26852 20750
rect 28476 23042 28532 23044
rect 28476 22990 28478 23042
rect 28478 22990 28530 23042
rect 28530 22990 28532 23042
rect 28476 22988 28532 22990
rect 27692 22876 27748 22932
rect 27692 21756 27748 21812
rect 28028 21196 28084 21252
rect 29932 23100 29988 23156
rect 29260 22370 29316 22372
rect 29260 22318 29262 22370
rect 29262 22318 29314 22370
rect 29314 22318 29316 22370
rect 29260 22316 29316 22318
rect 30044 22370 30100 22372
rect 30044 22318 30046 22370
rect 30046 22318 30098 22370
rect 30098 22318 30100 22370
rect 30044 22316 30100 22318
rect 28252 22146 28308 22148
rect 28252 22094 28254 22146
rect 28254 22094 28306 22146
rect 28306 22094 28308 22146
rect 28252 22092 28308 22094
rect 28140 21084 28196 21140
rect 28700 21980 28756 22036
rect 27580 20690 27636 20692
rect 27580 20638 27582 20690
rect 27582 20638 27634 20690
rect 27634 20638 27636 20690
rect 27580 20636 27636 20638
rect 27916 20524 27972 20580
rect 26908 20188 26964 20244
rect 27020 20130 27076 20132
rect 27020 20078 27022 20130
rect 27022 20078 27074 20130
rect 27074 20078 27076 20130
rect 27020 20076 27076 20078
rect 26684 20018 26740 20020
rect 26684 19966 26686 20018
rect 26686 19966 26738 20018
rect 26738 19966 26740 20018
rect 26684 19964 26740 19966
rect 26684 19180 26740 19236
rect 27244 18956 27300 19012
rect 27132 18732 27188 18788
rect 26796 18284 26852 18340
rect 26572 17836 26628 17892
rect 26796 16882 26852 16884
rect 26796 16830 26798 16882
rect 26798 16830 26850 16882
rect 26850 16830 26852 16882
rect 26796 16828 26852 16830
rect 26684 16098 26740 16100
rect 26684 16046 26686 16098
rect 26686 16046 26738 16098
rect 26738 16046 26740 16098
rect 26684 16044 26740 16046
rect 27692 19010 27748 19012
rect 27692 18958 27694 19010
rect 27694 18958 27746 19010
rect 27746 18958 27748 19010
rect 27692 18956 27748 18958
rect 27468 18620 27524 18676
rect 27468 17388 27524 17444
rect 27244 16492 27300 16548
rect 27244 15986 27300 15988
rect 27244 15934 27246 15986
rect 27246 15934 27298 15986
rect 27298 15934 27300 15986
rect 27244 15932 27300 15934
rect 27804 15986 27860 15988
rect 27804 15934 27806 15986
rect 27806 15934 27858 15986
rect 27858 15934 27860 15986
rect 27804 15932 27860 15934
rect 27356 15874 27412 15876
rect 27356 15822 27358 15874
rect 27358 15822 27410 15874
rect 27410 15822 27412 15874
rect 27356 15820 27412 15822
rect 27132 14476 27188 14532
rect 26012 14306 26068 14308
rect 26012 14254 26014 14306
rect 26014 14254 26066 14306
rect 26066 14254 26068 14306
rect 26012 14252 26068 14254
rect 25340 12796 25396 12852
rect 25564 12908 25620 12964
rect 25452 11788 25508 11844
rect 25788 11394 25844 11396
rect 25788 11342 25790 11394
rect 25790 11342 25842 11394
rect 25842 11342 25844 11394
rect 25788 11340 25844 11342
rect 26236 12962 26292 12964
rect 26236 12910 26238 12962
rect 26238 12910 26290 12962
rect 26290 12910 26292 12962
rect 26236 12908 26292 12910
rect 26012 12796 26068 12852
rect 26236 12460 26292 12516
rect 26012 12348 26068 12404
rect 26796 12684 26852 12740
rect 27132 12460 27188 12516
rect 28252 20690 28308 20692
rect 28252 20638 28254 20690
rect 28254 20638 28306 20690
rect 28306 20638 28308 20690
rect 28252 20636 28308 20638
rect 28140 20188 28196 20244
rect 28028 19964 28084 20020
rect 28588 20018 28644 20020
rect 28588 19966 28590 20018
rect 28590 19966 28642 20018
rect 28642 19966 28644 20018
rect 28588 19964 28644 19966
rect 28028 18956 28084 19012
rect 28028 15874 28084 15876
rect 28028 15822 28030 15874
rect 28030 15822 28082 15874
rect 28082 15822 28084 15874
rect 28028 15820 28084 15822
rect 29708 22092 29764 22148
rect 29372 21756 29428 21812
rect 29484 21868 29540 21924
rect 28700 14252 28756 14308
rect 27916 13580 27972 13636
rect 28140 12962 28196 12964
rect 28140 12910 28142 12962
rect 28142 12910 28194 12962
rect 28194 12910 28196 12962
rect 28140 12908 28196 12910
rect 28476 12908 28532 12964
rect 27804 12572 27860 12628
rect 27692 12348 27748 12404
rect 27468 12124 27524 12180
rect 26796 11900 26852 11956
rect 24892 10108 24948 10164
rect 26012 10108 26068 10164
rect 23548 9660 23604 9716
rect 24668 9042 24724 9044
rect 24668 8990 24670 9042
rect 24670 8990 24722 9042
rect 24722 8990 24724 9042
rect 24668 8988 24724 8990
rect 25340 9042 25396 9044
rect 25340 8990 25342 9042
rect 25342 8990 25394 9042
rect 25394 8990 25396 9042
rect 25340 8988 25396 8990
rect 26908 11900 26964 11956
rect 26460 11340 26516 11396
rect 26348 11116 26404 11172
rect 26572 11282 26628 11284
rect 26572 11230 26574 11282
rect 26574 11230 26626 11282
rect 26626 11230 26628 11282
rect 26572 11228 26628 11230
rect 26684 9884 26740 9940
rect 26124 8988 26180 9044
rect 25564 8092 25620 8148
rect 24444 7868 24500 7924
rect 22876 6690 22932 6692
rect 22876 6638 22878 6690
rect 22878 6638 22930 6690
rect 22930 6638 22932 6690
rect 22876 6636 22932 6638
rect 21756 6524 21812 6580
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19628 5852 19684 5908
rect 17948 5180 18004 5236
rect 16940 5122 16996 5124
rect 16940 5070 16942 5122
rect 16942 5070 16994 5122
rect 16994 5070 16996 5122
rect 16940 5068 16996 5070
rect 17612 5068 17668 5124
rect 16604 4396 16660 4452
rect 14924 4338 14980 4340
rect 14924 4286 14926 4338
rect 14926 4286 14978 4338
rect 14978 4286 14980 4338
rect 14924 4284 14980 4286
rect 14364 3500 14420 3556
rect 13916 3388 13972 3444
rect 14812 3388 14868 3444
rect 15260 3388 15316 3444
rect 17388 4450 17444 4452
rect 17388 4398 17390 4450
rect 17390 4398 17442 4450
rect 17442 4398 17444 4450
rect 17388 4396 17444 4398
rect 16940 3554 16996 3556
rect 16940 3502 16942 3554
rect 16942 3502 16994 3554
rect 16994 3502 16996 3554
rect 16940 3500 16996 3502
rect 21308 5292 21364 5348
rect 22876 6300 22932 6356
rect 21868 5906 21924 5908
rect 21868 5854 21870 5906
rect 21870 5854 21922 5906
rect 21922 5854 21924 5906
rect 21868 5852 21924 5854
rect 21756 5292 21812 5348
rect 22092 5292 22148 5348
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 23884 6636 23940 6692
rect 24220 6524 24276 6580
rect 24668 5964 24724 6020
rect 25340 6018 25396 6020
rect 25340 5966 25342 6018
rect 25342 5966 25394 6018
rect 25394 5966 25396 6018
rect 25340 5964 25396 5966
rect 25676 7586 25732 7588
rect 25676 7534 25678 7586
rect 25678 7534 25730 7586
rect 25730 7534 25732 7586
rect 25676 7532 25732 7534
rect 26572 7756 26628 7812
rect 26348 7644 26404 7700
rect 26124 7532 26180 7588
rect 27468 11788 27524 11844
rect 27244 11452 27300 11508
rect 27020 10610 27076 10612
rect 27020 10558 27022 10610
rect 27022 10558 27074 10610
rect 27074 10558 27076 10610
rect 27020 10556 27076 10558
rect 28588 12178 28644 12180
rect 28588 12126 28590 12178
rect 28590 12126 28642 12178
rect 28642 12126 28644 12178
rect 28588 12124 28644 12126
rect 27916 10556 27972 10612
rect 27356 9772 27412 9828
rect 27580 9884 27636 9940
rect 27244 8316 27300 8372
rect 28364 10108 28420 10164
rect 28140 9660 28196 9716
rect 28252 9826 28308 9828
rect 28252 9774 28254 9826
rect 28254 9774 28306 9826
rect 28306 9774 28308 9826
rect 28252 9772 28308 9774
rect 28252 9436 28308 9492
rect 23884 5122 23940 5124
rect 23884 5070 23886 5122
rect 23886 5070 23938 5122
rect 23938 5070 23940 5122
rect 23884 5068 23940 5070
rect 25452 5068 25508 5124
rect 27916 7474 27972 7476
rect 27916 7422 27918 7474
rect 27918 7422 27970 7474
rect 27970 7422 27972 7474
rect 27916 7420 27972 7422
rect 27580 6636 27636 6692
rect 28588 9714 28644 9716
rect 28588 9662 28590 9714
rect 28590 9662 28642 9714
rect 28642 9662 28644 9714
rect 28588 9660 28644 9662
rect 29596 16770 29652 16772
rect 29596 16718 29598 16770
rect 29598 16718 29650 16770
rect 29650 16718 29652 16770
rect 29596 16716 29652 16718
rect 29932 21756 29988 21812
rect 29820 20188 29876 20244
rect 29932 17106 29988 17108
rect 29932 17054 29934 17106
rect 29934 17054 29986 17106
rect 29986 17054 29988 17106
rect 29932 17052 29988 17054
rect 30044 16994 30100 16996
rect 30044 16942 30046 16994
rect 30046 16942 30098 16994
rect 30098 16942 30100 16994
rect 30044 16940 30100 16942
rect 30268 22988 30324 23044
rect 30492 22876 30548 22932
rect 30380 22764 30436 22820
rect 30492 22594 30548 22596
rect 30492 22542 30494 22594
rect 30494 22542 30546 22594
rect 30546 22542 30548 22594
rect 30492 22540 30548 22542
rect 30380 21868 30436 21924
rect 30492 21474 30548 21476
rect 30492 21422 30494 21474
rect 30494 21422 30546 21474
rect 30546 21422 30548 21474
rect 30492 21420 30548 21422
rect 30492 20578 30548 20580
rect 30492 20526 30494 20578
rect 30494 20526 30546 20578
rect 30546 20526 30548 20578
rect 30492 20524 30548 20526
rect 30380 16828 30436 16884
rect 30156 16156 30212 16212
rect 29484 15820 29540 15876
rect 29932 15820 29988 15876
rect 29932 15260 29988 15316
rect 29596 14642 29652 14644
rect 29596 14590 29598 14642
rect 29598 14590 29650 14642
rect 29650 14590 29652 14642
rect 29596 14588 29652 14590
rect 30156 15372 30212 15428
rect 32508 29986 32564 29988
rect 32508 29934 32510 29986
rect 32510 29934 32562 29986
rect 32562 29934 32564 29986
rect 32508 29932 32564 29934
rect 31948 29484 32004 29540
rect 32956 29708 33012 29764
rect 31276 29148 31332 29204
rect 32508 29148 32564 29204
rect 32620 28418 32676 28420
rect 32620 28366 32622 28418
rect 32622 28366 32674 28418
rect 32674 28366 32676 28418
rect 32620 28364 32676 28366
rect 32844 27916 32900 27972
rect 30716 25788 30772 25844
rect 31948 26908 32004 26964
rect 33404 28754 33460 28756
rect 33404 28702 33406 28754
rect 33406 28702 33458 28754
rect 33458 28702 33460 28754
rect 33404 28700 33460 28702
rect 33964 28364 34020 28420
rect 33628 27970 33684 27972
rect 33628 27918 33630 27970
rect 33630 27918 33682 27970
rect 33682 27918 33684 27970
rect 33628 27916 33684 27918
rect 31948 23938 32004 23940
rect 31948 23886 31950 23938
rect 31950 23886 32002 23938
rect 32002 23886 32004 23938
rect 31948 23884 32004 23886
rect 32172 25116 32228 25172
rect 31500 23772 31556 23828
rect 31276 23436 31332 23492
rect 31052 23212 31108 23268
rect 31164 23154 31220 23156
rect 31164 23102 31166 23154
rect 31166 23102 31218 23154
rect 31218 23102 31220 23154
rect 31164 23100 31220 23102
rect 31052 22540 31108 22596
rect 31612 22876 31668 22932
rect 30940 21980 30996 22036
rect 31164 20524 31220 20580
rect 30716 20188 30772 20244
rect 31388 21980 31444 22036
rect 31500 21868 31556 21924
rect 31948 22258 32004 22260
rect 31948 22206 31950 22258
rect 31950 22206 32002 22258
rect 32002 22206 32004 22258
rect 31948 22204 32004 22206
rect 31836 22146 31892 22148
rect 31836 22094 31838 22146
rect 31838 22094 31890 22146
rect 31890 22094 31892 22146
rect 31836 22092 31892 22094
rect 31724 21980 31780 22036
rect 32284 23938 32340 23940
rect 32284 23886 32286 23938
rect 32286 23886 32338 23938
rect 32338 23886 32340 23938
rect 32284 23884 32340 23886
rect 32844 23884 32900 23940
rect 32284 22988 32340 23044
rect 33068 23826 33124 23828
rect 33068 23774 33070 23826
rect 33070 23774 33122 23826
rect 33122 23774 33124 23826
rect 33068 23772 33124 23774
rect 32060 21980 32116 22036
rect 31836 21868 31892 21924
rect 31724 21644 31780 21700
rect 31836 21308 31892 21364
rect 32508 21868 32564 21924
rect 32508 21532 32564 21588
rect 31276 19628 31332 19684
rect 31164 19458 31220 19460
rect 31164 19406 31166 19458
rect 31166 19406 31218 19458
rect 31218 19406 31220 19458
rect 31164 19404 31220 19406
rect 31500 19458 31556 19460
rect 31500 19406 31502 19458
rect 31502 19406 31554 19458
rect 31554 19406 31556 19458
rect 31500 19404 31556 19406
rect 31612 18732 31668 18788
rect 32060 19234 32116 19236
rect 32060 19182 32062 19234
rect 32062 19182 32114 19234
rect 32114 19182 32116 19234
rect 32060 19180 32116 19182
rect 30268 15260 30324 15316
rect 30716 17052 30772 17108
rect 29708 14418 29764 14420
rect 29708 14366 29710 14418
rect 29710 14366 29762 14418
rect 29762 14366 29764 14418
rect 29708 14364 29764 14366
rect 29372 12796 29428 12852
rect 29148 12290 29204 12292
rect 29148 12238 29150 12290
rect 29150 12238 29202 12290
rect 29202 12238 29204 12290
rect 29148 12236 29204 12238
rect 29932 12962 29988 12964
rect 29932 12910 29934 12962
rect 29934 12910 29986 12962
rect 29986 12910 29988 12962
rect 29932 12908 29988 12910
rect 30044 12850 30100 12852
rect 30044 12798 30046 12850
rect 30046 12798 30098 12850
rect 30098 12798 30100 12850
rect 30044 12796 30100 12798
rect 30492 15484 30548 15540
rect 30940 16994 30996 16996
rect 30940 16942 30942 16994
rect 30942 16942 30994 16994
rect 30994 16942 30996 16994
rect 30940 16940 30996 16942
rect 31164 16828 31220 16884
rect 31388 16716 31444 16772
rect 31388 16156 31444 16212
rect 31164 16044 31220 16100
rect 31052 15372 31108 15428
rect 30940 14642 30996 14644
rect 30940 14590 30942 14642
rect 30942 14590 30994 14642
rect 30994 14590 30996 14642
rect 30940 14588 30996 14590
rect 30604 14418 30660 14420
rect 30604 14366 30606 14418
rect 30606 14366 30658 14418
rect 30658 14366 30660 14418
rect 30604 14364 30660 14366
rect 30380 14306 30436 14308
rect 30380 14254 30382 14306
rect 30382 14254 30434 14306
rect 30434 14254 30436 14306
rect 30380 14252 30436 14254
rect 31052 14306 31108 14308
rect 31052 14254 31054 14306
rect 31054 14254 31106 14306
rect 31106 14254 31108 14306
rect 31052 14252 31108 14254
rect 31388 15484 31444 15540
rect 30940 12962 30996 12964
rect 30940 12910 30942 12962
rect 30942 12910 30994 12962
rect 30994 12910 30996 12962
rect 30940 12908 30996 12910
rect 30716 12850 30772 12852
rect 30716 12798 30718 12850
rect 30718 12798 30770 12850
rect 30770 12798 30772 12850
rect 30716 12796 30772 12798
rect 30828 12572 30884 12628
rect 30268 12402 30324 12404
rect 30268 12350 30270 12402
rect 30270 12350 30322 12402
rect 30322 12350 30324 12402
rect 30268 12348 30324 12350
rect 30156 11452 30212 11508
rect 29708 11116 29764 11172
rect 29036 10610 29092 10612
rect 29036 10558 29038 10610
rect 29038 10558 29090 10610
rect 29090 10558 29092 10610
rect 29036 10556 29092 10558
rect 29148 9996 29204 10052
rect 29820 10610 29876 10612
rect 29820 10558 29822 10610
rect 29822 10558 29874 10610
rect 29874 10558 29876 10610
rect 29820 10556 29876 10558
rect 29596 10108 29652 10164
rect 29148 9826 29204 9828
rect 29148 9774 29150 9826
rect 29150 9774 29202 9826
rect 29202 9774 29204 9826
rect 29148 9772 29204 9774
rect 28588 7698 28644 7700
rect 28588 7646 28590 7698
rect 28590 7646 28642 7698
rect 28642 7646 28644 7698
rect 28588 7644 28644 7646
rect 28476 7532 28532 7588
rect 28140 6412 28196 6468
rect 28588 7362 28644 7364
rect 28588 7310 28590 7362
rect 28590 7310 28642 7362
rect 28642 7310 28644 7362
rect 28588 7308 28644 7310
rect 28364 6300 28420 6356
rect 28588 5404 28644 5460
rect 26796 5234 26852 5236
rect 26796 5182 26798 5234
rect 26798 5182 26850 5234
rect 26850 5182 26852 5234
rect 26796 5180 26852 5182
rect 27244 5234 27300 5236
rect 27244 5182 27246 5234
rect 27246 5182 27298 5234
rect 27298 5182 27300 5234
rect 27244 5180 27300 5182
rect 29932 10332 29988 10388
rect 29484 8764 29540 8820
rect 29820 9324 29876 9380
rect 30492 10050 30548 10052
rect 30492 9998 30494 10050
rect 30494 9998 30546 10050
rect 30546 9998 30548 10050
rect 30492 9996 30548 9998
rect 30156 8764 30212 8820
rect 30492 8316 30548 8372
rect 29932 8258 29988 8260
rect 29932 8206 29934 8258
rect 29934 8206 29986 8258
rect 29986 8206 29988 8258
rect 29932 8204 29988 8206
rect 29260 8092 29316 8148
rect 29596 7698 29652 7700
rect 29596 7646 29598 7698
rect 29598 7646 29650 7698
rect 29650 7646 29652 7698
rect 29596 7644 29652 7646
rect 30156 7586 30212 7588
rect 30156 7534 30158 7586
rect 30158 7534 30210 7586
rect 30210 7534 30212 7586
rect 30156 7532 30212 7534
rect 28812 7474 28868 7476
rect 28812 7422 28814 7474
rect 28814 7422 28866 7474
rect 28866 7422 28868 7474
rect 28812 7420 28868 7422
rect 29372 7474 29428 7476
rect 29372 7422 29374 7474
rect 29374 7422 29426 7474
rect 29426 7422 29428 7474
rect 29372 7420 29428 7422
rect 29820 7420 29876 7476
rect 29596 7362 29652 7364
rect 29596 7310 29598 7362
rect 29598 7310 29650 7362
rect 29650 7310 29652 7362
rect 29596 7308 29652 7310
rect 29708 6914 29764 6916
rect 29708 6862 29710 6914
rect 29710 6862 29762 6914
rect 29762 6862 29764 6914
rect 29708 6860 29764 6862
rect 29372 6690 29428 6692
rect 29372 6638 29374 6690
rect 29374 6638 29426 6690
rect 29426 6638 29428 6690
rect 29372 6636 29428 6638
rect 28588 5234 28644 5236
rect 28588 5182 28590 5234
rect 28590 5182 28642 5234
rect 28642 5182 28644 5234
rect 28588 5180 28644 5182
rect 26124 5068 26180 5124
rect 28364 4284 28420 4340
rect 28812 6412 28868 6468
rect 28812 5292 28868 5348
rect 29596 6466 29652 6468
rect 29596 6414 29598 6466
rect 29598 6414 29650 6466
rect 29650 6414 29652 6466
rect 29596 6412 29652 6414
rect 29260 5404 29316 5460
rect 29036 4338 29092 4340
rect 29036 4286 29038 4338
rect 29038 4286 29090 4338
rect 29090 4286 29092 4338
rect 29036 4284 29092 4286
rect 31276 9826 31332 9828
rect 31276 9774 31278 9826
rect 31278 9774 31330 9826
rect 31330 9774 31332 9826
rect 31276 9772 31332 9774
rect 31276 9548 31332 9604
rect 30828 9212 30884 9268
rect 31052 8540 31108 8596
rect 30828 8034 30884 8036
rect 30828 7982 30830 8034
rect 30830 7982 30882 8034
rect 30882 7982 30884 8034
rect 30828 7980 30884 7982
rect 31052 8034 31108 8036
rect 31052 7982 31054 8034
rect 31054 7982 31106 8034
rect 31106 7982 31108 8034
rect 31052 7980 31108 7982
rect 30940 7756 30996 7812
rect 30604 7420 30660 7476
rect 31276 7644 31332 7700
rect 31612 18226 31668 18228
rect 31612 18174 31614 18226
rect 31614 18174 31666 18226
rect 31666 18174 31668 18226
rect 31612 18172 31668 18174
rect 32284 18450 32340 18452
rect 32284 18398 32286 18450
rect 32286 18398 32338 18450
rect 32338 18398 32340 18450
rect 32284 18396 32340 18398
rect 33180 21698 33236 21700
rect 33180 21646 33182 21698
rect 33182 21646 33234 21698
rect 33234 21646 33236 21698
rect 33180 21644 33236 21646
rect 34748 34914 34804 34916
rect 34748 34862 34750 34914
rect 34750 34862 34802 34914
rect 34802 34862 34804 34914
rect 34748 34860 34804 34862
rect 34860 32508 34916 32564
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34748 32450 34804 32452
rect 34748 32398 34750 32450
rect 34750 32398 34802 32450
rect 34802 32398 34804 32450
rect 34748 32396 34804 32398
rect 34748 31724 34804 31780
rect 35308 33346 35364 33348
rect 35308 33294 35310 33346
rect 35310 33294 35362 33346
rect 35362 33294 35364 33346
rect 35308 33292 35364 33294
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35532 31890 35588 31892
rect 35532 31838 35534 31890
rect 35534 31838 35586 31890
rect 35586 31838 35588 31890
rect 35532 31836 35588 31838
rect 35644 31724 35700 31780
rect 35532 31666 35588 31668
rect 35532 31614 35534 31666
rect 35534 31614 35586 31666
rect 35586 31614 35588 31666
rect 35532 31612 35588 31614
rect 37548 34860 37604 34916
rect 36316 33516 36372 33572
rect 37212 33516 37268 33572
rect 37212 33292 37268 33348
rect 35868 32060 35924 32116
rect 37100 32396 37156 32452
rect 36988 31890 37044 31892
rect 36988 31838 36990 31890
rect 36990 31838 37042 31890
rect 37042 31838 37044 31890
rect 36988 31836 37044 31838
rect 34300 31164 34356 31220
rect 34188 29596 34244 29652
rect 35644 31554 35700 31556
rect 35644 31502 35646 31554
rect 35646 31502 35698 31554
rect 35698 31502 35700 31554
rect 35644 31500 35700 31502
rect 36540 31612 36596 31668
rect 35084 30828 35140 30884
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35868 30940 35924 30996
rect 37212 31554 37268 31556
rect 37212 31502 37214 31554
rect 37214 31502 37266 31554
rect 37266 31502 37268 31554
rect 37212 31500 37268 31502
rect 36988 30268 37044 30324
rect 39564 32450 39620 32452
rect 39564 32398 39566 32450
rect 39566 32398 39618 32450
rect 39618 32398 39620 32450
rect 39564 32396 39620 32398
rect 37772 30940 37828 30996
rect 39228 30940 39284 30996
rect 36988 30044 37044 30100
rect 35756 29596 35812 29652
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 27186 35252 27188
rect 35196 27134 35198 27186
rect 35198 27134 35250 27186
rect 35250 27134 35252 27186
rect 35196 27132 35252 27134
rect 34748 26908 34804 26964
rect 36428 29986 36484 29988
rect 36428 29934 36430 29986
rect 36430 29934 36482 29986
rect 36482 29934 36484 29986
rect 36428 29932 36484 29934
rect 36428 29484 36484 29540
rect 36764 29708 36820 29764
rect 36876 29650 36932 29652
rect 36876 29598 36878 29650
rect 36878 29598 36930 29650
rect 36930 29598 36932 29650
rect 36876 29596 36932 29598
rect 35980 27244 36036 27300
rect 36316 28476 36372 28532
rect 35532 26796 35588 26852
rect 34636 26514 34692 26516
rect 34636 26462 34638 26514
rect 34638 26462 34690 26514
rect 34690 26462 34692 26514
rect 34636 26460 34692 26462
rect 35756 27132 35812 27188
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34076 25452 34132 25508
rect 36092 27074 36148 27076
rect 36092 27022 36094 27074
rect 36094 27022 36146 27074
rect 36146 27022 36148 27074
rect 36092 27020 36148 27022
rect 35756 26908 35812 26964
rect 36204 26962 36260 26964
rect 36204 26910 36206 26962
rect 36206 26910 36258 26962
rect 36258 26910 36260 26962
rect 36204 26908 36260 26910
rect 37100 27916 37156 27972
rect 37324 30044 37380 30100
rect 37436 29932 37492 29988
rect 37660 29708 37716 29764
rect 38668 30098 38724 30100
rect 38668 30046 38670 30098
rect 38670 30046 38722 30098
rect 38722 30046 38724 30098
rect 38668 30044 38724 30046
rect 39004 29986 39060 29988
rect 39004 29934 39006 29986
rect 39006 29934 39058 29986
rect 39058 29934 39060 29986
rect 39004 29932 39060 29934
rect 37996 29538 38052 29540
rect 37996 29486 37998 29538
rect 37998 29486 38050 29538
rect 38050 29486 38052 29538
rect 37996 29484 38052 29486
rect 37660 28476 37716 28532
rect 36988 26962 37044 26964
rect 36988 26910 36990 26962
rect 36990 26910 37042 26962
rect 37042 26910 37044 26962
rect 36988 26908 37044 26910
rect 36428 26796 36484 26852
rect 35868 26236 35924 26292
rect 35644 24780 35700 24836
rect 36764 26290 36820 26292
rect 36764 26238 36766 26290
rect 36766 26238 36818 26290
rect 36818 26238 36820 26290
rect 36764 26236 36820 26238
rect 36092 24722 36148 24724
rect 36092 24670 36094 24722
rect 36094 24670 36146 24722
rect 36146 24670 36148 24722
rect 36092 24668 36148 24670
rect 36428 24780 36484 24836
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 24050 35252 24052
rect 35196 23998 35198 24050
rect 35198 23998 35250 24050
rect 35250 23998 35252 24050
rect 35196 23996 35252 23998
rect 35980 24108 36036 24164
rect 36092 23996 36148 24052
rect 35868 23884 35924 23940
rect 34076 23042 34132 23044
rect 34076 22990 34078 23042
rect 34078 22990 34130 23042
rect 34130 22990 34132 23042
rect 34076 22988 34132 22990
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35756 22482 35812 22484
rect 35756 22430 35758 22482
rect 35758 22430 35810 22482
rect 35810 22430 35812 22482
rect 35756 22428 35812 22430
rect 35532 22092 35588 22148
rect 36428 23772 36484 23828
rect 36428 23212 36484 23268
rect 37100 24722 37156 24724
rect 37100 24670 37102 24722
rect 37102 24670 37154 24722
rect 37154 24670 37156 24722
rect 37100 24668 37156 24670
rect 37100 23996 37156 24052
rect 36764 23100 36820 23156
rect 38556 27916 38612 27972
rect 37436 26796 37492 26852
rect 38108 27746 38164 27748
rect 38108 27694 38110 27746
rect 38110 27694 38162 27746
rect 38162 27694 38164 27746
rect 38108 27692 38164 27694
rect 38332 27074 38388 27076
rect 38332 27022 38334 27074
rect 38334 27022 38386 27074
rect 38386 27022 38388 27074
rect 38332 27020 38388 27022
rect 39004 27244 39060 27300
rect 39228 27692 39284 27748
rect 38332 26796 38388 26852
rect 37436 23938 37492 23940
rect 37436 23886 37438 23938
rect 37438 23886 37490 23938
rect 37490 23886 37492 23938
rect 37436 23884 37492 23886
rect 37548 23826 37604 23828
rect 37548 23774 37550 23826
rect 37550 23774 37602 23826
rect 37602 23774 37604 23826
rect 37548 23772 37604 23774
rect 36428 22428 36484 22484
rect 36092 22316 36148 22372
rect 37100 23266 37156 23268
rect 37100 23214 37102 23266
rect 37102 23214 37154 23266
rect 37154 23214 37156 23266
rect 37100 23212 37156 23214
rect 37324 23154 37380 23156
rect 37324 23102 37326 23154
rect 37326 23102 37378 23154
rect 37378 23102 37380 23154
rect 37324 23100 37380 23102
rect 37436 22370 37492 22372
rect 37436 22318 37438 22370
rect 37438 22318 37490 22370
rect 37490 22318 37492 22370
rect 37436 22316 37492 22318
rect 37772 23436 37828 23492
rect 38108 23996 38164 24052
rect 38892 23772 38948 23828
rect 37772 22540 37828 22596
rect 36092 21980 36148 22036
rect 36428 21474 36484 21476
rect 36428 21422 36430 21474
rect 36430 21422 36482 21474
rect 36482 21422 36484 21474
rect 36428 21420 36484 21422
rect 35868 21308 35924 21364
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 33740 20578 33796 20580
rect 33740 20526 33742 20578
rect 33742 20526 33794 20578
rect 33794 20526 33796 20578
rect 33740 20524 33796 20526
rect 37100 20578 37156 20580
rect 37100 20526 37102 20578
rect 37102 20526 37154 20578
rect 37154 20526 37156 20578
rect 37100 20524 37156 20526
rect 37772 20524 37828 20580
rect 35756 20076 35812 20132
rect 35980 19852 36036 19908
rect 37548 19852 37604 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 33404 19458 33460 19460
rect 33404 19406 33406 19458
rect 33406 19406 33458 19458
rect 33458 19406 33460 19458
rect 33404 19404 33460 19406
rect 33404 19234 33460 19236
rect 33404 19182 33406 19234
rect 33406 19182 33458 19234
rect 33458 19182 33460 19234
rect 33404 19180 33460 19182
rect 36204 19122 36260 19124
rect 36204 19070 36206 19122
rect 36206 19070 36258 19122
rect 36258 19070 36260 19122
rect 36204 19068 36260 19070
rect 37548 19346 37604 19348
rect 37548 19294 37550 19346
rect 37550 19294 37602 19346
rect 37602 19294 37604 19346
rect 37548 19292 37604 19294
rect 38332 19292 38388 19348
rect 37324 19068 37380 19124
rect 33068 18396 33124 18452
rect 31724 17052 31780 17108
rect 31612 16492 31668 16548
rect 32060 17106 32116 17108
rect 32060 17054 32062 17106
rect 32062 17054 32114 17106
rect 32114 17054 32116 17106
rect 32060 17052 32116 17054
rect 32284 16604 32340 16660
rect 31836 16268 31892 16324
rect 31948 15484 32004 15540
rect 32620 15932 32676 15988
rect 31724 15036 31780 15092
rect 31500 12348 31556 12404
rect 31612 12572 31668 12628
rect 32620 12962 32676 12964
rect 32620 12910 32622 12962
rect 32622 12910 32674 12962
rect 32674 12910 32676 12962
rect 32620 12908 32676 12910
rect 32732 15036 32788 15092
rect 32396 12738 32452 12740
rect 32396 12686 32398 12738
rect 32398 12686 32450 12738
rect 32450 12686 32452 12738
rect 32396 12684 32452 12686
rect 31724 12348 31780 12404
rect 33068 15036 33124 15092
rect 33292 17724 33348 17780
rect 33292 16940 33348 16996
rect 33964 18338 34020 18340
rect 33964 18286 33966 18338
rect 33966 18286 34018 18338
rect 34018 18286 34020 18338
rect 33964 18284 34020 18286
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 33628 16492 33684 16548
rect 35980 18338 36036 18340
rect 35980 18286 35982 18338
rect 35982 18286 36034 18338
rect 36034 18286 36036 18338
rect 35980 18284 36036 18286
rect 36316 18450 36372 18452
rect 36316 18398 36318 18450
rect 36318 18398 36370 18450
rect 36370 18398 36372 18450
rect 36316 18396 36372 18398
rect 36092 18060 36148 18116
rect 36540 17836 36596 17892
rect 37324 18508 37380 18564
rect 37100 18284 37156 18340
rect 37212 18060 37268 18116
rect 37212 17836 37268 17892
rect 37100 17778 37156 17780
rect 37100 17726 37102 17778
rect 37102 17726 37154 17778
rect 37154 17726 37156 17778
rect 37100 17724 37156 17726
rect 37212 17666 37268 17668
rect 37212 17614 37214 17666
rect 37214 17614 37266 17666
rect 37266 17614 37268 17666
rect 37212 17612 37268 17614
rect 35756 17388 35812 17444
rect 38108 18562 38164 18564
rect 38108 18510 38110 18562
rect 38110 18510 38162 18562
rect 38162 18510 38164 18562
rect 38108 18508 38164 18510
rect 38220 18450 38276 18452
rect 38220 18398 38222 18450
rect 38222 18398 38274 18450
rect 38274 18398 38276 18450
rect 38220 18396 38276 18398
rect 37436 18060 37492 18116
rect 37996 17554 38052 17556
rect 37996 17502 37998 17554
rect 37998 17502 38050 17554
rect 38050 17502 38052 17554
rect 37996 17500 38052 17502
rect 37660 17442 37716 17444
rect 37660 17390 37662 17442
rect 37662 17390 37714 17442
rect 37714 17390 37716 17442
rect 37660 17388 37716 17390
rect 35308 16828 35364 16884
rect 35868 16716 35924 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34636 16268 34692 16324
rect 34412 16098 34468 16100
rect 34412 16046 34414 16098
rect 34414 16046 34466 16098
rect 34466 16046 34468 16098
rect 34412 16044 34468 16046
rect 33404 15932 33460 15988
rect 33292 13804 33348 13860
rect 34412 13804 34468 13860
rect 33180 13468 33236 13524
rect 33628 13244 33684 13300
rect 33404 12908 33460 12964
rect 33068 12738 33124 12740
rect 33068 12686 33070 12738
rect 33070 12686 33122 12738
rect 33122 12686 33124 12738
rect 33068 12684 33124 12686
rect 33404 12684 33460 12740
rect 32060 11170 32116 11172
rect 32060 11118 32062 11170
rect 32062 11118 32114 11170
rect 32114 11118 32116 11170
rect 32060 11116 32116 11118
rect 31836 10108 31892 10164
rect 32508 10610 32564 10612
rect 32508 10558 32510 10610
rect 32510 10558 32562 10610
rect 32562 10558 32564 10610
rect 32508 10556 32564 10558
rect 33180 11116 33236 11172
rect 34188 12962 34244 12964
rect 34188 12910 34190 12962
rect 34190 12910 34242 12962
rect 34242 12910 34244 12962
rect 34188 12908 34244 12910
rect 34300 12796 34356 12852
rect 33964 12348 34020 12404
rect 34076 12290 34132 12292
rect 34076 12238 34078 12290
rect 34078 12238 34130 12290
rect 34130 12238 34132 12290
rect 34076 12236 34132 12238
rect 34524 12572 34580 12628
rect 32172 9884 32228 9940
rect 31724 9436 31780 9492
rect 32508 10220 32564 10276
rect 33516 10722 33572 10724
rect 33516 10670 33518 10722
rect 33518 10670 33570 10722
rect 33570 10670 33572 10722
rect 33516 10668 33572 10670
rect 33740 10610 33796 10612
rect 33740 10558 33742 10610
rect 33742 10558 33794 10610
rect 33794 10558 33796 10610
rect 33740 10556 33796 10558
rect 33516 10332 33572 10388
rect 33628 10220 33684 10276
rect 32508 9772 32564 9828
rect 32284 9660 32340 9716
rect 32172 9548 32228 9604
rect 31836 9100 31892 9156
rect 31724 7756 31780 7812
rect 32620 9714 32676 9716
rect 32620 9662 32622 9714
rect 32622 9662 32674 9714
rect 32674 9662 32676 9714
rect 32620 9660 32676 9662
rect 33068 9660 33124 9716
rect 32732 9324 32788 9380
rect 32844 9548 32900 9604
rect 32620 8316 32676 8372
rect 32732 8092 32788 8148
rect 32172 7698 32228 7700
rect 32172 7646 32174 7698
rect 32174 7646 32226 7698
rect 32226 7646 32228 7698
rect 32172 7644 32228 7646
rect 32508 7474 32564 7476
rect 32508 7422 32510 7474
rect 32510 7422 32562 7474
rect 32562 7422 32564 7474
rect 32508 7420 32564 7422
rect 31948 6860 32004 6916
rect 31612 6524 31668 6580
rect 31276 5068 31332 5124
rect 31500 3500 31556 3556
rect 18508 3442 18564 3444
rect 18508 3390 18510 3442
rect 18510 3390 18562 3442
rect 18562 3390 18564 3442
rect 18508 3388 18564 3390
rect 31052 3442 31108 3444
rect 31052 3390 31054 3442
rect 31054 3390 31106 3442
rect 31106 3390 31108 3442
rect 31052 3388 31108 3390
rect 32284 6188 32340 6244
rect 32060 5852 32116 5908
rect 32732 5740 32788 5796
rect 32060 5180 32116 5236
rect 31948 4450 32004 4452
rect 31948 4398 31950 4450
rect 31950 4398 32002 4450
rect 32002 4398 32004 4450
rect 31948 4396 32004 4398
rect 32620 4620 32676 4676
rect 33292 9884 33348 9940
rect 33292 9602 33348 9604
rect 33292 9550 33294 9602
rect 33294 9550 33346 9602
rect 33346 9550 33348 9602
rect 33292 9548 33348 9550
rect 33180 7756 33236 7812
rect 33404 8258 33460 8260
rect 33404 8206 33406 8258
rect 33406 8206 33458 8258
rect 33458 8206 33460 8258
rect 33404 8204 33460 8206
rect 33516 7756 33572 7812
rect 33964 10444 34020 10500
rect 34076 9154 34132 9156
rect 34076 9102 34078 9154
rect 34078 9102 34130 9154
rect 34130 9102 34132 9154
rect 34076 9100 34132 9102
rect 33852 7532 33908 7588
rect 33628 7420 33684 7476
rect 33852 6412 33908 6468
rect 34300 9436 34356 9492
rect 35532 16268 35588 16324
rect 34860 15986 34916 15988
rect 34860 15934 34862 15986
rect 34862 15934 34914 15986
rect 34914 15934 34916 15986
rect 34860 15932 34916 15934
rect 35196 15986 35252 15988
rect 35196 15934 35198 15986
rect 35198 15934 35250 15986
rect 35250 15934 35252 15986
rect 35196 15932 35252 15934
rect 35868 15986 35924 15988
rect 35868 15934 35870 15986
rect 35870 15934 35922 15986
rect 35922 15934 35924 15986
rect 35868 15932 35924 15934
rect 36316 16044 36372 16100
rect 37212 16770 37268 16772
rect 37212 16718 37214 16770
rect 37214 16718 37266 16770
rect 37266 16718 37268 16770
rect 37212 16716 37268 16718
rect 35308 15036 35364 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35532 14364 35588 14420
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 34748 12796 34804 12852
rect 34972 12908 35028 12964
rect 34860 12572 34916 12628
rect 34860 9772 34916 9828
rect 34636 9042 34692 9044
rect 34636 8990 34638 9042
rect 34638 8990 34690 9042
rect 34690 8990 34692 9042
rect 34636 8988 34692 8990
rect 34524 8258 34580 8260
rect 34524 8206 34526 8258
rect 34526 8206 34578 8258
rect 34578 8206 34580 8258
rect 34524 8204 34580 8206
rect 34412 6860 34468 6916
rect 35196 12738 35252 12740
rect 35196 12686 35198 12738
rect 35198 12686 35250 12738
rect 35250 12686 35252 12738
rect 35196 12684 35252 12686
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35868 13858 35924 13860
rect 35868 13806 35870 13858
rect 35870 13806 35922 13858
rect 35922 13806 35924 13858
rect 35868 13804 35924 13806
rect 35644 12908 35700 12964
rect 35868 12572 35924 12628
rect 36428 13916 36484 13972
rect 35532 11564 35588 11620
rect 35420 11116 35476 11172
rect 35308 10610 35364 10612
rect 35308 10558 35310 10610
rect 35310 10558 35362 10610
rect 35362 10558 35364 10610
rect 35308 10556 35364 10558
rect 35084 10444 35140 10500
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35756 10556 35812 10612
rect 35644 9548 35700 9604
rect 36204 10780 36260 10836
rect 36764 13468 36820 13524
rect 36540 10892 36596 10948
rect 35980 10498 36036 10500
rect 35980 10446 35982 10498
rect 35982 10446 36034 10498
rect 36034 10446 36036 10498
rect 35980 10444 36036 10446
rect 36428 10108 36484 10164
rect 36316 9772 36372 9828
rect 36316 9436 36372 9492
rect 35532 8988 35588 9044
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 36204 9042 36260 9044
rect 36204 8990 36206 9042
rect 36206 8990 36258 9042
rect 36258 8990 36260 9042
rect 36204 8988 36260 8990
rect 35980 8764 36036 8820
rect 36540 9884 36596 9940
rect 36652 9772 36708 9828
rect 36540 9100 36596 9156
rect 35868 8316 35924 8372
rect 34972 8092 35028 8148
rect 35756 8204 35812 8260
rect 35644 7586 35700 7588
rect 35644 7534 35646 7586
rect 35646 7534 35698 7586
rect 35698 7534 35700 7586
rect 35644 7532 35700 7534
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34860 6636 34916 6692
rect 34300 6578 34356 6580
rect 34300 6526 34302 6578
rect 34302 6526 34354 6578
rect 34354 6526 34356 6578
rect 34300 6524 34356 6526
rect 35532 6188 35588 6244
rect 36428 8428 36484 8484
rect 36316 8204 36372 8260
rect 35980 7586 36036 7588
rect 35980 7534 35982 7586
rect 35982 7534 36034 7586
rect 36034 7534 36036 7586
rect 35980 7532 36036 7534
rect 36204 6748 36260 6804
rect 36316 7868 36372 7924
rect 35868 6636 35924 6692
rect 33628 5794 33684 5796
rect 33628 5742 33630 5794
rect 33630 5742 33682 5794
rect 33682 5742 33684 5794
rect 33628 5740 33684 5742
rect 33852 5682 33908 5684
rect 33852 5630 33854 5682
rect 33854 5630 33906 5682
rect 33906 5630 33908 5682
rect 33852 5628 33908 5630
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35644 5292 35700 5348
rect 34524 5068 34580 5124
rect 35308 5068 35364 5124
rect 34076 4956 34132 5012
rect 33516 4450 33572 4452
rect 33516 4398 33518 4450
rect 33518 4398 33570 4450
rect 33570 4398 33572 4450
rect 33516 4396 33572 4398
rect 33404 3500 33460 3556
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 34524 4732 34580 4788
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35980 6300 36036 6356
rect 35868 5628 35924 5684
rect 35980 5740 36036 5796
rect 36204 5068 36260 5124
rect 35980 4898 36036 4900
rect 35980 4846 35982 4898
rect 35982 4846 36034 4898
rect 36034 4846 36036 4898
rect 35980 4844 36036 4846
rect 36652 8204 36708 8260
rect 36652 7980 36708 8036
rect 37436 16098 37492 16100
rect 37436 16046 37438 16098
rect 37438 16046 37490 16098
rect 37490 16046 37492 16098
rect 37436 16044 37492 16046
rect 37100 14252 37156 14308
rect 37660 13916 37716 13972
rect 37436 13858 37492 13860
rect 37436 13806 37438 13858
rect 37438 13806 37490 13858
rect 37490 13806 37492 13858
rect 37436 13804 37492 13806
rect 37324 13692 37380 13748
rect 36988 12908 37044 12964
rect 37212 12290 37268 12292
rect 37212 12238 37214 12290
rect 37214 12238 37266 12290
rect 37266 12238 37268 12290
rect 37212 12236 37268 12238
rect 37772 12850 37828 12852
rect 37772 12798 37774 12850
rect 37774 12798 37826 12850
rect 37826 12798 37828 12850
rect 37772 12796 37828 12798
rect 37884 14476 37940 14532
rect 37324 12012 37380 12068
rect 38108 14140 38164 14196
rect 38108 13468 38164 13524
rect 37996 11564 38052 11620
rect 37436 11170 37492 11172
rect 37436 11118 37438 11170
rect 37438 11118 37490 11170
rect 37490 11118 37492 11170
rect 37436 11116 37492 11118
rect 38108 11452 38164 11508
rect 37436 10834 37492 10836
rect 37436 10782 37438 10834
rect 37438 10782 37490 10834
rect 37490 10782 37492 10834
rect 37436 10780 37492 10782
rect 37660 11116 37716 11172
rect 37884 10892 37940 10948
rect 38108 10892 38164 10948
rect 38332 14252 38388 14308
rect 39116 22540 39172 22596
rect 38892 21420 38948 21476
rect 39564 21474 39620 21476
rect 39564 21422 39566 21474
rect 39566 21422 39618 21474
rect 39618 21422 39620 21474
rect 39564 21420 39620 21422
rect 38556 20524 38612 20580
rect 38556 15148 38612 15204
rect 39564 15202 39620 15204
rect 39564 15150 39566 15202
rect 39566 15150 39618 15202
rect 39618 15150 39620 15202
rect 39564 15148 39620 15150
rect 39676 14306 39732 14308
rect 39676 14254 39678 14306
rect 39678 14254 39730 14306
rect 39730 14254 39732 14306
rect 39676 14252 39732 14254
rect 38556 14140 38612 14196
rect 38444 13916 38500 13972
rect 38556 13858 38612 13860
rect 38556 13806 38558 13858
rect 38558 13806 38610 13858
rect 38610 13806 38612 13858
rect 38556 13804 38612 13806
rect 38892 13746 38948 13748
rect 38892 13694 38894 13746
rect 38894 13694 38946 13746
rect 38946 13694 38948 13746
rect 38892 13692 38948 13694
rect 39340 13468 39396 13524
rect 38444 12850 38500 12852
rect 38444 12798 38446 12850
rect 38446 12798 38498 12850
rect 38498 12798 38500 12850
rect 38444 12796 38500 12798
rect 38332 12012 38388 12068
rect 38556 11452 38612 11508
rect 38444 10780 38500 10836
rect 37212 9884 37268 9940
rect 37548 9826 37604 9828
rect 37548 9774 37550 9826
rect 37550 9774 37602 9826
rect 37602 9774 37604 9826
rect 37548 9772 37604 9774
rect 37212 9602 37268 9604
rect 37212 9550 37214 9602
rect 37214 9550 37266 9602
rect 37266 9550 37268 9602
rect 37212 9548 37268 9550
rect 37436 9602 37492 9604
rect 37436 9550 37438 9602
rect 37438 9550 37490 9602
rect 37490 9550 37492 9602
rect 37436 9548 37492 9550
rect 37100 9324 37156 9380
rect 37772 9324 37828 9380
rect 36988 9154 37044 9156
rect 36988 9102 36990 9154
rect 36990 9102 37042 9154
rect 37042 9102 37044 9154
rect 36988 9100 37044 9102
rect 36876 8764 36932 8820
rect 36988 8146 37044 8148
rect 36988 8094 36990 8146
rect 36990 8094 37042 8146
rect 37042 8094 37044 8146
rect 36988 8092 37044 8094
rect 37324 9154 37380 9156
rect 37324 9102 37326 9154
rect 37326 9102 37378 9154
rect 37378 9102 37380 9154
rect 37324 9100 37380 9102
rect 37324 8258 37380 8260
rect 37324 8206 37326 8258
rect 37326 8206 37378 8258
rect 37378 8206 37380 8258
rect 37324 8204 37380 8206
rect 36764 6412 36820 6468
rect 36876 6748 36932 6804
rect 36540 5852 36596 5908
rect 37212 7532 37268 7588
rect 36652 6188 36708 6244
rect 37324 6076 37380 6132
rect 37100 5010 37156 5012
rect 37100 4958 37102 5010
rect 37102 4958 37154 5010
rect 37154 4958 37156 5010
rect 37100 4956 37156 4958
rect 36764 4844 36820 4900
rect 38108 10108 38164 10164
rect 38780 10722 38836 10724
rect 38780 10670 38782 10722
rect 38782 10670 38834 10722
rect 38834 10670 38836 10722
rect 38780 10668 38836 10670
rect 38220 9772 38276 9828
rect 37996 9714 38052 9716
rect 37996 9662 37998 9714
rect 37998 9662 38050 9714
rect 38050 9662 38052 9714
rect 37996 9660 38052 9662
rect 38108 9324 38164 9380
rect 39116 10108 39172 10164
rect 39228 9826 39284 9828
rect 39228 9774 39230 9826
rect 39230 9774 39282 9826
rect 39282 9774 39284 9826
rect 39228 9772 39284 9774
rect 38892 9602 38948 9604
rect 38892 9550 38894 9602
rect 38894 9550 38946 9602
rect 38946 9550 38948 9602
rect 38892 9548 38948 9550
rect 39004 9436 39060 9492
rect 38332 9154 38388 9156
rect 38332 9102 38334 9154
rect 38334 9102 38386 9154
rect 38386 9102 38388 9154
rect 38332 9100 38388 9102
rect 37772 8316 37828 8372
rect 37996 8370 38052 8372
rect 37996 8318 37998 8370
rect 37998 8318 38050 8370
rect 38050 8318 38052 8370
rect 37996 8316 38052 8318
rect 37548 6524 37604 6580
rect 37660 5180 37716 5236
rect 38108 8092 38164 8148
rect 37996 7532 38052 7588
rect 37884 6188 37940 6244
rect 37772 4956 37828 5012
rect 37436 4844 37492 4900
rect 38332 8428 38388 8484
rect 38556 8204 38612 8260
rect 39228 8316 39284 8372
rect 38108 4620 38164 4676
rect 39228 8034 39284 8036
rect 39228 7982 39230 8034
rect 39230 7982 39282 8034
rect 39282 7982 39284 8034
rect 39228 7980 39284 7982
rect 39004 6860 39060 6916
rect 38892 6636 38948 6692
rect 36764 4396 36820 4452
rect 35420 3388 35476 3444
rect 37436 4226 37492 4228
rect 37436 4174 37438 4226
rect 37438 4174 37490 4226
rect 37490 4174 37492 4226
rect 37436 4172 37492 4174
rect 37996 3442 38052 3444
rect 37996 3390 37998 3442
rect 37998 3390 38050 3442
rect 38050 3390 38052 3442
rect 37996 3388 38052 3390
rect 39116 6300 39172 6356
rect 39340 6076 39396 6132
rect 39004 5292 39060 5348
rect 38780 4956 38836 5012
rect 38892 4172 38948 4228
rect 39228 5234 39284 5236
rect 39228 5182 39230 5234
rect 39230 5182 39282 5234
rect 39282 5182 39284 5234
rect 39228 5180 39284 5182
rect 39116 4732 39172 4788
rect 39452 3388 39508 3444
<< metal3 >>
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 17714 39676 17724 39732
rect 17780 39676 18620 39732
rect 18676 39676 18686 39732
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 11778 39004 11788 39060
rect 11844 39004 12908 39060
rect 12964 39004 13580 39060
rect 13636 39004 15372 39060
rect 15428 39004 15438 39060
rect 21298 38892 21308 38948
rect 21364 38892 22876 38948
rect 22932 38892 22942 38948
rect 9986 38780 9996 38836
rect 10052 38780 11340 38836
rect 11396 38780 12684 38836
rect 12740 38780 12750 38836
rect 16594 38780 16604 38836
rect 16660 38780 18172 38836
rect 18228 38780 18238 38836
rect 18386 38780 18396 38836
rect 18452 38780 20300 38836
rect 20356 38780 20972 38836
rect 21028 38780 21038 38836
rect 11666 38668 11676 38724
rect 11732 38668 12012 38724
rect 12068 38668 12078 38724
rect 12226 38556 12236 38612
rect 12292 38556 13804 38612
rect 13860 38556 13870 38612
rect 13122 38444 13132 38500
rect 13188 38444 16492 38500
rect 16548 38444 16558 38500
rect 20850 38444 20860 38500
rect 20916 38444 21644 38500
rect 21700 38444 21710 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16818 38332 16828 38388
rect 16884 38332 20076 38388
rect 20132 38332 20142 38388
rect 9650 38220 9660 38276
rect 9716 38220 10556 38276
rect 10612 38220 12012 38276
rect 12068 38220 17164 38276
rect 17220 38220 17836 38276
rect 17892 38220 17902 38276
rect 9986 38108 9996 38164
rect 10052 38108 14700 38164
rect 14756 38108 16156 38164
rect 16212 38108 16222 38164
rect 16482 38108 16492 38164
rect 16548 38108 17388 38164
rect 17444 38108 19292 38164
rect 19348 38108 19358 38164
rect 11554 37996 11564 38052
rect 11620 37996 13916 38052
rect 13972 37996 13982 38052
rect 14130 37996 14140 38052
rect 14196 37996 15932 38052
rect 15988 37996 21924 38052
rect 21868 37940 21924 37996
rect 12338 37884 12348 37940
rect 12404 37884 13468 37940
rect 13524 37884 13534 37940
rect 18162 37884 18172 37940
rect 18228 37884 18956 37940
rect 19012 37884 19022 37940
rect 21858 37884 21868 37940
rect 21924 37884 24108 37940
rect 24164 37884 24174 37940
rect 13010 37772 13020 37828
rect 13076 37772 13692 37828
rect 13748 37772 13758 37828
rect 16258 37772 16268 37828
rect 16324 37772 17388 37828
rect 17444 37772 17454 37828
rect 18722 37772 18732 37828
rect 18788 37772 19628 37828
rect 19684 37772 20524 37828
rect 20580 37772 20590 37828
rect 21746 37772 21756 37828
rect 21812 37772 22428 37828
rect 22484 37772 23100 37828
rect 23156 37772 23166 37828
rect 12786 37660 12796 37716
rect 12852 37660 13580 37716
rect 13636 37660 13646 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 15026 37548 15036 37604
rect 15092 37548 16828 37604
rect 16884 37548 16894 37604
rect 12226 37436 12236 37492
rect 12292 37436 13468 37492
rect 13524 37436 13534 37492
rect 16706 37436 16716 37492
rect 16772 37436 17500 37492
rect 17556 37436 17566 37492
rect 17602 37324 17612 37380
rect 17668 37324 22652 37380
rect 22708 37324 24444 37380
rect 24500 37324 24510 37380
rect 24658 37324 24668 37380
rect 24724 37324 28252 37380
rect 28308 37324 28812 37380
rect 28868 37324 28878 37380
rect 13906 37212 13916 37268
rect 13972 37212 14364 37268
rect 14420 37212 18060 37268
rect 18116 37212 18126 37268
rect 18274 37100 18284 37156
rect 18340 37100 19068 37156
rect 19124 37100 20412 37156
rect 20468 37100 21756 37156
rect 21812 37100 21822 37156
rect 24546 37100 24556 37156
rect 24612 37100 27580 37156
rect 27636 37100 27646 37156
rect 22194 36988 22204 37044
rect 22260 36988 25340 37044
rect 25396 36988 26236 37044
rect 26292 36988 26302 37044
rect 18386 36876 18396 36932
rect 18452 36876 20524 36932
rect 20580 36876 22428 36932
rect 22484 36876 22494 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 13346 36428 13356 36484
rect 13412 36428 14028 36484
rect 14084 36428 14094 36484
rect 22754 36428 22764 36484
rect 22820 36428 23436 36484
rect 23492 36428 23502 36484
rect 11554 36316 11564 36372
rect 11620 36316 13468 36372
rect 13524 36316 13534 36372
rect 24770 36316 24780 36372
rect 24836 36316 25564 36372
rect 25620 36316 25630 36372
rect 24210 36204 24220 36260
rect 24276 36204 24892 36260
rect 24948 36204 24958 36260
rect 33058 36204 33068 36260
rect 33124 36204 33740 36260
rect 33796 36204 33806 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 14700 35868 16604 35924
rect 16660 35868 16670 35924
rect 14700 35812 14756 35868
rect 13794 35756 13804 35812
rect 13860 35756 14476 35812
rect 14532 35756 14542 35812
rect 14690 35756 14700 35812
rect 14756 35756 14766 35812
rect 15092 35756 24332 35812
rect 24388 35756 25004 35812
rect 25060 35756 25070 35812
rect 25778 35756 25788 35812
rect 25844 35756 26684 35812
rect 26740 35756 33404 35812
rect 33460 35756 35084 35812
rect 35140 35756 35150 35812
rect 15092 35700 15148 35756
rect 14130 35644 14140 35700
rect 14196 35644 15148 35700
rect 19842 35644 19852 35700
rect 19908 35644 21420 35700
rect 21476 35644 22204 35700
rect 22260 35644 22270 35700
rect 12338 35532 12348 35588
rect 12404 35532 14364 35588
rect 14420 35532 14430 35588
rect 21186 35532 21196 35588
rect 21252 35532 21868 35588
rect 21924 35532 23212 35588
rect 23268 35532 23278 35588
rect 17490 35308 17500 35364
rect 17556 35308 18396 35364
rect 18452 35308 18462 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 5618 35196 5628 35252
rect 5684 35196 6188 35252
rect 6244 35196 9660 35252
rect 9716 35196 11788 35252
rect 11844 35196 11854 35252
rect 8978 35084 8988 35140
rect 9044 35084 12124 35140
rect 12180 35084 12190 35140
rect 6402 34972 6412 35028
rect 6468 34972 12012 35028
rect 12068 34972 12078 35028
rect 22866 34972 22876 35028
rect 22932 34972 23996 35028
rect 24052 34972 24062 35028
rect 25330 34972 25340 35028
rect 25396 34972 28364 35028
rect 28420 34972 31164 35028
rect 31220 34972 31230 35028
rect 14914 34860 14924 34916
rect 14980 34860 17276 34916
rect 17332 34860 17948 34916
rect 18004 34860 18014 34916
rect 31714 34860 31724 34916
rect 31780 34860 34748 34916
rect 34804 34860 37548 34916
rect 37604 34860 37614 34916
rect 12898 34748 12908 34804
rect 12964 34748 14812 34804
rect 14868 34748 14878 34804
rect 14914 34636 14924 34692
rect 14980 34636 16156 34692
rect 16212 34636 17612 34692
rect 17668 34636 17678 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 12450 34412 12460 34468
rect 12516 34412 14140 34468
rect 14196 34412 18620 34468
rect 18676 34412 18686 34468
rect 11554 34300 11564 34356
rect 11620 34300 12796 34356
rect 12852 34300 13468 34356
rect 13524 34300 13534 34356
rect 26852 34300 29148 34356
rect 29204 34300 29214 34356
rect 13570 34188 13580 34244
rect 13636 34188 14700 34244
rect 14756 34188 14766 34244
rect 14130 34076 14140 34132
rect 14196 34076 14588 34132
rect 14644 34076 14654 34132
rect 15026 34076 15036 34132
rect 15092 34076 15596 34132
rect 15652 34076 19628 34132
rect 19684 34076 19694 34132
rect 26852 34020 26908 34300
rect 30818 34188 30828 34244
rect 30884 34188 32172 34244
rect 32228 34188 32238 34244
rect 31154 34076 31164 34132
rect 31220 34076 34076 34132
rect 34132 34076 34142 34132
rect 9538 33964 9548 34020
rect 9604 33964 10444 34020
rect 10500 33964 11340 34020
rect 11396 33964 11406 34020
rect 18274 33964 18284 34020
rect 18340 33964 19180 34020
rect 19236 33964 19246 34020
rect 20962 33964 20972 34020
rect 21028 33964 21644 34020
rect 21700 33964 26908 34020
rect 29922 33964 29932 34020
rect 29988 33964 31052 34020
rect 31108 33964 31276 34020
rect 31332 33964 31342 34020
rect 16594 33852 16604 33908
rect 16660 33852 17836 33908
rect 17892 33852 21308 33908
rect 21364 33852 21756 33908
rect 21812 33852 21822 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 11330 33516 11340 33572
rect 11396 33516 12796 33572
rect 12852 33516 13916 33572
rect 13972 33516 13982 33572
rect 34066 33516 34076 33572
rect 34132 33516 36316 33572
rect 36372 33516 37212 33572
rect 37268 33516 37278 33572
rect 6850 33404 6860 33460
rect 6916 33404 17388 33460
rect 17444 33404 17454 33460
rect 19618 33404 19628 33460
rect 19684 33404 20300 33460
rect 20356 33404 20366 33460
rect 9314 33292 9324 33348
rect 9380 33292 12628 33348
rect 14242 33292 14252 33348
rect 14308 33292 15708 33348
rect 15764 33292 15774 33348
rect 18722 33292 18732 33348
rect 18788 33292 19068 33348
rect 19124 33292 20188 33348
rect 20244 33292 20254 33348
rect 20514 33292 20524 33348
rect 20580 33292 21308 33348
rect 21364 33292 21374 33348
rect 33170 33292 33180 33348
rect 33236 33292 35308 33348
rect 35364 33292 37212 33348
rect 37268 33292 37278 33348
rect 12572 33236 12628 33292
rect 8194 33180 8204 33236
rect 8260 33180 9660 33236
rect 9716 33180 9996 33236
rect 10052 33180 10062 33236
rect 12562 33180 12572 33236
rect 12628 33180 14140 33236
rect 14196 33180 14206 33236
rect 17238 33180 17276 33236
rect 17332 33180 17342 33236
rect 18274 33180 18284 33236
rect 18340 33180 19852 33236
rect 19908 33180 20636 33236
rect 20692 33180 20702 33236
rect 14578 33068 14588 33124
rect 14644 33068 15596 33124
rect 15652 33068 19516 33124
rect 19572 33068 19582 33124
rect 21410 33068 21420 33124
rect 21476 33068 22316 33124
rect 22372 33068 22382 33124
rect 24434 33068 24444 33124
rect 24500 33068 25452 33124
rect 25508 33068 25518 33124
rect 28242 33068 28252 33124
rect 28308 33068 29820 33124
rect 29876 33068 29886 33124
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 19618 32732 19628 32788
rect 19684 32732 21308 32788
rect 21364 32732 21374 32788
rect 23090 32732 23100 32788
rect 23156 32732 23548 32788
rect 23604 32732 25340 32788
rect 25396 32732 25406 32788
rect 29250 32732 29260 32788
rect 29316 32732 30380 32788
rect 30436 32732 30446 32788
rect 30594 32732 30604 32788
rect 30660 32732 32956 32788
rect 33012 32732 33022 32788
rect 23650 32620 23660 32676
rect 23716 32620 25116 32676
rect 25172 32620 25182 32676
rect 26450 32508 26460 32564
rect 26516 32508 28140 32564
rect 28196 32508 28206 32564
rect 29474 32508 29484 32564
rect 29540 32508 30492 32564
rect 30548 32508 30558 32564
rect 31826 32508 31836 32564
rect 31892 32508 33292 32564
rect 33348 32508 34076 32564
rect 34132 32508 34860 32564
rect 34916 32508 34926 32564
rect 27570 32396 27580 32452
rect 27636 32396 29596 32452
rect 29652 32396 30268 32452
rect 30324 32396 30334 32452
rect 32274 32396 32284 32452
rect 32340 32396 33180 32452
rect 33236 32396 33246 32452
rect 34738 32396 34748 32452
rect 34804 32396 37100 32452
rect 37156 32396 39564 32452
rect 39620 32396 39630 32452
rect 19506 32284 19516 32340
rect 19572 32284 21644 32340
rect 21700 32284 21710 32340
rect 17266 32172 17276 32228
rect 17332 32172 17724 32228
rect 17780 32172 17790 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 31378 32060 31388 32116
rect 31444 32060 31454 32116
rect 35858 32060 35868 32116
rect 35924 32060 37268 32116
rect 28578 31948 28588 32004
rect 28644 31948 30828 32004
rect 30884 31948 30894 32004
rect 31388 31892 31444 32060
rect 11218 31836 11228 31892
rect 11284 31836 11788 31892
rect 11844 31836 11854 31892
rect 12002 31836 12012 31892
rect 12068 31836 12572 31892
rect 12628 31836 12638 31892
rect 14018 31836 14028 31892
rect 14084 31836 17388 31892
rect 17444 31836 17948 31892
rect 18004 31836 18014 31892
rect 31388 31836 32004 31892
rect 35522 31836 35532 31892
rect 35588 31836 36988 31892
rect 37044 31836 37054 31892
rect 31948 31780 32004 31836
rect 11554 31724 11564 31780
rect 11620 31724 12124 31780
rect 12180 31724 12190 31780
rect 12674 31724 12684 31780
rect 12740 31724 14924 31780
rect 14980 31724 14990 31780
rect 30594 31724 30604 31780
rect 30660 31724 30940 31780
rect 30996 31724 31006 31780
rect 31266 31724 31276 31780
rect 31332 31724 31724 31780
rect 31780 31724 31790 31780
rect 31938 31724 31948 31780
rect 32004 31724 34748 31780
rect 34804 31724 35644 31780
rect 35700 31724 35710 31780
rect 14802 31612 14812 31668
rect 14868 31612 16156 31668
rect 16212 31612 16222 31668
rect 18050 31612 18060 31668
rect 18116 31612 18620 31668
rect 18676 31612 18686 31668
rect 34066 31612 34076 31668
rect 34132 31612 35532 31668
rect 35588 31612 36540 31668
rect 36596 31612 36606 31668
rect 37212 31556 37268 32060
rect 13570 31500 13580 31556
rect 13636 31500 14700 31556
rect 14756 31500 14766 31556
rect 16258 31500 16268 31556
rect 16324 31500 17276 31556
rect 17332 31500 17342 31556
rect 17490 31500 17500 31556
rect 17556 31500 18956 31556
rect 19012 31500 19022 31556
rect 31892 31500 35644 31556
rect 35700 31500 35710 31556
rect 37202 31500 37212 31556
rect 37268 31500 37278 31556
rect 31892 31444 31948 31500
rect 26002 31388 26012 31444
rect 26068 31388 31948 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 30940 31332 30996 31388
rect 30930 31276 30940 31332
rect 30996 31276 31006 31332
rect 8754 31164 8764 31220
rect 8820 31164 11228 31220
rect 11284 31164 13804 31220
rect 13860 31164 15372 31220
rect 15428 31164 15438 31220
rect 28690 31164 28700 31220
rect 28756 31164 29708 31220
rect 29764 31164 31836 31220
rect 31892 31164 33180 31220
rect 33236 31164 34300 31220
rect 34356 31164 34366 31220
rect 7186 31052 7196 31108
rect 7252 31052 8428 31108
rect 8484 31052 9660 31108
rect 9716 31052 9726 31108
rect 16594 31052 16604 31108
rect 16660 31052 17388 31108
rect 17444 31052 17454 31108
rect 19170 31052 19180 31108
rect 19236 31052 23212 31108
rect 23268 31052 28476 31108
rect 28532 31052 28542 31108
rect 8530 30940 8540 30996
rect 8596 30940 9996 30996
rect 10052 30940 13692 30996
rect 13748 30940 13758 30996
rect 18610 30940 18620 30996
rect 18676 30940 18686 30996
rect 27794 30940 27804 30996
rect 27860 30940 31836 30996
rect 31892 30940 31902 30996
rect 32050 30940 32060 30996
rect 32116 30940 33404 30996
rect 33460 30940 35868 30996
rect 35924 30940 37772 30996
rect 37828 30940 39228 30996
rect 39284 30940 39294 30996
rect 18620 30884 18676 30940
rect 18620 30828 24108 30884
rect 24164 30828 35084 30884
rect 35140 30828 35150 30884
rect 27458 30716 27468 30772
rect 27524 30716 30268 30772
rect 30324 30716 30334 30772
rect 25778 30604 25788 30660
rect 25844 30604 31948 30660
rect 32004 30604 32014 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 3602 30380 3612 30436
rect 3668 30380 3678 30436
rect 3612 30324 3668 30380
rect 3612 30268 8372 30324
rect 8754 30268 8764 30324
rect 8820 30268 10108 30324
rect 10164 30268 10174 30324
rect 14018 30268 14028 30324
rect 14084 30268 14924 30324
rect 14980 30268 14990 30324
rect 17602 30268 17612 30324
rect 17668 30268 18396 30324
rect 18452 30268 18462 30324
rect 22642 30268 22652 30324
rect 22708 30268 23996 30324
rect 24052 30268 24062 30324
rect 28252 30268 30156 30324
rect 30212 30268 31164 30324
rect 31220 30268 31230 30324
rect 36978 30268 36988 30324
rect 37044 30268 37054 30324
rect 8316 29876 8372 30268
rect 28252 30212 28308 30268
rect 36988 30212 37044 30268
rect 9314 30156 9324 30212
rect 9380 30156 10220 30212
rect 10276 30156 10286 30212
rect 14354 30156 14364 30212
rect 14420 30156 17724 30212
rect 17780 30156 17790 30212
rect 18284 30156 18620 30212
rect 18676 30156 18686 30212
rect 20402 30156 20412 30212
rect 20468 30156 25004 30212
rect 25060 30156 25070 30212
rect 26338 30156 26348 30212
rect 26404 30156 27468 30212
rect 27524 30156 28252 30212
rect 28308 30156 28318 30212
rect 30370 30156 30380 30212
rect 30436 30156 31388 30212
rect 31444 30156 32564 30212
rect 18284 30100 18340 30156
rect 11666 30044 11676 30100
rect 11732 30044 14476 30100
rect 14532 30044 18340 30100
rect 18722 30044 18732 30100
rect 18788 30044 27356 30100
rect 27412 30044 27422 30100
rect 28466 30044 28476 30100
rect 28532 30044 31948 30100
rect 10098 29932 10108 29988
rect 10164 29932 11228 29988
rect 11284 29932 11294 29988
rect 13794 29932 13804 29988
rect 13860 29932 14252 29988
rect 14308 29932 14318 29988
rect 15092 29932 17164 29988
rect 17220 29932 17230 29988
rect 17714 29932 17724 29988
rect 17780 29932 18060 29988
rect 18116 29932 18126 29988
rect 18386 29932 18396 29988
rect 18452 29932 19068 29988
rect 19124 29932 19134 29988
rect 26226 29932 26236 29988
rect 26292 29932 26460 29988
rect 26516 29932 27132 29988
rect 27188 29932 27692 29988
rect 27748 29932 27758 29988
rect 15092 29876 15148 29932
rect 8316 29820 15148 29876
rect 16706 29820 16716 29876
rect 16772 29820 17500 29876
rect 17556 29820 17566 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 31892 29764 31948 30044
rect 32508 29988 32564 30156
rect 36428 30156 37044 30212
rect 36428 29988 36484 30156
rect 36978 30044 36988 30100
rect 37044 30044 37324 30100
rect 37380 30044 38668 30100
rect 38724 30044 38734 30100
rect 32498 29932 32508 29988
rect 32564 29932 32574 29988
rect 36418 29932 36428 29988
rect 36484 29932 36494 29988
rect 37426 29932 37436 29988
rect 37492 29932 39004 29988
rect 39060 29932 39070 29988
rect 10546 29708 10556 29764
rect 10612 29708 11564 29764
rect 11620 29708 11630 29764
rect 31892 29708 32956 29764
rect 33012 29708 33022 29764
rect 36754 29708 36764 29764
rect 36820 29708 37660 29764
rect 37716 29708 37726 29764
rect 10658 29596 10668 29652
rect 10724 29596 11340 29652
rect 11396 29596 11406 29652
rect 26786 29596 26796 29652
rect 26852 29596 27356 29652
rect 27412 29596 34188 29652
rect 34244 29596 34254 29652
rect 35746 29596 35756 29652
rect 35812 29596 36876 29652
rect 36932 29596 36942 29652
rect 6738 29484 6748 29540
rect 6804 29484 14420 29540
rect 17714 29484 17724 29540
rect 17780 29484 18172 29540
rect 18228 29484 18238 29540
rect 19170 29484 19180 29540
rect 19236 29484 26684 29540
rect 26740 29484 26750 29540
rect 27010 29484 27020 29540
rect 27076 29484 28476 29540
rect 28532 29484 28542 29540
rect 31154 29484 31164 29540
rect 31220 29484 31948 29540
rect 32004 29484 32014 29540
rect 36418 29484 36428 29540
rect 36484 29484 37996 29540
rect 38052 29484 38062 29540
rect 14364 29428 14420 29484
rect 1922 29372 1932 29428
rect 1988 29372 2828 29428
rect 2884 29372 5180 29428
rect 5236 29372 5246 29428
rect 8642 29372 8652 29428
rect 8708 29372 9884 29428
rect 9940 29372 10332 29428
rect 10388 29372 10398 29428
rect 14354 29372 14364 29428
rect 14420 29372 14430 29428
rect 20626 29372 20636 29428
rect 20692 29372 23548 29428
rect 23604 29372 23996 29428
rect 24052 29372 24062 29428
rect 26562 29372 26572 29428
rect 26628 29372 27132 29428
rect 27188 29372 27580 29428
rect 27636 29372 27646 29428
rect 4722 29260 4732 29316
rect 4788 29260 6636 29316
rect 6692 29260 6702 29316
rect 8418 29260 8428 29316
rect 8484 29260 9100 29316
rect 9156 29260 10108 29316
rect 10164 29260 10174 29316
rect 11106 29260 11116 29316
rect 11172 29260 13804 29316
rect 13860 29260 13870 29316
rect 17266 29260 17276 29316
rect 17332 29260 21196 29316
rect 21252 29260 21262 29316
rect 11666 29148 11676 29204
rect 11732 29148 13692 29204
rect 13748 29148 13758 29204
rect 31266 29148 31276 29204
rect 31332 29148 32508 29204
rect 32564 29148 32574 29204
rect 14354 29036 14364 29092
rect 14420 29036 17612 29092
rect 17668 29036 17678 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 11890 28924 11900 28980
rect 11956 28924 14588 28980
rect 14644 28924 14654 28980
rect 7970 28812 7980 28868
rect 8036 28812 8876 28868
rect 8932 28812 10724 28868
rect 10882 28812 10892 28868
rect 10948 28812 11452 28868
rect 11508 28812 11518 28868
rect 10668 28756 10724 28812
rect 8530 28700 8540 28756
rect 8596 28700 9436 28756
rect 9492 28700 9502 28756
rect 10658 28700 10668 28756
rect 10724 28700 10734 28756
rect 11218 28700 11228 28756
rect 11284 28700 12124 28756
rect 12180 28700 12190 28756
rect 21298 28700 21308 28756
rect 21364 28700 22764 28756
rect 22820 28700 22830 28756
rect 22988 28700 33404 28756
rect 33460 28700 33470 28756
rect 22988 28644 23044 28700
rect 8754 28588 8764 28644
rect 8820 28588 9548 28644
rect 9604 28588 10220 28644
rect 10276 28588 10286 28644
rect 12002 28588 12012 28644
rect 12068 28588 13468 28644
rect 13524 28588 13534 28644
rect 13906 28588 13916 28644
rect 13972 28588 14700 28644
rect 14756 28588 14766 28644
rect 20178 28588 20188 28644
rect 20244 28588 20748 28644
rect 20804 28588 23044 28644
rect 25890 28588 25900 28644
rect 25956 28588 26572 28644
rect 26628 28588 26638 28644
rect 28018 28588 28028 28644
rect 28084 28588 28364 28644
rect 28420 28588 28430 28644
rect 20188 28532 20244 28588
rect 9426 28476 9436 28532
rect 9492 28476 10332 28532
rect 10388 28476 10398 28532
rect 12338 28476 12348 28532
rect 12404 28476 13804 28532
rect 13860 28476 13870 28532
rect 15362 28476 15372 28532
rect 15428 28476 20244 28532
rect 21746 28476 21756 28532
rect 21812 28476 23772 28532
rect 23828 28476 23838 28532
rect 27458 28476 27468 28532
rect 27524 28476 28140 28532
rect 28196 28476 28206 28532
rect 28690 28476 28700 28532
rect 28756 28476 29708 28532
rect 29764 28476 29774 28532
rect 36306 28476 36316 28532
rect 36372 28476 37660 28532
rect 37716 28476 37726 28532
rect 10882 28364 10892 28420
rect 10948 28364 13468 28420
rect 13524 28364 13534 28420
rect 26898 28364 26908 28420
rect 26964 28364 28588 28420
rect 28644 28364 30044 28420
rect 30100 28364 30492 28420
rect 30548 28364 30558 28420
rect 32610 28364 32620 28420
rect 32676 28364 33964 28420
rect 34020 28364 34030 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 22866 28140 22876 28196
rect 22932 28140 22942 28196
rect 22876 28084 22932 28140
rect 8418 28028 8428 28084
rect 8484 28028 8988 28084
rect 9044 28028 17948 28084
rect 18004 28028 18014 28084
rect 22642 28028 22652 28084
rect 22708 28028 22932 28084
rect 21634 27916 21644 27972
rect 21700 27916 23100 27972
rect 23156 27916 30268 27972
rect 30324 27916 30334 27972
rect 32834 27916 32844 27972
rect 32900 27916 33628 27972
rect 33684 27916 37100 27972
rect 37156 27916 38556 27972
rect 38612 27916 38622 27972
rect 9202 27804 9212 27860
rect 9268 27804 10444 27860
rect 10500 27804 10510 27860
rect 26898 27804 26908 27860
rect 26964 27804 28252 27860
rect 28308 27804 29148 27860
rect 29204 27804 29214 27860
rect 6738 27692 6748 27748
rect 6804 27692 9436 27748
rect 9492 27692 9502 27748
rect 38098 27692 38108 27748
rect 38164 27692 39228 27748
rect 39284 27692 39294 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 15362 27356 15372 27412
rect 15428 27356 16716 27412
rect 16772 27356 16782 27412
rect 30034 27244 30044 27300
rect 30100 27244 35980 27300
rect 36036 27244 39004 27300
rect 39060 27244 39070 27300
rect 9762 27132 9772 27188
rect 9828 27132 10444 27188
rect 10500 27132 12236 27188
rect 12292 27132 12302 27188
rect 28130 27132 28140 27188
rect 28196 27132 29372 27188
rect 29428 27132 29438 27188
rect 35186 27132 35196 27188
rect 35252 27132 35756 27188
rect 35812 27132 35822 27188
rect 25666 27020 25676 27076
rect 25732 27020 26236 27076
rect 26292 27020 26796 27076
rect 26852 27020 26862 27076
rect 36082 27020 36092 27076
rect 36148 27020 38332 27076
rect 38388 27020 38398 27076
rect 1810 26908 1820 26964
rect 1876 26908 3836 26964
rect 3892 26908 5068 26964
rect 5124 26908 7196 26964
rect 7252 26908 7262 26964
rect 12450 26908 12460 26964
rect 12516 26908 14252 26964
rect 14308 26908 14812 26964
rect 14868 26908 14878 26964
rect 31938 26908 31948 26964
rect 32004 26908 34748 26964
rect 34804 26908 35756 26964
rect 35812 26908 35822 26964
rect 36194 26908 36204 26964
rect 36260 26908 36988 26964
rect 37044 26908 37054 26964
rect 35522 26796 35532 26852
rect 35588 26796 36428 26852
rect 36484 26796 36494 26852
rect 37426 26796 37436 26852
rect 37492 26796 38332 26852
rect 38388 26796 38398 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 6850 26572 6860 26628
rect 6916 26572 7532 26628
rect 7588 26572 7598 26628
rect 26562 26572 26572 26628
rect 26628 26572 27468 26628
rect 27524 26572 27804 26628
rect 27860 26572 27870 26628
rect 18274 26460 18284 26516
rect 18340 26460 34636 26516
rect 34692 26460 34702 26516
rect 4610 26236 4620 26292
rect 4676 26236 6412 26292
rect 6468 26236 6478 26292
rect 26226 26236 26236 26292
rect 26292 26236 27020 26292
rect 27076 26236 27086 26292
rect 35858 26236 35868 26292
rect 35924 26236 36764 26292
rect 36820 26236 36830 26292
rect 13010 26124 13020 26180
rect 13076 26124 15484 26180
rect 15540 26124 17500 26180
rect 17556 26124 17566 26180
rect 18834 26124 18844 26180
rect 18900 26124 20748 26180
rect 20804 26124 20814 26180
rect 22866 26124 22876 26180
rect 22932 26124 25228 26180
rect 25284 26124 25294 26180
rect 26684 26012 28252 26068
rect 28308 26012 28318 26068
rect 26684 25956 26740 26012
rect 26674 25900 26684 25956
rect 26740 25900 26750 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 17490 25788 17500 25844
rect 17556 25788 23100 25844
rect 23156 25788 26908 25844
rect 26964 25788 26974 25844
rect 28242 25788 28252 25844
rect 28308 25788 29484 25844
rect 29540 25788 30716 25844
rect 30772 25788 30782 25844
rect 14018 25564 14028 25620
rect 14084 25564 15596 25620
rect 15652 25564 15662 25620
rect 20738 25564 20748 25620
rect 20804 25564 25452 25620
rect 25508 25564 25518 25620
rect 6402 25452 6412 25508
rect 6468 25452 7308 25508
rect 7364 25452 7374 25508
rect 25778 25452 25788 25508
rect 25844 25452 34076 25508
rect 34132 25452 34142 25508
rect 16258 25228 16268 25284
rect 16324 25228 16828 25284
rect 16884 25228 17500 25284
rect 17556 25228 17948 25284
rect 18004 25228 18014 25284
rect 27346 25116 27356 25172
rect 27412 25116 29148 25172
rect 29204 25116 32172 25172
rect 32228 25116 32238 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 28130 25004 28140 25060
rect 28196 25004 28924 25060
rect 28980 25004 28990 25060
rect 5730 24892 5740 24948
rect 5796 24892 7868 24948
rect 7924 24892 7934 24948
rect 4946 24780 4956 24836
rect 5012 24780 5964 24836
rect 6020 24780 6030 24836
rect 28354 24780 28364 24836
rect 28420 24780 29372 24836
rect 29428 24780 29438 24836
rect 35634 24780 35644 24836
rect 35700 24780 36428 24836
rect 36484 24780 36494 24836
rect 3490 24668 3500 24724
rect 3556 24668 6524 24724
rect 6580 24668 6590 24724
rect 6962 24668 6972 24724
rect 7028 24668 7644 24724
rect 7700 24668 7710 24724
rect 18834 24668 18844 24724
rect 18900 24668 19292 24724
rect 19348 24668 22428 24724
rect 22484 24668 22494 24724
rect 24658 24668 24668 24724
rect 24724 24668 25564 24724
rect 25620 24668 25630 24724
rect 26226 24668 26236 24724
rect 26292 24668 28588 24724
rect 28644 24668 29708 24724
rect 29764 24668 29774 24724
rect 36082 24668 36092 24724
rect 36148 24668 37100 24724
rect 37156 24668 37166 24724
rect 7186 24556 7196 24612
rect 7252 24556 8316 24612
rect 8372 24556 8382 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 24546 24108 24556 24164
rect 24612 24108 25564 24164
rect 25620 24108 26012 24164
rect 26068 24108 26078 24164
rect 35970 24108 35980 24164
rect 36036 24108 37156 24164
rect 37100 24052 37156 24108
rect 12786 23996 12796 24052
rect 12852 23996 13804 24052
rect 13860 23996 13870 24052
rect 35186 23996 35196 24052
rect 35252 23996 36092 24052
rect 36148 23996 36158 24052
rect 37090 23996 37100 24052
rect 37156 23996 38108 24052
rect 38164 23996 38174 24052
rect 3266 23884 3276 23940
rect 3332 23884 4396 23940
rect 4452 23884 4462 23940
rect 4834 23884 4844 23940
rect 4900 23884 5628 23940
rect 5684 23884 5694 23940
rect 8418 23884 8428 23940
rect 8484 23884 11900 23940
rect 11956 23884 15148 23940
rect 15204 23884 15214 23940
rect 20290 23884 20300 23940
rect 20356 23884 21756 23940
rect 21812 23884 23548 23940
rect 23604 23884 25004 23940
rect 25060 23884 31948 23940
rect 32004 23884 32284 23940
rect 32340 23884 32844 23940
rect 32900 23884 32910 23940
rect 35858 23884 35868 23940
rect 35924 23884 37436 23940
rect 37492 23884 38668 23940
rect 38612 23828 38668 23884
rect 21634 23772 21644 23828
rect 21700 23772 22428 23828
rect 22484 23772 22494 23828
rect 26898 23772 26908 23828
rect 26964 23772 27132 23828
rect 27188 23772 27198 23828
rect 31490 23772 31500 23828
rect 31556 23772 33068 23828
rect 33124 23772 33134 23828
rect 36418 23772 36428 23828
rect 36484 23772 37548 23828
rect 37604 23772 37614 23828
rect 38612 23772 38892 23828
rect 38948 23772 38958 23828
rect 12898 23660 12908 23716
rect 12964 23660 13916 23716
rect 13972 23660 13982 23716
rect 19506 23548 19516 23604
rect 19572 23548 19582 23604
rect 7074 23436 7084 23492
rect 7140 23436 7980 23492
rect 8036 23436 8046 23492
rect 19516 23380 19572 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 31266 23436 31276 23492
rect 31332 23436 37772 23492
rect 37828 23436 37838 23492
rect 17042 23324 17052 23380
rect 17108 23324 17500 23380
rect 17556 23324 17566 23380
rect 18162 23324 18172 23380
rect 18228 23324 23660 23380
rect 23716 23324 23726 23380
rect 31276 23268 31332 23436
rect 14018 23212 14028 23268
rect 14084 23212 15596 23268
rect 15652 23212 15662 23268
rect 17602 23212 17612 23268
rect 17668 23212 26908 23268
rect 26964 23212 26974 23268
rect 31042 23212 31052 23268
rect 31108 23212 31332 23268
rect 36418 23212 36428 23268
rect 36484 23212 37100 23268
rect 37156 23212 37166 23268
rect 6066 23100 6076 23156
rect 6132 23100 7980 23156
rect 8036 23100 8046 23156
rect 18498 23100 18508 23156
rect 18564 23100 19180 23156
rect 19236 23100 19246 23156
rect 21970 23100 21980 23156
rect 22036 23100 22764 23156
rect 22820 23100 22830 23156
rect 22978 23100 22988 23156
rect 23044 23100 23436 23156
rect 23492 23100 23502 23156
rect 29922 23100 29932 23156
rect 29988 23100 31164 23156
rect 31220 23100 31230 23156
rect 36754 23100 36764 23156
rect 36820 23100 37324 23156
rect 37380 23100 37390 23156
rect 22764 23044 22820 23100
rect 7746 22988 7756 23044
rect 7812 22988 10332 23044
rect 10388 22988 10398 23044
rect 19506 22988 19516 23044
rect 19572 22988 19964 23044
rect 20020 22988 20412 23044
rect 20468 22988 22092 23044
rect 22148 22988 22158 23044
rect 22764 22988 23884 23044
rect 23940 22988 23950 23044
rect 28466 22988 28476 23044
rect 28532 22988 30268 23044
rect 30324 22988 30334 23044
rect 32274 22988 32284 23044
rect 32340 22988 34076 23044
rect 34132 22988 34142 23044
rect 3490 22876 3500 22932
rect 3556 22876 8316 22932
rect 8372 22876 11564 22932
rect 11620 22876 11630 22932
rect 14802 22876 14812 22932
rect 14868 22876 16828 22932
rect 16884 22876 17948 22932
rect 18004 22876 18396 22932
rect 18452 22876 18462 22932
rect 22530 22876 22540 22932
rect 22596 22876 26908 22932
rect 27682 22876 27692 22932
rect 27748 22876 30492 22932
rect 30548 22876 31612 22932
rect 31668 22876 31678 22932
rect 26852 22820 26908 22876
rect 15092 22764 15932 22820
rect 15988 22764 17388 22820
rect 17444 22764 17454 22820
rect 26852 22764 30380 22820
rect 30436 22764 30446 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 8166 22652 8204 22708
rect 8260 22652 8270 22708
rect 15092 22596 15148 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 7186 22540 7196 22596
rect 7252 22540 7756 22596
rect 7812 22540 7822 22596
rect 14018 22540 14028 22596
rect 14084 22540 15148 22596
rect 30482 22540 30492 22596
rect 30548 22540 31052 22596
rect 31108 22540 31118 22596
rect 37762 22540 37772 22596
rect 37828 22540 39116 22596
rect 39172 22540 39182 22596
rect 5842 22428 5852 22484
rect 5908 22428 6300 22484
rect 6356 22428 8204 22484
rect 8260 22428 8270 22484
rect 15250 22428 15260 22484
rect 15316 22428 16156 22484
rect 16212 22428 16222 22484
rect 16930 22428 16940 22484
rect 16996 22428 18172 22484
rect 18228 22428 18238 22484
rect 35746 22428 35756 22484
rect 35812 22428 36428 22484
rect 36484 22428 36494 22484
rect 16940 22372 16996 22428
rect 5954 22316 5964 22372
rect 6020 22316 6748 22372
rect 6804 22316 6814 22372
rect 9874 22316 9884 22372
rect 9940 22316 12460 22372
rect 12516 22316 15708 22372
rect 15764 22316 15774 22372
rect 16034 22316 16044 22372
rect 16100 22316 16996 22372
rect 18274 22316 18284 22372
rect 18340 22316 18956 22372
rect 19012 22316 19022 22372
rect 29250 22316 29260 22372
rect 29316 22316 30044 22372
rect 30100 22316 30110 22372
rect 36082 22316 36092 22372
rect 36148 22316 37436 22372
rect 37492 22316 37502 22372
rect 7074 22204 7084 22260
rect 7140 22204 9996 22260
rect 10052 22204 10062 22260
rect 10770 22204 10780 22260
rect 10836 22204 12796 22260
rect 12852 22204 13356 22260
rect 13412 22204 13422 22260
rect 14578 22204 14588 22260
rect 14644 22204 15596 22260
rect 15652 22204 15662 22260
rect 19058 22204 19068 22260
rect 19124 22204 19628 22260
rect 19684 22204 20412 22260
rect 20468 22204 20478 22260
rect 30940 22204 31948 22260
rect 32004 22204 32014 22260
rect 5058 22092 5068 22148
rect 5124 22092 5852 22148
rect 5908 22092 5918 22148
rect 7298 22092 7308 22148
rect 7364 22092 14140 22148
rect 14196 22092 14700 22148
rect 14756 22092 14766 22148
rect 15092 22092 18956 22148
rect 19012 22092 19022 22148
rect 28242 22092 28252 22148
rect 28308 22092 29708 22148
rect 29764 22092 29774 22148
rect 15092 22036 15148 22092
rect 30940 22036 30996 22204
rect 31826 22092 31836 22148
rect 31892 22092 35532 22148
rect 35588 22092 35598 22148
rect 9202 21980 9212 22036
rect 9268 21980 9548 22036
rect 9604 21980 9614 22036
rect 11442 21980 11452 22036
rect 11508 21980 15148 22036
rect 18722 21980 18732 22036
rect 18788 21980 19628 22036
rect 19684 21980 19694 22036
rect 23426 21980 23436 22036
rect 23492 21980 28700 22036
rect 28756 21980 30940 22036
rect 30996 21980 31006 22036
rect 31378 21980 31388 22036
rect 31444 21980 31724 22036
rect 31780 21980 32060 22036
rect 32116 21980 36092 22036
rect 36148 21980 36158 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 6850 21868 6860 21924
rect 6916 21868 12516 21924
rect 29474 21868 29484 21924
rect 29540 21868 30380 21924
rect 30436 21868 31500 21924
rect 31556 21868 31566 21924
rect 31826 21868 31836 21924
rect 31892 21868 32508 21924
rect 32564 21868 32574 21924
rect 10434 21756 10444 21812
rect 10500 21756 11340 21812
rect 11396 21756 11406 21812
rect 7970 21644 7980 21700
rect 8036 21644 8764 21700
rect 8820 21644 9548 21700
rect 9604 21644 9614 21700
rect 3714 21532 3724 21588
rect 3780 21532 5068 21588
rect 5124 21532 7084 21588
rect 7140 21532 7150 21588
rect 12460 21476 12516 21868
rect 14354 21756 14364 21812
rect 14420 21756 27692 21812
rect 27748 21756 29372 21812
rect 29428 21756 29932 21812
rect 29988 21756 29998 21812
rect 14466 21644 14476 21700
rect 14532 21644 15652 21700
rect 31714 21644 31724 21700
rect 31780 21644 33180 21700
rect 33236 21644 33246 21700
rect 12674 21532 12684 21588
rect 12740 21532 13468 21588
rect 13524 21532 14588 21588
rect 14644 21532 14654 21588
rect 15596 21476 15652 21644
rect 19058 21532 19068 21588
rect 19124 21532 20076 21588
rect 20132 21532 25900 21588
rect 25956 21532 32508 21588
rect 32564 21532 32574 21588
rect 12460 21420 14028 21476
rect 14084 21420 14094 21476
rect 15586 21420 15596 21476
rect 15652 21420 15662 21476
rect 18722 21420 18732 21476
rect 18788 21420 19964 21476
rect 20020 21420 20030 21476
rect 27010 21420 27020 21476
rect 27076 21420 30492 21476
rect 30548 21420 36428 21476
rect 36484 21420 36494 21476
rect 38882 21420 38892 21476
rect 38948 21420 39564 21476
rect 39620 21420 39630 21476
rect 4946 21308 4956 21364
rect 5012 21308 5404 21364
rect 5460 21308 7644 21364
rect 7700 21308 8540 21364
rect 8596 21308 8606 21364
rect 25218 21308 25228 21364
rect 25284 21308 25676 21364
rect 25732 21308 25742 21364
rect 31826 21308 31836 21364
rect 31892 21308 35868 21364
rect 35924 21308 35934 21364
rect 14914 21196 14924 21252
rect 14980 21196 28028 21252
rect 28084 21196 28094 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 15138 21084 15148 21140
rect 15204 21084 26124 21140
rect 26180 21084 28140 21140
rect 28196 21084 28206 21140
rect 8866 20972 8876 21028
rect 8932 20972 9548 21028
rect 9604 20972 9772 21028
rect 9828 20972 9838 21028
rect 7410 20860 7420 20916
rect 7476 20860 10500 20916
rect 10444 20804 10500 20860
rect 7746 20748 7756 20804
rect 7812 20748 8652 20804
rect 8708 20748 8718 20804
rect 10434 20748 10444 20804
rect 10500 20748 12908 20804
rect 12964 20748 12974 20804
rect 22866 20748 22876 20804
rect 22932 20748 26796 20804
rect 26852 20748 26862 20804
rect 5506 20636 5516 20692
rect 5572 20636 8316 20692
rect 8372 20636 8382 20692
rect 26002 20636 26012 20692
rect 26068 20636 27580 20692
rect 27636 20636 28252 20692
rect 28308 20636 28318 20692
rect 26012 20580 26068 20636
rect 6402 20524 6412 20580
rect 6468 20524 7084 20580
rect 7140 20524 7150 20580
rect 10322 20524 10332 20580
rect 10388 20524 18844 20580
rect 18900 20524 18910 20580
rect 25218 20524 25228 20580
rect 25284 20524 26068 20580
rect 27906 20524 27916 20580
rect 27972 20524 30492 20580
rect 30548 20524 31164 20580
rect 31220 20524 31230 20580
rect 33730 20524 33740 20580
rect 33796 20524 37100 20580
rect 37156 20524 37772 20580
rect 37828 20524 38556 20580
rect 38612 20524 38622 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 21634 20300 21644 20356
rect 21700 20300 25452 20356
rect 25508 20300 25900 20356
rect 25956 20300 25966 20356
rect 8754 20188 8764 20244
rect 8820 20188 9772 20244
rect 9828 20188 9838 20244
rect 19058 20188 19068 20244
rect 19124 20188 19740 20244
rect 19796 20188 19806 20244
rect 25330 20188 25340 20244
rect 25396 20188 25406 20244
rect 26898 20188 26908 20244
rect 26964 20188 27300 20244
rect 28130 20188 28140 20244
rect 28196 20188 29820 20244
rect 29876 20188 29886 20244
rect 30706 20188 30716 20244
rect 30772 20188 30782 20244
rect 25340 20132 25396 20188
rect 27244 20132 27300 20188
rect 30716 20132 30772 20188
rect 3938 20076 3948 20132
rect 4004 20076 5628 20132
rect 5684 20076 8204 20132
rect 8260 20076 8270 20132
rect 10770 20076 10780 20132
rect 10836 20076 11340 20132
rect 11396 20076 11676 20132
rect 11732 20076 11742 20132
rect 13794 20076 13804 20132
rect 13860 20076 14924 20132
rect 14980 20076 14990 20132
rect 15138 20076 15148 20132
rect 15204 20076 15932 20132
rect 15988 20076 16380 20132
rect 16436 20076 17052 20132
rect 17108 20076 17388 20132
rect 17444 20076 17454 20132
rect 20514 20076 20524 20132
rect 20580 20076 22652 20132
rect 22708 20076 23772 20132
rect 23828 20076 23838 20132
rect 25340 20076 26124 20132
rect 26180 20076 27020 20132
rect 27076 20076 27086 20132
rect 27244 20076 35756 20132
rect 35812 20076 35822 20132
rect 5058 19964 5068 20020
rect 5124 19964 6524 20020
rect 6580 19964 6590 20020
rect 11554 19964 11564 20020
rect 11620 19964 13356 20020
rect 13412 19964 15540 20020
rect 16706 19964 16716 20020
rect 16772 19964 19292 20020
rect 19348 19964 19628 20020
rect 19684 19964 19694 20020
rect 23090 19964 23100 20020
rect 23156 19964 24276 20020
rect 24434 19964 24444 20020
rect 24500 19964 26684 20020
rect 26740 19964 26750 20020
rect 28018 19964 28028 20020
rect 28084 19964 28588 20020
rect 28644 19964 28654 20020
rect 12450 19852 12460 19908
rect 12516 19852 13692 19908
rect 13748 19852 13758 19908
rect 15484 19796 15540 19964
rect 24220 19908 24276 19964
rect 18386 19852 18396 19908
rect 18452 19852 21196 19908
rect 21252 19852 21644 19908
rect 21700 19852 21710 19908
rect 21858 19852 21868 19908
rect 21924 19852 23996 19908
rect 24052 19852 24062 19908
rect 24210 19852 24220 19908
rect 24276 19852 35980 19908
rect 36036 19852 37548 19908
rect 37604 19852 37614 19908
rect 15474 19740 15484 19796
rect 15540 19740 15550 19796
rect 20626 19628 20636 19684
rect 20692 19628 31276 19684
rect 31332 19628 31342 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 9426 19516 9436 19572
rect 9492 19516 9502 19572
rect 9436 19236 9492 19516
rect 14802 19404 14812 19460
rect 14868 19404 15932 19460
rect 15988 19404 21868 19460
rect 21924 19404 21934 19460
rect 23650 19404 23660 19460
rect 23716 19404 31164 19460
rect 31220 19404 31230 19460
rect 31490 19404 31500 19460
rect 31556 19404 33404 19460
rect 33460 19404 33470 19460
rect 13570 19292 13580 19348
rect 13636 19292 14588 19348
rect 14644 19292 14654 19348
rect 18834 19292 18844 19348
rect 18900 19292 25228 19348
rect 25284 19292 25294 19348
rect 37538 19292 37548 19348
rect 37604 19292 38332 19348
rect 38388 19292 38398 19348
rect 4722 19180 4732 19236
rect 4788 19180 6188 19236
rect 6244 19180 7756 19236
rect 7812 19180 7822 19236
rect 8418 19180 8428 19236
rect 8484 19180 11116 19236
rect 11172 19180 11182 19236
rect 19506 19180 19516 19236
rect 19572 19180 21308 19236
rect 21364 19180 21374 19236
rect 25442 19180 25452 19236
rect 25508 19180 26684 19236
rect 26740 19180 26750 19236
rect 32050 19180 32060 19236
rect 32116 19180 33404 19236
rect 33460 19180 33470 19236
rect 2482 19068 2492 19124
rect 2548 19068 3500 19124
rect 3556 19068 3566 19124
rect 8194 19068 8204 19124
rect 8260 19068 9212 19124
rect 9268 19068 10220 19124
rect 10276 19068 10286 19124
rect 19618 19068 19628 19124
rect 19684 19068 20076 19124
rect 20132 19068 21644 19124
rect 21700 19068 21710 19124
rect 36194 19068 36204 19124
rect 36260 19068 37324 19124
rect 37380 19068 37390 19124
rect 15474 18956 15484 19012
rect 15540 18956 18956 19012
rect 19012 18956 20188 19012
rect 20244 18956 20254 19012
rect 27234 18956 27244 19012
rect 27300 18956 27692 19012
rect 27748 18956 28028 19012
rect 28084 18956 28094 19012
rect 3602 18844 3612 18900
rect 3668 18844 4396 18900
rect 4452 18844 16716 18900
rect 16772 18844 16782 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 21858 18732 21868 18788
rect 21924 18732 23212 18788
rect 23268 18732 23278 18788
rect 27122 18732 27132 18788
rect 27188 18732 31612 18788
rect 31668 18732 31678 18788
rect 18274 18620 18284 18676
rect 18340 18620 18844 18676
rect 18900 18620 18910 18676
rect 19842 18620 19852 18676
rect 19908 18620 21532 18676
rect 21588 18620 27468 18676
rect 27524 18620 27534 18676
rect 5058 18508 5068 18564
rect 5124 18508 5964 18564
rect 6020 18508 6030 18564
rect 17378 18508 17388 18564
rect 17444 18508 23548 18564
rect 23604 18508 24556 18564
rect 24612 18508 24622 18564
rect 37314 18508 37324 18564
rect 37380 18508 38108 18564
rect 38164 18508 38174 18564
rect 12786 18396 12796 18452
rect 12852 18396 17780 18452
rect 17938 18396 17948 18452
rect 18004 18396 18508 18452
rect 18564 18396 19292 18452
rect 19348 18396 19358 18452
rect 32274 18396 32284 18452
rect 32340 18396 33068 18452
rect 33124 18396 33134 18452
rect 36306 18396 36316 18452
rect 36372 18396 38220 18452
rect 38276 18396 38286 18452
rect 17724 18340 17780 18396
rect 17724 18284 19628 18340
rect 19684 18284 19694 18340
rect 26450 18284 26460 18340
rect 26516 18284 26796 18340
rect 26852 18284 31892 18340
rect 33954 18284 33964 18340
rect 34020 18284 35980 18340
rect 36036 18284 36046 18340
rect 37090 18284 37100 18340
rect 37156 18284 37166 18340
rect 31836 18228 31892 18284
rect 37100 18228 37156 18284
rect 14802 18172 14812 18228
rect 14868 18172 19068 18228
rect 19124 18172 19740 18228
rect 19796 18172 19806 18228
rect 26852 18172 31612 18228
rect 31668 18172 31678 18228
rect 31836 18172 37156 18228
rect 26852 18116 26908 18172
rect 16594 18060 16604 18116
rect 16660 18060 26908 18116
rect 36082 18060 36092 18116
rect 36148 18060 37212 18116
rect 37268 18060 37436 18116
rect 37492 18060 37502 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 11778 17948 11788 18004
rect 11844 17948 21868 18004
rect 21924 17948 21934 18004
rect 11666 17836 11676 17892
rect 11732 17836 17276 17892
rect 17332 17836 17342 17892
rect 22866 17836 22876 17892
rect 22932 17836 23772 17892
rect 23828 17836 26572 17892
rect 26628 17836 26638 17892
rect 36530 17836 36540 17892
rect 36596 17836 37212 17892
rect 37268 17836 37278 17892
rect 4610 17724 4620 17780
rect 4676 17724 5796 17780
rect 18386 17724 18396 17780
rect 18452 17724 18732 17780
rect 18788 17724 19740 17780
rect 19796 17724 19806 17780
rect 33282 17724 33292 17780
rect 33348 17724 37100 17780
rect 37156 17724 37166 17780
rect 5740 17668 5796 17724
rect 1810 17612 1820 17668
rect 1876 17612 5068 17668
rect 5124 17612 5134 17668
rect 5730 17612 5740 17668
rect 5796 17612 8540 17668
rect 8596 17612 8606 17668
rect 19618 17612 19628 17668
rect 19684 17612 22540 17668
rect 22596 17612 23100 17668
rect 23156 17612 23166 17668
rect 37202 17612 37212 17668
rect 37268 17612 38052 17668
rect 37996 17556 38052 17612
rect 7634 17500 7644 17556
rect 7700 17500 8428 17556
rect 8484 17500 8494 17556
rect 23426 17500 23436 17556
rect 23492 17500 24332 17556
rect 24388 17500 24398 17556
rect 37986 17500 37996 17556
rect 38052 17500 38062 17556
rect 24434 17388 24444 17444
rect 24500 17388 27468 17444
rect 27524 17388 27534 17444
rect 35746 17388 35756 17444
rect 35812 17388 37660 17444
rect 37716 17388 37726 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 23202 17164 23212 17220
rect 23268 17164 23278 17220
rect 23212 17108 23268 17164
rect 10434 17052 10444 17108
rect 10500 17052 11676 17108
rect 11732 17052 11742 17108
rect 17826 17052 17836 17108
rect 17892 17052 18844 17108
rect 18900 17052 18910 17108
rect 22866 17052 22876 17108
rect 22932 17052 23268 17108
rect 24882 17052 24892 17108
rect 24948 17052 29932 17108
rect 29988 17052 30716 17108
rect 30772 17052 30782 17108
rect 31714 17052 31724 17108
rect 31780 17052 32060 17108
rect 32116 17052 32126 17108
rect 23212 16996 23268 17052
rect 23212 16940 23548 16996
rect 23604 16940 25228 16996
rect 25284 16940 25294 16996
rect 30034 16940 30044 16996
rect 30100 16940 30940 16996
rect 30996 16940 33292 16996
rect 33348 16940 33358 16996
rect 1922 16828 1932 16884
rect 1988 16828 10332 16884
rect 10388 16828 10398 16884
rect 17378 16828 17388 16884
rect 17444 16828 17836 16884
rect 17892 16828 17902 16884
rect 18162 16828 18172 16884
rect 18228 16828 19292 16884
rect 19348 16828 19358 16884
rect 24098 16828 24108 16884
rect 24164 16828 24174 16884
rect 24546 16828 24556 16884
rect 24612 16828 25620 16884
rect 26786 16828 26796 16884
rect 26852 16828 30380 16884
rect 30436 16828 31164 16884
rect 31220 16828 31230 16884
rect 32284 16828 35308 16884
rect 35364 16828 35374 16884
rect 3042 16716 3052 16772
rect 3108 16716 4172 16772
rect 4228 16716 5852 16772
rect 5908 16716 7308 16772
rect 7364 16716 7374 16772
rect 7746 16716 7756 16772
rect 7812 16716 12236 16772
rect 12292 16716 12302 16772
rect 18172 16660 18228 16828
rect 24108 16772 24164 16828
rect 25564 16772 25620 16828
rect 22530 16716 22540 16772
rect 22596 16716 24164 16772
rect 25554 16716 25564 16772
rect 25620 16716 29596 16772
rect 29652 16716 31388 16772
rect 31444 16716 31454 16772
rect 32284 16660 32340 16828
rect 35858 16716 35868 16772
rect 35924 16716 37212 16772
rect 37268 16716 37278 16772
rect 9874 16604 9884 16660
rect 9940 16604 10892 16660
rect 10948 16604 10958 16660
rect 12562 16604 12572 16660
rect 12628 16604 18228 16660
rect 32274 16604 32284 16660
rect 32340 16604 32350 16660
rect 20738 16492 20748 16548
rect 20804 16492 27244 16548
rect 27300 16492 31612 16548
rect 31668 16492 33628 16548
rect 33684 16492 33694 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 18162 16380 18172 16436
rect 18228 16380 22092 16436
rect 22148 16380 22158 16436
rect 6066 16268 6076 16324
rect 6132 16268 6972 16324
rect 7028 16268 7038 16324
rect 7634 16268 7644 16324
rect 7700 16268 18508 16324
rect 18564 16268 18574 16324
rect 19282 16268 19292 16324
rect 19348 16268 19852 16324
rect 19908 16268 24668 16324
rect 24724 16268 24734 16324
rect 31826 16268 31836 16324
rect 31892 16268 34636 16324
rect 34692 16268 35532 16324
rect 35588 16268 35598 16324
rect 9762 16156 9772 16212
rect 9828 16156 10444 16212
rect 10500 16156 11788 16212
rect 11844 16156 11854 16212
rect 14354 16156 14364 16212
rect 14420 16156 15708 16212
rect 15764 16156 15774 16212
rect 18162 16156 18172 16212
rect 18228 16156 18620 16212
rect 18676 16156 20188 16212
rect 20244 16156 30156 16212
rect 30212 16156 30222 16212
rect 31378 16156 31388 16212
rect 31444 16156 37492 16212
rect 37436 16100 37492 16156
rect 15250 16044 15260 16100
rect 15316 16044 22540 16100
rect 22596 16044 22606 16100
rect 23762 16044 23772 16100
rect 23828 16044 26684 16100
rect 26740 16044 26750 16100
rect 31154 16044 31164 16100
rect 31220 16044 34412 16100
rect 34468 16044 36316 16100
rect 36372 16044 36382 16100
rect 37426 16044 37436 16100
rect 37492 16044 37502 16100
rect 14578 15932 14588 15988
rect 14644 15932 17836 15988
rect 17892 15932 17902 15988
rect 18946 15932 18956 15988
rect 19012 15932 22204 15988
rect 22260 15932 22270 15988
rect 22418 15932 22428 15988
rect 22484 15932 23324 15988
rect 23380 15932 27244 15988
rect 27300 15932 27804 15988
rect 27860 15932 27870 15988
rect 32610 15932 32620 15988
rect 32676 15932 33404 15988
rect 33460 15932 34860 15988
rect 34916 15932 34926 15988
rect 35186 15932 35196 15988
rect 35252 15932 35868 15988
rect 35924 15932 35934 15988
rect 3266 15820 3276 15876
rect 3332 15820 4060 15876
rect 4116 15820 4126 15876
rect 4274 15820 4284 15876
rect 4340 15820 4956 15876
rect 5012 15820 5022 15876
rect 6178 15820 6188 15876
rect 6244 15820 7420 15876
rect 7476 15820 7486 15876
rect 12674 15820 12684 15876
rect 12740 15820 14924 15876
rect 14980 15820 14990 15876
rect 17714 15820 17724 15876
rect 17780 15820 19404 15876
rect 19460 15820 22876 15876
rect 22932 15820 22942 15876
rect 23090 15820 23100 15876
rect 23156 15820 23436 15876
rect 23492 15820 23996 15876
rect 24052 15820 24062 15876
rect 27346 15820 27356 15876
rect 27412 15820 28028 15876
rect 28084 15820 29484 15876
rect 29540 15820 29932 15876
rect 29988 15820 29998 15876
rect 18386 15708 18396 15764
rect 18452 15708 18676 15764
rect 18620 15652 18676 15708
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 18610 15596 18620 15652
rect 18676 15596 18686 15652
rect 4946 15484 4956 15540
rect 5012 15484 6076 15540
rect 6132 15484 6142 15540
rect 7298 15484 7308 15540
rect 7364 15484 10220 15540
rect 10276 15484 10286 15540
rect 19058 15484 19068 15540
rect 19124 15484 20076 15540
rect 20132 15484 20142 15540
rect 22194 15484 22204 15540
rect 22260 15484 23100 15540
rect 23156 15484 23772 15540
rect 23828 15484 23838 15540
rect 30482 15484 30492 15540
rect 30548 15484 31388 15540
rect 31444 15484 31948 15540
rect 32004 15484 32014 15540
rect 5058 15372 5068 15428
rect 5124 15372 5628 15428
rect 5684 15372 5694 15428
rect 8978 15372 8988 15428
rect 9044 15372 10332 15428
rect 10388 15372 10398 15428
rect 18498 15372 18508 15428
rect 18564 15372 19740 15428
rect 19796 15372 19806 15428
rect 30146 15372 30156 15428
rect 30212 15372 31052 15428
rect 31108 15372 32788 15428
rect 5068 15316 5124 15372
rect 2818 15260 2828 15316
rect 2884 15260 3500 15316
rect 3556 15260 3566 15316
rect 4386 15260 4396 15316
rect 4452 15260 5124 15316
rect 6850 15260 6860 15316
rect 6916 15260 9212 15316
rect 9268 15260 9278 15316
rect 18844 15260 19404 15316
rect 19460 15260 20300 15316
rect 20356 15260 20366 15316
rect 23874 15260 23884 15316
rect 23940 15260 24668 15316
rect 24724 15260 24734 15316
rect 29922 15260 29932 15316
rect 29988 15260 30268 15316
rect 30324 15260 31780 15316
rect 4050 15148 4060 15204
rect 4116 15148 5292 15204
rect 5348 15148 5852 15204
rect 5908 15148 6524 15204
rect 6580 15148 6590 15204
rect 6860 15148 7196 15204
rect 7252 15148 7262 15204
rect 10098 15148 10108 15204
rect 10164 15148 11788 15204
rect 11844 15148 11854 15204
rect 16146 15148 16156 15204
rect 16212 15148 18396 15204
rect 18452 15148 18462 15204
rect 6860 15092 6916 15148
rect 18844 15092 18900 15260
rect 19506 15148 19516 15204
rect 19572 15148 20748 15204
rect 20804 15148 20814 15204
rect 31724 15092 31780 15260
rect 32732 15092 32788 15372
rect 37772 15148 38556 15204
rect 38612 15148 39564 15204
rect 39620 15148 39630 15204
rect 6738 15036 6748 15092
rect 6804 15036 6916 15092
rect 18834 15036 18844 15092
rect 18900 15036 18910 15092
rect 31714 15036 31724 15092
rect 31780 15036 31790 15092
rect 32722 15036 32732 15092
rect 32788 15036 32798 15092
rect 33058 15036 33068 15092
rect 33124 15036 35308 15092
rect 35364 15036 35374 15092
rect 11890 14924 11900 14980
rect 11956 14924 17612 14980
rect 17668 14924 17678 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 13570 14812 13580 14868
rect 13636 14812 15260 14868
rect 15316 14812 15326 14868
rect 3490 14700 3500 14756
rect 3556 14700 4508 14756
rect 4564 14700 4574 14756
rect 17938 14700 17948 14756
rect 18004 14700 18620 14756
rect 18676 14700 18686 14756
rect 29586 14588 29596 14644
rect 29652 14588 30940 14644
rect 30996 14588 31006 14644
rect 37772 14532 37828 15148
rect 4946 14476 4956 14532
rect 5012 14476 7308 14532
rect 7364 14476 7374 14532
rect 19506 14476 19516 14532
rect 19572 14476 19684 14532
rect 23874 14476 23884 14532
rect 23940 14476 27132 14532
rect 27188 14476 27198 14532
rect 37772 14476 37884 14532
rect 37940 14476 37950 14532
rect 19628 14420 19684 14476
rect 19628 14364 23772 14420
rect 23828 14364 25228 14420
rect 25284 14364 25294 14420
rect 29698 14364 29708 14420
rect 29764 14364 30604 14420
rect 30660 14364 35532 14420
rect 35588 14364 35598 14420
rect 11666 14252 11676 14308
rect 11732 14252 13468 14308
rect 13524 14252 14588 14308
rect 14644 14252 14654 14308
rect 16258 14252 16268 14308
rect 16324 14252 22988 14308
rect 23044 14252 26012 14308
rect 26068 14252 26078 14308
rect 28690 14252 28700 14308
rect 28756 14252 30380 14308
rect 30436 14252 30446 14308
rect 31042 14252 31052 14308
rect 31108 14252 37100 14308
rect 37156 14252 37166 14308
rect 38322 14252 38332 14308
rect 38388 14252 39676 14308
rect 39732 14252 39742 14308
rect 17826 14140 17836 14196
rect 17892 14140 18284 14196
rect 18340 14140 18732 14196
rect 18788 14140 18798 14196
rect 19394 14140 19404 14196
rect 19460 14140 19684 14196
rect 38098 14140 38108 14196
rect 38164 14140 38556 14196
rect 38612 14140 38622 14196
rect 19628 14084 19684 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 19618 14028 19628 14084
rect 19684 14028 19694 14084
rect 8194 13916 8204 13972
rect 8260 13916 9660 13972
rect 9716 13916 12348 13972
rect 12404 13916 12414 13972
rect 15138 13916 15148 13972
rect 15204 13916 17612 13972
rect 17668 13916 18396 13972
rect 18452 13916 18462 13972
rect 19954 13916 19964 13972
rect 20020 13916 20300 13972
rect 20356 13916 20366 13972
rect 36418 13916 36428 13972
rect 36484 13916 37660 13972
rect 37716 13916 38444 13972
rect 38500 13916 38510 13972
rect 33254 13804 33292 13860
rect 33348 13804 33358 13860
rect 34402 13804 34412 13860
rect 34468 13804 35868 13860
rect 35924 13804 35934 13860
rect 37426 13804 37436 13860
rect 37492 13804 38556 13860
rect 38612 13804 38622 13860
rect 12002 13692 12012 13748
rect 12068 13692 16268 13748
rect 16324 13692 16334 13748
rect 17938 13692 17948 13748
rect 18004 13692 19180 13748
rect 19236 13692 24780 13748
rect 24836 13692 24846 13748
rect 37314 13692 37324 13748
rect 37380 13692 38892 13748
rect 38948 13692 38958 13748
rect 1922 13580 1932 13636
rect 1988 13580 2268 13636
rect 2324 13580 2334 13636
rect 5170 13580 5180 13636
rect 5236 13580 5628 13636
rect 5684 13580 15036 13636
rect 15092 13580 15596 13636
rect 15652 13580 15662 13636
rect 18582 13580 18620 13636
rect 18676 13580 18686 13636
rect 20178 13580 20188 13636
rect 20244 13580 21420 13636
rect 21476 13580 22652 13636
rect 22708 13580 22718 13636
rect 22866 13580 22876 13636
rect 22932 13580 27916 13636
rect 27972 13580 27982 13636
rect 7186 13468 7196 13524
rect 7252 13468 8092 13524
rect 8148 13468 8158 13524
rect 9538 13468 9548 13524
rect 9604 13468 10668 13524
rect 10724 13468 11452 13524
rect 11508 13468 11518 13524
rect 22754 13468 22764 13524
rect 22820 13468 23884 13524
rect 23940 13468 23950 13524
rect 33170 13468 33180 13524
rect 33236 13468 33684 13524
rect 36754 13468 36764 13524
rect 36820 13468 36932 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 33628 13300 33684 13468
rect 36876 13412 36932 13468
rect 37324 13468 38108 13524
rect 38164 13468 39340 13524
rect 39396 13468 39406 13524
rect 37324 13412 37380 13468
rect 36876 13356 37380 13412
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 33618 13244 33628 13300
rect 33684 13244 33694 13300
rect 17938 12908 17948 12964
rect 18004 12908 19068 12964
rect 19124 12908 19134 12964
rect 21970 12908 21980 12964
rect 22036 12908 22316 12964
rect 22372 12908 22764 12964
rect 22820 12908 22830 12964
rect 25554 12908 25564 12964
rect 25620 12908 26236 12964
rect 26292 12908 28140 12964
rect 28196 12908 28206 12964
rect 28466 12908 28476 12964
rect 28532 12908 29932 12964
rect 29988 12908 30940 12964
rect 30996 12908 31006 12964
rect 32610 12908 32620 12964
rect 32676 12908 33404 12964
rect 33460 12908 33470 12964
rect 34178 12908 34188 12964
rect 34244 12908 34972 12964
rect 35028 12908 35038 12964
rect 35634 12908 35644 12964
rect 35700 12908 36988 12964
rect 37044 12908 37054 12964
rect 11106 12796 11116 12852
rect 11172 12796 13580 12852
rect 13636 12796 13646 12852
rect 19506 12796 19516 12852
rect 19572 12796 22988 12852
rect 23044 12796 25340 12852
rect 25396 12796 26012 12852
rect 26068 12796 26078 12852
rect 19404 12684 19740 12740
rect 19796 12684 23436 12740
rect 23492 12684 23502 12740
rect 26786 12684 26796 12740
rect 26852 12684 26908 12908
rect 29372 12852 29428 12908
rect 29362 12796 29372 12852
rect 29428 12796 29438 12852
rect 30034 12796 30044 12852
rect 30100 12796 30716 12852
rect 30772 12796 30782 12852
rect 34290 12796 34300 12852
rect 34356 12796 34748 12852
rect 34804 12796 34814 12852
rect 37762 12796 37772 12852
rect 37828 12796 38444 12852
rect 38500 12796 38510 12852
rect 32386 12684 32396 12740
rect 32452 12684 33068 12740
rect 33124 12684 33134 12740
rect 33394 12684 33404 12740
rect 33460 12684 35196 12740
rect 35252 12684 35262 12740
rect 19404 12516 19460 12684
rect 27794 12572 27804 12628
rect 27860 12572 30828 12628
rect 30884 12572 30894 12628
rect 31602 12572 31612 12628
rect 31668 12572 34524 12628
rect 34580 12572 34860 12628
rect 34916 12572 35868 12628
rect 35924 12572 35934 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 18946 12460 18956 12516
rect 19012 12460 19460 12516
rect 23090 12460 23100 12516
rect 23156 12460 26236 12516
rect 26292 12460 27132 12516
rect 27188 12460 27198 12516
rect 15810 12348 15820 12404
rect 15876 12348 18284 12404
rect 18340 12348 18350 12404
rect 18834 12348 18844 12404
rect 18900 12348 19404 12404
rect 19460 12348 21420 12404
rect 21476 12348 21486 12404
rect 26002 12348 26012 12404
rect 26068 12348 27692 12404
rect 27748 12348 27758 12404
rect 30258 12348 30268 12404
rect 30324 12348 31500 12404
rect 31556 12348 31566 12404
rect 31714 12348 31724 12404
rect 31780 12348 33964 12404
rect 34020 12348 34030 12404
rect 26852 12236 29148 12292
rect 29204 12236 29214 12292
rect 34066 12236 34076 12292
rect 34132 12236 37212 12292
rect 37268 12236 37660 12292
rect 37716 12236 37726 12292
rect 8194 12124 8204 12180
rect 8260 12124 8876 12180
rect 8932 12124 8942 12180
rect 13794 12124 13804 12180
rect 13860 12124 22204 12180
rect 22260 12124 22764 12180
rect 22820 12124 22830 12180
rect 26852 12068 26908 12236
rect 27458 12124 27468 12180
rect 27524 12124 28588 12180
rect 28644 12124 28654 12180
rect 24770 12012 24780 12068
rect 24836 12012 26908 12068
rect 37314 12012 37324 12068
rect 37380 12012 38332 12068
rect 38388 12012 38398 12068
rect 19058 11900 19068 11956
rect 19124 11900 19516 11956
rect 19572 11900 19582 11956
rect 22194 11900 22204 11956
rect 22260 11900 24444 11956
rect 24500 11900 24510 11956
rect 26786 11900 26796 11956
rect 26852 11900 26908 11956
rect 26964 11900 26974 11956
rect 17714 11788 17724 11844
rect 17780 11788 18620 11844
rect 18676 11788 18686 11844
rect 25442 11788 25452 11844
rect 25508 11788 27468 11844
rect 27524 11788 27534 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 5954 11564 5964 11620
rect 6020 11564 6748 11620
rect 6804 11564 11452 11620
rect 11508 11564 12236 11620
rect 12292 11564 12302 11620
rect 17826 11564 17836 11620
rect 17892 11564 18844 11620
rect 18900 11564 18910 11620
rect 35522 11564 35532 11620
rect 35588 11564 37996 11620
rect 38052 11564 38062 11620
rect 12450 11452 12460 11508
rect 12516 11452 13692 11508
rect 13748 11452 14700 11508
rect 14756 11452 14766 11508
rect 18610 11452 18620 11508
rect 18676 11452 18732 11508
rect 18788 11452 19404 11508
rect 19460 11452 19470 11508
rect 23202 11452 23212 11508
rect 23268 11452 27244 11508
rect 27300 11452 30156 11508
rect 30212 11452 30222 11508
rect 38098 11452 38108 11508
rect 38164 11452 38556 11508
rect 38612 11452 38622 11508
rect 17602 11340 17612 11396
rect 17668 11340 18060 11396
rect 18116 11340 19068 11396
rect 19124 11340 19964 11396
rect 20020 11340 20030 11396
rect 20738 11340 20748 11396
rect 20804 11340 21868 11396
rect 21924 11340 21934 11396
rect 22082 11340 22092 11396
rect 22148 11340 22988 11396
rect 23044 11340 23054 11396
rect 23426 11340 23436 11396
rect 23492 11340 25788 11396
rect 25844 11340 26460 11396
rect 26516 11340 26526 11396
rect 22988 11284 23044 11340
rect 9986 11228 9996 11284
rect 10052 11228 11564 11284
rect 11620 11228 15148 11284
rect 17938 11228 17948 11284
rect 18004 11228 21644 11284
rect 21700 11228 21710 11284
rect 22988 11228 23660 11284
rect 23716 11228 23726 11284
rect 24098 11228 24108 11284
rect 24164 11228 26572 11284
rect 26628 11228 26638 11284
rect 15092 11172 15148 11228
rect 23660 11172 23716 11228
rect 6178 11116 6188 11172
rect 6244 11116 7084 11172
rect 7140 11116 7150 11172
rect 8082 11116 8092 11172
rect 8148 11116 12348 11172
rect 12404 11116 12414 11172
rect 15026 11116 15036 11172
rect 15092 11116 21756 11172
rect 21812 11116 22092 11172
rect 22148 11116 22158 11172
rect 23660 11116 26348 11172
rect 26404 11116 29708 11172
rect 29764 11116 29774 11172
rect 32050 11116 32060 11172
rect 32116 11116 33180 11172
rect 33236 11116 33246 11172
rect 35410 11116 35420 11172
rect 35476 11116 37436 11172
rect 37492 11116 37502 11172
rect 37650 11116 37660 11172
rect 37716 11116 37754 11172
rect 18162 11004 18172 11060
rect 18228 11004 19516 11060
rect 19572 11004 19582 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 36530 10892 36540 10948
rect 36596 10892 37884 10948
rect 37940 10892 38108 10948
rect 38164 10892 38174 10948
rect 6514 10780 6524 10836
rect 6580 10780 7308 10836
rect 7364 10780 7374 10836
rect 19394 10780 19404 10836
rect 19460 10780 19740 10836
rect 19796 10780 20188 10836
rect 20244 10780 20254 10836
rect 36194 10780 36204 10836
rect 36260 10780 37436 10836
rect 37492 10780 38444 10836
rect 38500 10780 38510 10836
rect 33506 10668 33516 10724
rect 33572 10668 37324 10724
rect 37380 10668 38780 10724
rect 38836 10668 38846 10724
rect 19618 10556 19628 10612
rect 19684 10556 21196 10612
rect 21252 10556 22876 10612
rect 22932 10556 24556 10612
rect 24612 10556 24622 10612
rect 27010 10556 27020 10612
rect 27076 10556 27916 10612
rect 27972 10556 29036 10612
rect 29092 10556 29820 10612
rect 29876 10556 29886 10612
rect 32498 10556 32508 10612
rect 32564 10556 33740 10612
rect 33796 10556 33806 10612
rect 35298 10556 35308 10612
rect 35364 10556 35756 10612
rect 35812 10556 35822 10612
rect 7410 10444 7420 10500
rect 7476 10444 8316 10500
rect 8372 10444 8382 10500
rect 23090 10444 23100 10500
rect 23156 10444 23996 10500
rect 24052 10444 24062 10500
rect 33954 10444 33964 10500
rect 34020 10444 35084 10500
rect 35140 10444 35980 10500
rect 36036 10444 36046 10500
rect 29922 10332 29932 10388
rect 29988 10332 33516 10388
rect 33572 10332 33582 10388
rect 32498 10220 32508 10276
rect 32564 10220 33628 10276
rect 33684 10220 33694 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 13234 10108 13244 10164
rect 13300 10108 13310 10164
rect 24882 10108 24892 10164
rect 24948 10108 26012 10164
rect 26068 10108 26078 10164
rect 28354 10108 28364 10164
rect 28420 10108 29596 10164
rect 29652 10108 29662 10164
rect 31826 10108 31836 10164
rect 31892 10108 32004 10164
rect 36418 10108 36428 10164
rect 36484 10108 38108 10164
rect 38164 10108 39116 10164
rect 39172 10108 39182 10164
rect 13244 10052 13300 10108
rect 7522 9996 7532 10052
rect 7588 9996 8652 10052
rect 8708 9996 8718 10052
rect 13244 9996 16940 10052
rect 16996 9996 17006 10052
rect 29138 9996 29148 10052
rect 29204 9996 30492 10052
rect 30548 9996 30558 10052
rect 26674 9884 26684 9940
rect 26740 9884 27580 9940
rect 27636 9884 27646 9940
rect 31948 9828 32004 10108
rect 32162 9884 32172 9940
rect 32228 9884 33292 9940
rect 33348 9884 33358 9940
rect 36530 9884 36540 9940
rect 36596 9884 37212 9940
rect 37268 9884 37278 9940
rect 27346 9772 27356 9828
rect 27412 9772 28252 9828
rect 28308 9772 28318 9828
rect 29138 9772 29148 9828
rect 29204 9772 31276 9828
rect 31332 9772 31342 9828
rect 31948 9772 32508 9828
rect 32564 9772 34860 9828
rect 34916 9772 36316 9828
rect 36372 9772 36382 9828
rect 36642 9772 36652 9828
rect 36708 9772 37548 9828
rect 37604 9772 37614 9828
rect 38210 9772 38220 9828
rect 38276 9772 39228 9828
rect 39284 9772 39294 9828
rect 3154 9660 3164 9716
rect 3220 9660 4060 9716
rect 4116 9660 4126 9716
rect 13794 9660 13804 9716
rect 13860 9660 18396 9716
rect 18452 9660 20076 9716
rect 20132 9660 22540 9716
rect 22596 9660 23548 9716
rect 23604 9660 23614 9716
rect 28130 9660 28140 9716
rect 28196 9660 28588 9716
rect 28644 9660 32284 9716
rect 32340 9660 32620 9716
rect 32676 9660 33068 9716
rect 33124 9660 33134 9716
rect 37212 9660 37996 9716
rect 38052 9660 38062 9716
rect 37212 9604 37268 9660
rect 9986 9548 9996 9604
rect 10052 9548 13244 9604
rect 13300 9548 13310 9604
rect 31266 9548 31276 9604
rect 31332 9548 32172 9604
rect 32228 9548 32238 9604
rect 32834 9548 32844 9604
rect 32900 9548 33292 9604
rect 33348 9548 35644 9604
rect 35700 9548 35710 9604
rect 37202 9548 37212 9604
rect 37268 9548 37278 9604
rect 37426 9548 37436 9604
rect 37492 9548 38892 9604
rect 38948 9548 38958 9604
rect 9202 9436 9212 9492
rect 9268 9436 15372 9492
rect 15428 9436 17388 9492
rect 17444 9436 17454 9492
rect 28242 9436 28252 9492
rect 28308 9436 31724 9492
rect 31780 9436 34300 9492
rect 34356 9436 34366 9492
rect 36306 9436 36316 9492
rect 36372 9436 39004 9492
rect 39060 9436 39070 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 29810 9324 29820 9380
rect 29876 9324 31052 9380
rect 31108 9324 32732 9380
rect 32788 9324 37100 9380
rect 37156 9324 37166 9380
rect 37762 9324 37772 9380
rect 37828 9324 38108 9380
rect 38164 9324 38174 9380
rect 8642 9212 8652 9268
rect 8708 9212 9660 9268
rect 9716 9212 9726 9268
rect 30818 9212 30828 9268
rect 30884 9212 38388 9268
rect 38332 9156 38388 9212
rect 31826 9100 31836 9156
rect 31892 9100 34076 9156
rect 34132 9100 34142 9156
rect 36530 9100 36540 9156
rect 36596 9100 36988 9156
rect 37044 9100 37054 9156
rect 37286 9100 37324 9156
rect 37380 9100 37390 9156
rect 38322 9100 38332 9156
rect 38388 9100 38398 9156
rect 5954 8988 5964 9044
rect 6020 8988 6300 9044
rect 6356 8988 9436 9044
rect 9492 8988 9502 9044
rect 16930 8988 16940 9044
rect 16996 8988 24668 9044
rect 24724 8988 25340 9044
rect 25396 8988 26124 9044
rect 26180 8988 26190 9044
rect 34626 8988 34636 9044
rect 34692 8988 35532 9044
rect 35588 8988 36204 9044
rect 36260 8988 36270 9044
rect 11778 8876 11788 8932
rect 11844 8876 14140 8932
rect 14196 8876 14206 8932
rect 4610 8764 4620 8820
rect 4676 8764 6972 8820
rect 7028 8764 8876 8820
rect 8932 8764 8942 8820
rect 29474 8764 29484 8820
rect 29540 8764 30156 8820
rect 30212 8764 30222 8820
rect 35970 8764 35980 8820
rect 36036 8764 36876 8820
rect 36932 8764 36942 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 11330 8540 11340 8596
rect 11396 8540 12460 8596
rect 12516 8540 12526 8596
rect 31042 8540 31052 8596
rect 31108 8540 32004 8596
rect 5506 8428 5516 8484
rect 5572 8428 12124 8484
rect 12180 8428 12190 8484
rect 31948 8372 32004 8540
rect 36418 8428 36428 8484
rect 36484 8428 38332 8484
rect 38388 8428 38398 8484
rect 8418 8316 8428 8372
rect 8484 8316 9324 8372
rect 9380 8316 9390 8372
rect 12674 8316 12684 8372
rect 12740 8316 15932 8372
rect 15988 8316 16492 8372
rect 16548 8316 18732 8372
rect 18788 8316 18798 8372
rect 27234 8316 27244 8372
rect 27300 8316 30492 8372
rect 30548 8316 30558 8372
rect 31948 8316 32620 8372
rect 32676 8316 32686 8372
rect 35858 8316 35868 8372
rect 35924 8316 37772 8372
rect 37828 8316 37838 8372
rect 37986 8316 37996 8372
rect 38052 8316 39228 8372
rect 39284 8316 39294 8372
rect 31948 8260 32004 8316
rect 11666 8204 11676 8260
rect 11732 8204 13692 8260
rect 13748 8204 13758 8260
rect 13906 8204 13916 8260
rect 13972 8204 15260 8260
rect 15316 8204 15326 8260
rect 16034 8204 16044 8260
rect 16100 8204 20748 8260
rect 20804 8204 20814 8260
rect 29922 8204 29932 8260
rect 29988 8204 32004 8260
rect 33394 8204 33404 8260
rect 33460 8204 34524 8260
rect 34580 8204 35756 8260
rect 35812 8204 35822 8260
rect 35980 8204 36316 8260
rect 36372 8204 36652 8260
rect 36708 8204 36718 8260
rect 37314 8204 37324 8260
rect 37380 8204 38556 8260
rect 38612 8204 38622 8260
rect 35980 8148 36036 8204
rect 5058 8092 5068 8148
rect 5124 8092 5628 8148
rect 5684 8092 5694 8148
rect 9874 8092 9884 8148
rect 9940 8092 10556 8148
rect 10612 8092 12236 8148
rect 12292 8092 12302 8148
rect 14690 8092 14700 8148
rect 14756 8092 15372 8148
rect 15428 8092 15438 8148
rect 25554 8092 25564 8148
rect 25620 8092 29260 8148
rect 29316 8092 29326 8148
rect 32722 8092 32732 8148
rect 32788 8092 34972 8148
rect 35028 8092 36036 8148
rect 36316 8092 36988 8148
rect 37044 8092 38108 8148
rect 38164 8092 38174 8148
rect 8866 7980 8876 8036
rect 8932 7980 13580 8036
rect 13636 7980 13646 8036
rect 26852 7980 30828 8036
rect 30884 7980 30894 8036
rect 31042 7980 31052 8036
rect 31108 7980 31146 8036
rect 26852 7924 26908 7980
rect 36316 7924 36372 8092
rect 36642 7980 36652 8036
rect 36708 7980 39228 8036
rect 39284 7980 39294 8036
rect 11218 7868 11228 7924
rect 11284 7868 16156 7924
rect 16212 7868 16222 7924
rect 24434 7868 24444 7924
rect 24500 7868 26908 7924
rect 36306 7868 36316 7924
rect 36372 7868 36382 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 26562 7756 26572 7812
rect 26628 7756 30940 7812
rect 30996 7756 31724 7812
rect 31780 7756 33180 7812
rect 33236 7756 33516 7812
rect 33572 7756 33582 7812
rect 3714 7644 3724 7700
rect 3780 7644 4956 7700
rect 5012 7644 9660 7700
rect 9716 7644 9726 7700
rect 17042 7644 17052 7700
rect 17108 7644 17724 7700
rect 17780 7644 22652 7700
rect 22708 7644 22718 7700
rect 26338 7644 26348 7700
rect 26404 7644 28588 7700
rect 28644 7644 28654 7700
rect 29586 7644 29596 7700
rect 29652 7644 31108 7700
rect 31266 7644 31276 7700
rect 31332 7644 32172 7700
rect 32228 7644 32238 7700
rect 31052 7588 31108 7644
rect 8082 7532 8092 7588
rect 8148 7532 8652 7588
rect 8708 7532 8718 7588
rect 9762 7532 9772 7588
rect 9828 7532 10668 7588
rect 10724 7532 10734 7588
rect 17938 7532 17948 7588
rect 18004 7532 25676 7588
rect 25732 7532 26124 7588
rect 26180 7532 26190 7588
rect 28466 7532 28476 7588
rect 28532 7532 30156 7588
rect 30212 7532 30222 7588
rect 31052 7532 33852 7588
rect 33908 7532 35644 7588
rect 35700 7532 35710 7588
rect 35970 7532 35980 7588
rect 36036 7532 37212 7588
rect 37268 7532 37996 7588
rect 38052 7532 38062 7588
rect 10210 7420 10220 7476
rect 10276 7420 13692 7476
rect 13748 7420 13758 7476
rect 20962 7420 20972 7476
rect 21028 7420 22092 7476
rect 22148 7420 22158 7476
rect 27906 7420 27916 7476
rect 27972 7420 28812 7476
rect 28868 7420 29372 7476
rect 29428 7420 29438 7476
rect 29810 7420 29820 7476
rect 29876 7420 30604 7476
rect 30660 7420 32508 7476
rect 32564 7420 33628 7476
rect 33684 7420 33694 7476
rect 28578 7308 28588 7364
rect 28644 7308 29596 7364
rect 29652 7308 29662 7364
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 7186 6860 7196 6916
rect 7252 6860 8428 6916
rect 8484 6860 8494 6916
rect 8642 6860 8652 6916
rect 8708 6860 11004 6916
rect 11060 6860 11676 6916
rect 11732 6860 11742 6916
rect 13682 6860 13692 6916
rect 13748 6860 15820 6916
rect 15876 6860 16716 6916
rect 16772 6860 16782 6916
rect 29698 6860 29708 6916
rect 29764 6860 31948 6916
rect 32004 6860 32014 6916
rect 34402 6860 34412 6916
rect 34468 6860 39004 6916
rect 39060 6860 39070 6916
rect 5394 6748 5404 6804
rect 5460 6748 6860 6804
rect 6916 6748 7980 6804
rect 8036 6748 8046 6804
rect 10658 6748 10668 6804
rect 10724 6748 11452 6804
rect 11508 6748 11518 6804
rect 12898 6748 12908 6804
rect 12964 6748 15484 6804
rect 15540 6748 15550 6804
rect 36194 6748 36204 6804
rect 36260 6748 36876 6804
rect 36932 6748 36942 6804
rect 6290 6636 6300 6692
rect 6356 6636 8092 6692
rect 8148 6636 8158 6692
rect 13458 6636 13468 6692
rect 13524 6636 14364 6692
rect 14420 6636 14430 6692
rect 15334 6636 15372 6692
rect 15428 6636 15438 6692
rect 15586 6636 15596 6692
rect 15652 6636 21084 6692
rect 21140 6636 21150 6692
rect 22866 6636 22876 6692
rect 22932 6636 23884 6692
rect 23940 6636 23950 6692
rect 27570 6636 27580 6692
rect 27636 6636 29372 6692
rect 29428 6636 29438 6692
rect 34850 6636 34860 6692
rect 34916 6636 35868 6692
rect 35924 6636 35934 6692
rect 38612 6636 38892 6692
rect 38948 6636 38958 6692
rect 15596 6580 15652 6636
rect 5618 6524 5628 6580
rect 5684 6524 6748 6580
rect 6804 6524 6814 6580
rect 7746 6524 7756 6580
rect 7812 6524 8764 6580
rect 8820 6524 8830 6580
rect 14130 6524 14140 6580
rect 14196 6524 15652 6580
rect 16146 6524 16156 6580
rect 16212 6524 16940 6580
rect 16996 6524 19628 6580
rect 19684 6524 19694 6580
rect 21746 6524 21756 6580
rect 21812 6524 24220 6580
rect 24276 6524 24286 6580
rect 31602 6524 31612 6580
rect 31668 6524 34300 6580
rect 34356 6524 37548 6580
rect 37604 6524 37614 6580
rect 38612 6468 38668 6636
rect 1922 6412 1932 6468
rect 1988 6412 4956 6468
rect 5012 6412 5292 6468
rect 5348 6412 8876 6468
rect 8932 6412 9548 6468
rect 9604 6412 12684 6468
rect 12740 6412 16380 6468
rect 16436 6412 17836 6468
rect 17892 6412 17902 6468
rect 28130 6412 28140 6468
rect 28196 6412 28812 6468
rect 28868 6412 29596 6468
rect 29652 6412 29662 6468
rect 33842 6412 33852 6468
rect 33908 6412 36764 6468
rect 36820 6412 38668 6468
rect 14130 6300 14140 6356
rect 14196 6300 15372 6356
rect 15428 6300 15438 6356
rect 22866 6300 22876 6356
rect 22932 6300 28364 6356
rect 28420 6300 28430 6356
rect 35970 6300 35980 6356
rect 36036 6300 39116 6356
rect 39172 6300 39182 6356
rect 15372 6244 15428 6300
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 15362 6188 15372 6244
rect 15428 6188 15438 6244
rect 32274 6188 32284 6244
rect 32340 6188 35532 6244
rect 35588 6188 36652 6244
rect 36708 6188 36718 6244
rect 36876 6188 37884 6244
rect 37940 6188 37950 6244
rect 36876 6132 36932 6188
rect 10882 6076 10892 6132
rect 10948 6076 12012 6132
rect 12068 6076 12078 6132
rect 13122 6076 13132 6132
rect 13188 6076 13916 6132
rect 13972 6076 36932 6132
rect 37314 6076 37324 6132
rect 37380 6076 39340 6132
rect 39396 6076 39406 6132
rect 5730 5964 5740 6020
rect 5796 5964 7644 6020
rect 7700 5964 9660 6020
rect 9716 5964 9726 6020
rect 11778 5964 11788 6020
rect 11844 5964 12460 6020
rect 12516 5964 15036 6020
rect 15092 5964 15102 6020
rect 24658 5964 24668 6020
rect 24724 5964 25340 6020
rect 25396 5964 25406 6020
rect 4946 5852 4956 5908
rect 5012 5852 6076 5908
rect 6132 5852 6142 5908
rect 10322 5852 10332 5908
rect 10388 5852 17388 5908
rect 17444 5852 17454 5908
rect 19618 5852 19628 5908
rect 19684 5852 21868 5908
rect 21924 5852 21934 5908
rect 32050 5852 32060 5908
rect 32116 5852 36540 5908
rect 36596 5852 36606 5908
rect 5842 5740 5852 5796
rect 5908 5740 7308 5796
rect 7364 5740 7374 5796
rect 10546 5740 10556 5796
rect 10612 5740 12908 5796
rect 12964 5740 12974 5796
rect 16258 5740 16268 5796
rect 16324 5740 17612 5796
rect 17668 5740 17678 5796
rect 32722 5740 32732 5796
rect 32788 5740 33628 5796
rect 33684 5740 35980 5796
rect 36036 5740 36046 5796
rect 6066 5628 6076 5684
rect 6132 5628 7084 5684
rect 7140 5628 7150 5684
rect 33842 5628 33852 5684
rect 33908 5628 35868 5684
rect 35924 5628 35934 5684
rect 5618 5516 5628 5572
rect 5684 5516 8092 5572
rect 8148 5516 8158 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 28578 5404 28588 5460
rect 28644 5404 29260 5460
rect 29316 5404 29326 5460
rect 8642 5292 8652 5348
rect 8708 5292 12796 5348
rect 12852 5292 12862 5348
rect 15092 5292 21308 5348
rect 21364 5292 21756 5348
rect 21812 5292 22092 5348
rect 22148 5292 22158 5348
rect 26852 5292 28812 5348
rect 28868 5292 28878 5348
rect 35634 5292 35644 5348
rect 35700 5292 39004 5348
rect 39060 5292 39070 5348
rect 15092 5236 15148 5292
rect 4722 5180 4732 5236
rect 4788 5180 5516 5236
rect 5572 5180 5582 5236
rect 7746 5180 7756 5236
rect 7812 5180 8988 5236
rect 9044 5180 9054 5236
rect 9202 5180 9212 5236
rect 9268 5180 9660 5236
rect 9716 5180 15148 5236
rect 16258 5180 16268 5236
rect 16324 5180 17948 5236
rect 18004 5180 18014 5236
rect 26786 5180 26796 5236
rect 26852 5180 26908 5292
rect 27234 5180 27244 5236
rect 27300 5180 28588 5236
rect 28644 5180 32060 5236
rect 32116 5180 32126 5236
rect 37650 5180 37660 5236
rect 37716 5180 39228 5236
rect 39284 5180 39294 5236
rect 27244 5124 27300 5180
rect 8530 5068 8540 5124
rect 8596 5068 9548 5124
rect 9604 5068 9614 5124
rect 16930 5068 16940 5124
rect 16996 5068 17612 5124
rect 17668 5068 17678 5124
rect 23874 5068 23884 5124
rect 23940 5068 25452 5124
rect 25508 5068 26124 5124
rect 26180 5068 27300 5124
rect 31266 5068 31276 5124
rect 31332 5068 34524 5124
rect 34580 5068 34590 5124
rect 35298 5068 35308 5124
rect 35364 5068 36204 5124
rect 36260 5068 36270 5124
rect 2594 4956 2604 5012
rect 2660 4956 5964 5012
rect 6020 4956 6030 5012
rect 34066 4956 34076 5012
rect 34132 4956 37100 5012
rect 37156 4956 37772 5012
rect 37828 4956 37838 5012
rect 38612 4956 38780 5012
rect 38836 4956 38846 5012
rect 38612 4900 38668 4956
rect 35970 4844 35980 4900
rect 36036 4844 36764 4900
rect 36820 4844 36830 4900
rect 37426 4844 37436 4900
rect 37492 4844 38668 4900
rect 34514 4732 34524 4788
rect 34580 4732 39116 4788
rect 39172 4732 39182 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 32610 4620 32620 4676
rect 32676 4620 38108 4676
rect 38164 4620 38174 4676
rect 3938 4508 3948 4564
rect 4004 4508 10556 4564
rect 10612 4508 10622 4564
rect 16594 4396 16604 4452
rect 16660 4396 17388 4452
rect 17444 4396 17454 4452
rect 31938 4396 31948 4452
rect 32004 4396 33516 4452
rect 33572 4396 36764 4452
rect 36820 4396 36830 4452
rect 4722 4284 4732 4340
rect 4788 4284 5516 4340
rect 5572 4284 5582 4340
rect 13794 4284 13804 4340
rect 13860 4284 14924 4340
rect 14980 4284 14990 4340
rect 28354 4284 28364 4340
rect 28420 4284 29036 4340
rect 29092 4284 29102 4340
rect 37426 4172 37436 4228
rect 37492 4172 38892 4228
rect 38948 4172 38958 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 7746 3612 7756 3668
rect 7812 3612 8540 3668
rect 8596 3612 8606 3668
rect 12114 3612 12124 3668
rect 12180 3612 13132 3668
rect 13188 3612 13198 3668
rect 5058 3500 5068 3556
rect 5124 3500 5740 3556
rect 5796 3500 5806 3556
rect 14354 3500 14364 3556
rect 14420 3500 16940 3556
rect 16996 3500 17006 3556
rect 31490 3500 31500 3556
rect 31556 3500 33404 3556
rect 33460 3500 38668 3556
rect 38612 3444 38668 3500
rect 13906 3388 13916 3444
rect 13972 3388 14812 3444
rect 14868 3388 14878 3444
rect 15250 3388 15260 3444
rect 15316 3388 18508 3444
rect 18564 3388 18574 3444
rect 31042 3388 31052 3444
rect 31108 3388 35420 3444
rect 35476 3388 37996 3444
rect 38052 3388 38062 3444
rect 38612 3388 39452 3444
rect 39508 3388 39518 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 17276 33180 17332 33236
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 17276 32172 17332 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 8204 22652 8260 22708
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 8204 19068 8260 19124
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 33292 13804 33348 13860
rect 18620 13580 18676 13636
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 37660 12236 37716 12292
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 18620 11452 18676 11508
rect 37660 11116 37716 11172
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 37324 10668 37380 10724
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 33292 9548 33348 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 31052 9324 31108 9380
rect 37324 9100 37380 9156
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 31052 7980 31108 8036
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 15372 6636 15428 6692
rect 15372 6300 15428 6356
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 41612
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 19808 40796 20128 41612
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 17276 33236 17332 33246
rect 17276 32228 17332 33180
rect 17276 32162 17332 32172
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 8204 22708 8260 22718
rect 8204 19124 8260 22652
rect 8204 19058 8260 19068
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 18620 13636 18676 13646
rect 18620 11508 18676 13580
rect 18620 11442 18676 11452
rect 19808 12572 20128 14084
rect 35168 41580 35488 41612
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 33292 13860 33348 13870
rect 33292 9604 33348 13804
rect 33292 9538 33348 9548
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 37660 12292 37716 12302
rect 37660 11172 37716 12236
rect 37660 11106 37716 11116
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 31052 9380 31108 9390
rect 31052 8036 31108 9324
rect 31052 7970 31108 7980
rect 35168 8652 35488 10164
rect 37324 10724 37380 10734
rect 37324 9156 37380 10668
rect 37324 9090 37380 9100
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 15372 6692 15428 6702
rect 15372 6356 15428 6636
rect 15372 6290 15428 6300
rect 19808 6300 20128 7812
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0553_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0554_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12768 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0555_
timestamp 1698431365
transform -1 0 14896 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0556_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14672 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0557_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16240 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0558_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25760 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0559_
timestamp 1698431365
transform -1 0 21840 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0560_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0561_
timestamp 1698431365
transform 1 0 26208 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0562_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26544 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0563_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20048 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0564_
timestamp 1698431365
transform 1 0 8176 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0565_
timestamp 1698431365
transform -1 0 7392 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0566_
timestamp 1698431365
transform 1 0 6160 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0567_
timestamp 1698431365
transform -1 0 7056 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0568_
timestamp 1698431365
transform 1 0 5488 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0569_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0570_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0571_
timestamp 1698431365
transform -1 0 7840 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0572_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8400 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0573_
timestamp 1698431365
transform 1 0 31136 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0574_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0575_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26544 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0576_
timestamp 1698431365
transform -1 0 27440 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0577_
timestamp 1698431365
transform -1 0 15344 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0578_
timestamp 1698431365
transform 1 0 14784 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0579_
timestamp 1698431365
transform -1 0 13776 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0580_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14448 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0581_
timestamp 1698431365
transform 1 0 14560 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0582_
timestamp 1698431365
transform -1 0 21952 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0583_
timestamp 1698431365
transform 1 0 15680 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0584_
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0585_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0586_
timestamp 1698431365
transform 1 0 23632 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0587_
timestamp 1698431365
transform -1 0 24528 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0588_
timestamp 1698431365
transform 1 0 22400 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0589_
timestamp 1698431365
transform -1 0 19600 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0590_
timestamp 1698431365
transform 1 0 22512 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0591_
timestamp 1698431365
transform -1 0 24080 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0592_
timestamp 1698431365
transform 1 0 18592 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0593_
timestamp 1698431365
transform 1 0 19488 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0594_
timestamp 1698431365
transform -1 0 20496 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0595_
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0596_
timestamp 1698431365
transform -1 0 6384 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0597_
timestamp 1698431365
transform 1 0 6160 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0598_
timestamp 1698431365
transform -1 0 7056 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0599_
timestamp 1698431365
transform -1 0 5264 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0600_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0601_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6496 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0602_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0603_
timestamp 1698431365
transform 1 0 7056 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0604_
timestamp 1698431365
transform -1 0 5600 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0605_
timestamp 1698431365
transform -1 0 10640 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0606_
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0607_
timestamp 1698431365
transform 1 0 7504 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0608_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9632 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0609_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0610_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0611_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14112 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0612_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0613_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13104 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0614_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0615_
timestamp 1698431365
transform -1 0 19712 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0616_
timestamp 1698431365
transform -1 0 11424 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0617_
timestamp 1698431365
transform 1 0 8400 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0618_
timestamp 1698431365
transform -1 0 5264 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0619_
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _0620_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8176 0 -1 21952
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0621_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7840 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0622_
timestamp 1698431365
transform 1 0 7952 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0623_
timestamp 1698431365
transform -1 0 11984 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0624_
timestamp 1698431365
transform -1 0 10864 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0625_
timestamp 1698431365
transform 1 0 20832 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0626_
timestamp 1698431365
transform -1 0 15792 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0627_
timestamp 1698431365
transform 1 0 12208 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0628_
timestamp 1698431365
transform -1 0 6944 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0629_
timestamp 1698431365
transform 1 0 12096 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0630_
timestamp 1698431365
transform 1 0 11312 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0631_
timestamp 1698431365
transform -1 0 12768 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0632_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10416 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0633_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0634_
timestamp 1698431365
transform 1 0 12208 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0635_
timestamp 1698431365
transform 1 0 11312 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0636_
timestamp 1698431365
transform 1 0 7056 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0637_
timestamp 1698431365
transform 1 0 7728 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0638_
timestamp 1698431365
transform 1 0 6272 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0639_
timestamp 1698431365
transform -1 0 5264 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0640_
timestamp 1698431365
transform 1 0 8736 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0641_
timestamp 1698431365
transform -1 0 15680 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0642_
timestamp 1698431365
transform -1 0 10416 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0643_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0644_
timestamp 1698431365
transform 1 0 5712 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0645_
timestamp 1698431365
transform -1 0 7728 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0646_
timestamp 1698431365
transform -1 0 7616 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0647_
timestamp 1698431365
transform -1 0 8512 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0648_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7840 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0649_
timestamp 1698431365
transform -1 0 12544 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0650_
timestamp 1698431365
transform 1 0 7952 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0651_
timestamp 1698431365
transform -1 0 9072 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0652_
timestamp 1698431365
transform -1 0 10752 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0653_
timestamp 1698431365
transform 1 0 7616 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0654_
timestamp 1698431365
transform 1 0 7616 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0655_
timestamp 1698431365
transform 1 0 11536 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0656_
timestamp 1698431365
transform 1 0 21952 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0657_
timestamp 1698431365
transform 1 0 13328 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0658_
timestamp 1698431365
transform 1 0 13440 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0659_
timestamp 1698431365
transform 1 0 15008 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0660_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0661_
timestamp 1698431365
transform -1 0 14560 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0662_
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0663_
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0664_
timestamp 1698431365
transform -1 0 30128 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0665_
timestamp 1698431365
transform -1 0 34944 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0666_
timestamp 1698431365
transform -1 0 26656 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0667_
timestamp 1698431365
transform -1 0 31024 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0668_
timestamp 1698431365
transform 1 0 29680 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0669_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26992 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0670_
timestamp 1698431365
transform 1 0 6272 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0671_
timestamp 1698431365
transform -1 0 19040 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0672_
timestamp 1698431365
transform -1 0 17920 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0673_
timestamp 1698431365
transform 1 0 9408 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0674_
timestamp 1698431365
transform -1 0 11760 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0675_
timestamp 1698431365
transform 1 0 13552 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0676_
timestamp 1698431365
transform -1 0 14112 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0677_
timestamp 1698431365
transform 1 0 11088 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0678_
timestamp 1698431365
transform 1 0 8736 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0679_
timestamp 1698431365
transform 1 0 12432 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0680_
timestamp 1698431365
transform 1 0 14112 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0681_
timestamp 1698431365
transform 1 0 34272 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0682_
timestamp 1698431365
transform -1 0 31696 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0683_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28112 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0684_
timestamp 1698431365
transform 1 0 18032 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0685_
timestamp 1698431365
transform 1 0 18928 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0686_
timestamp 1698431365
transform 1 0 25200 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0687_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20272 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0688_
timestamp 1698431365
transform -1 0 13104 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0689_
timestamp 1698431365
transform -1 0 14672 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0690_
timestamp 1698431365
transform 1 0 21280 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0691_
timestamp 1698431365
transform 1 0 6608 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0692_
timestamp 1698431365
transform 1 0 8288 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0693_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8512 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0694_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8960 0 1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0695_
timestamp 1698431365
transform 1 0 22400 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0696_
timestamp 1698431365
transform 1 0 21504 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0697_
timestamp 1698431365
transform 1 0 23968 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0698_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23744 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0699_
timestamp 1698431365
transform -1 0 23632 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0700_
timestamp 1698431365
transform 1 0 26656 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0701_
timestamp 1698431365
transform 1 0 27888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0702_
timestamp 1698431365
transform -1 0 22624 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0703_
timestamp 1698431365
transform -1 0 21840 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0704_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0705_
timestamp 1698431365
transform -1 0 23632 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0706_
timestamp 1698431365
transform -1 0 22624 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0707_
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0708_
timestamp 1698431365
transform -1 0 16576 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0709_
timestamp 1698431365
transform 1 0 16576 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0710_
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0711_
timestamp 1698431365
transform -1 0 10752 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0712_
timestamp 1698431365
transform 1 0 15008 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0713_
timestamp 1698431365
transform 1 0 13104 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0714_
timestamp 1698431365
transform 1 0 10192 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0715_
timestamp 1698431365
transform -1 0 10192 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0716_
timestamp 1698431365
transform -1 0 7840 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0717_
timestamp 1698431365
transform -1 0 5936 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0718_
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0719_
timestamp 1698431365
transform -1 0 6272 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0720_
timestamp 1698431365
transform 1 0 6608 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0721_
timestamp 1698431365
transform 1 0 8736 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0722_
timestamp 1698431365
transform -1 0 31248 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0723_
timestamp 1698431365
transform -1 0 39648 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0724_
timestamp 1698431365
transform -1 0 38304 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0725_
timestamp 1698431365
transform -1 0 36624 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0726_
timestamp 1698431365
transform 1 0 35728 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0727_
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0728_
timestamp 1698431365
transform -1 0 29904 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0729_
timestamp 1698431365
transform -1 0 30128 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0730_
timestamp 1698431365
transform -1 0 23408 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0731_
timestamp 1698431365
transform -1 0 22624 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0732_
timestamp 1698431365
transform -1 0 28784 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0733_
timestamp 1698431365
transform 1 0 28000 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0734_
timestamp 1698431365
transform -1 0 30800 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0735_
timestamp 1698431365
transform 1 0 18704 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0736_
timestamp 1698431365
transform -1 0 30352 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0737_
timestamp 1698431365
transform -1 0 31472 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0738_
timestamp 1698431365
transform 1 0 28784 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0739_
timestamp 1698431365
transform 1 0 26768 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0740_
timestamp 1698431365
transform 1 0 34160 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0741_
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0742_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38752 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0743_
timestamp 1698431365
transform 1 0 36064 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0744_
timestamp 1698431365
transform 1 0 36848 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0745_
timestamp 1698431365
transform -1 0 36176 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0746_
timestamp 1698431365
transform 1 0 29232 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0747_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29232 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0748_
timestamp 1698431365
transform 1 0 27440 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0749_
timestamp 1698431365
transform 1 0 26544 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0750_
timestamp 1698431365
transform -1 0 26768 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0751_
timestamp 1698431365
transform 1 0 27888 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0752_
timestamp 1698431365
transform -1 0 30240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0753_
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0754_
timestamp 1698431365
transform -1 0 37520 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0755_
timestamp 1698431365
transform 1 0 28672 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0756_
timestamp 1698431365
transform -1 0 29456 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0757_
timestamp 1698431365
transform -1 0 30912 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0758_
timestamp 1698431365
transform -1 0 39536 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0759_
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0760_
timestamp 1698431365
transform 1 0 32144 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0761_
timestamp 1698431365
transform -1 0 30352 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0762_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30352 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0763_
timestamp 1698431365
transform 1 0 22624 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0764_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0765_
timestamp 1698431365
transform -1 0 25760 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0766_
timestamp 1698431365
transform 1 0 26096 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0767_
timestamp 1698431365
transform -1 0 31920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0768_
timestamp 1698431365
transform -1 0 32704 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0769_
timestamp 1698431365
transform -1 0 31472 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0770_
timestamp 1698431365
transform -1 0 32032 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0771_
timestamp 1698431365
transform 1 0 30352 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0772_
timestamp 1698431365
transform -1 0 24640 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0773_
timestamp 1698431365
transform 1 0 14560 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0774_
timestamp 1698431365
transform 1 0 33264 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0775_
timestamp 1698431365
transform -1 0 34832 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0776_
timestamp 1698431365
transform 1 0 28112 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0777_
timestamp 1698431365
transform 1 0 33040 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0778_
timestamp 1698431365
transform -1 0 35392 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0779_
timestamp 1698431365
transform -1 0 33936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0780_
timestamp 1698431365
transform 1 0 31808 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0781_
timestamp 1698431365
transform -1 0 32144 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0782_
timestamp 1698431365
transform -1 0 32032 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0783_
timestamp 1698431365
transform 1 0 31584 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0784_
timestamp 1698431365
transform 1 0 32144 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0785_
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0786_
timestamp 1698431365
transform 1 0 32032 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0787_
timestamp 1698431365
transform 1 0 33152 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0788_
timestamp 1698431365
transform 1 0 20048 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0789_
timestamp 1698431365
transform 1 0 35392 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0790_
timestamp 1698431365
transform -1 0 35392 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0791_
timestamp 1698431365
transform 1 0 33488 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0792_
timestamp 1698431365
transform 1 0 34720 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0793_
timestamp 1698431365
transform 1 0 33040 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0794_
timestamp 1698431365
transform -1 0 34720 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0795_
timestamp 1698431365
transform -1 0 34496 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0796_
timestamp 1698431365
transform 1 0 31472 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0797_
timestamp 1698431365
transform 1 0 32032 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0798_
timestamp 1698431365
transform 1 0 32928 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0799_
timestamp 1698431365
transform 1 0 31808 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0800_
timestamp 1698431365
transform -1 0 32368 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0801_
timestamp 1698431365
transform -1 0 38528 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0802_
timestamp 1698431365
transform 1 0 35728 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0803_
timestamp 1698431365
transform 1 0 33936 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0804_
timestamp 1698431365
transform 1 0 36064 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0805_
timestamp 1698431365
transform 1 0 38416 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0806_
timestamp 1698431365
transform 1 0 38416 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0807_
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0808_
timestamp 1698431365
transform 1 0 37296 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0809_
timestamp 1698431365
transform -1 0 39424 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0810_
timestamp 1698431365
transform -1 0 19040 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0811_
timestamp 1698431365
transform 1 0 34832 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0812_
timestamp 1698431365
transform -1 0 37856 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0813_
timestamp 1698431365
transform 1 0 38640 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0814_
timestamp 1698431365
transform -1 0 38864 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0815_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37296 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0816_
timestamp 1698431365
transform -1 0 36064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0817_
timestamp 1698431365
transform -1 0 35728 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0818_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0819_
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0820_
timestamp 1698431365
transform -1 0 38192 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0821_
timestamp 1698431365
transform 1 0 36848 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0822_
timestamp 1698431365
transform -1 0 39088 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0823_
timestamp 1698431365
transform -1 0 37856 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0824_
timestamp 1698431365
transform -1 0 38528 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0825_
timestamp 1698431365
transform -1 0 36624 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0826_
timestamp 1698431365
transform 1 0 29792 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0827_
timestamp 1698431365
transform -1 0 32144 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0828_
timestamp 1698431365
transform 1 0 31584 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0829_
timestamp 1698431365
transform -1 0 24640 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0830_
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0831_
timestamp 1698431365
transform 1 0 35616 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0832_
timestamp 1698431365
transform -1 0 38192 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0833_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0834_
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0835_
timestamp 1698431365
transform 1 0 33152 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0836_
timestamp 1698431365
transform -1 0 39536 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0837_
timestamp 1698431365
transform 1 0 36960 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0838_
timestamp 1698431365
transform -1 0 38416 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0839_
timestamp 1698431365
transform -1 0 39312 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0840_
timestamp 1698431365
transform -1 0 38416 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0841_
timestamp 1698431365
transform -1 0 38192 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0842_
timestamp 1698431365
transform -1 0 36624 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0843_
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0844_
timestamp 1698431365
transform -1 0 37296 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0845_
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0846_
timestamp 1698431365
transform -1 0 36512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0847_
timestamp 1698431365
transform 1 0 37296 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0848_
timestamp 1698431365
transform -1 0 33712 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0849_
timestamp 1698431365
transform -1 0 39536 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0850_
timestamp 1698431365
transform 1 0 36624 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0851_
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0852_
timestamp 1698431365
transform -1 0 33936 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0853_
timestamp 1698431365
transform 1 0 34944 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0854_
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0855_
timestamp 1698431365
transform -1 0 38192 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0856_
timestamp 1698431365
transform -1 0 36624 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0857_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0858_
timestamp 1698431365
transform -1 0 35280 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0859_
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0860_
timestamp 1698431365
transform 1 0 34944 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0861_
timestamp 1698431365
transform 1 0 35280 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0862_
timestamp 1698431365
transform -1 0 32144 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0863_
timestamp 1698431365
transform -1 0 33488 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0864_
timestamp 1698431365
transform 1 0 31024 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0865_
timestamp 1698431365
transform 1 0 30128 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0866_
timestamp 1698431365
transform -1 0 31584 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0867_
timestamp 1698431365
transform -1 0 28784 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0868_
timestamp 1698431365
transform 1 0 29680 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0869_
timestamp 1698431365
transform -1 0 29456 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0870_
timestamp 1698431365
transform -1 0 32368 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0871_
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0872_
timestamp 1698431365
transform -1 0 32704 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0873_
timestamp 1698431365
transform 1 0 31808 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0874_
timestamp 1698431365
transform -1 0 31696 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0875_
timestamp 1698431365
transform -1 0 31808 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0876_
timestamp 1698431365
transform 1 0 32368 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0877_
timestamp 1698431365
transform -1 0 20944 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0878_
timestamp 1698431365
transform 1 0 29456 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0879_
timestamp 1698431365
transform -1 0 30576 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0880_
timestamp 1698431365
transform -1 0 29232 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0881_
timestamp 1698431365
transform -1 0 26880 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0882_
timestamp 1698431365
transform -1 0 25872 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0883_
timestamp 1698431365
transform -1 0 23520 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0884_
timestamp 1698431365
transform -1 0 23184 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0885_
timestamp 1698431365
transform 1 0 21504 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0886_
timestamp 1698431365
transform -1 0 24640 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0887_
timestamp 1698431365
transform 1 0 19376 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0888_
timestamp 1698431365
transform 1 0 21616 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0889_
timestamp 1698431365
transform 1 0 23632 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0890_
timestamp 1698431365
transform -1 0 25984 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0891_
timestamp 1698431365
transform -1 0 24864 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0892_
timestamp 1698431365
transform -1 0 23072 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0893_
timestamp 1698431365
transform -1 0 22176 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0894_
timestamp 1698431365
transform 1 0 21280 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0895_
timestamp 1698431365
transform 1 0 22176 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0896_
timestamp 1698431365
transform 1 0 19488 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0897_
timestamp 1698431365
transform -1 0 22288 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0898_
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0899_
timestamp 1698431365
transform 1 0 22176 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0900_
timestamp 1698431365
transform -1 0 20832 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0901_
timestamp 1698431365
transform -1 0 19824 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0902_
timestamp 1698431365
transform 1 0 16352 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0903_
timestamp 1698431365
transform -1 0 20384 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0904_
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0905_
timestamp 1698431365
transform 1 0 14448 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0906_
timestamp 1698431365
transform -1 0 16800 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0907_
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0908_
timestamp 1698431365
transform -1 0 18256 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0909_
timestamp 1698431365
transform -1 0 17920 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0910_
timestamp 1698431365
transform 1 0 17920 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0911_
timestamp 1698431365
transform -1 0 19152 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0912_
timestamp 1698431365
transform -1 0 19152 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0913_
timestamp 1698431365
transform 1 0 11760 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0914_
timestamp 1698431365
transform 1 0 14672 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0915_
timestamp 1698431365
transform -1 0 18704 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0916_
timestamp 1698431365
transform -1 0 17696 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0917_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0918_
timestamp 1698431365
transform -1 0 17696 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0919_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0920_
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0921_
timestamp 1698431365
transform 1 0 17808 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0922_
timestamp 1698431365
transform -1 0 20048 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0923_
timestamp 1698431365
transform -1 0 20832 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0924_
timestamp 1698431365
transform -1 0 20832 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0925_
timestamp 1698431365
transform 1 0 19376 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0926_
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0927_
timestamp 1698431365
transform -1 0 15344 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0928_
timestamp 1698431365
transform 1 0 12432 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0929_
timestamp 1698431365
transform 1 0 15456 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0930_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13776 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0931_
timestamp 1698431365
transform 1 0 12544 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0932_
timestamp 1698431365
transform 1 0 13216 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0933_
timestamp 1698431365
transform 1 0 12096 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0934_
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0935_
timestamp 1698431365
transform -1 0 12432 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0936_
timestamp 1698431365
transform 1 0 12320 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0937_
timestamp 1698431365
transform 1 0 10304 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0938_
timestamp 1698431365
transform 1 0 11088 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0939_
timestamp 1698431365
transform -1 0 14224 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0940_
timestamp 1698431365
transform -1 0 14672 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0941_
timestamp 1698431365
transform 1 0 12544 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0942_
timestamp 1698431365
transform -1 0 14896 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0943_
timestamp 1698431365
transform -1 0 12544 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0944_
timestamp 1698431365
transform -1 0 17920 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0945_
timestamp 1698431365
transform 1 0 12992 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0946_
timestamp 1698431365
transform 1 0 14448 0 -1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0947_
timestamp 1698431365
transform -1 0 15120 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0948_
timestamp 1698431365
transform -1 0 18592 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0949_
timestamp 1698431365
transform 1 0 16016 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0950_
timestamp 1698431365
transform 1 0 15904 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0951_
timestamp 1698431365
transform 1 0 16912 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0952_
timestamp 1698431365
transform 1 0 16912 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0953_
timestamp 1698431365
transform -1 0 18480 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0954_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _0955_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0956_
timestamp 1698431365
transform -1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0957_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25872 0 1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0958_
timestamp 1698431365
transform 1 0 25200 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0959_
timestamp 1698431365
transform 1 0 26432 0 -1 10976
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0960_
timestamp 1698431365
transform 1 0 22848 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _0961_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25200 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0962_
timestamp 1698431365
transform 1 0 24528 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0963_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25200 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0964_
timestamp 1698431365
transform 1 0 25648 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0965_
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0966_
timestamp 1698431365
transform -1 0 33264 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0967_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0968_
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0969_
timestamp 1698431365
transform 1 0 35504 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0970_
timestamp 1698431365
transform -1 0 37744 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0971_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0972_
timestamp 1698431365
transform -1 0 33936 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0973_
timestamp 1698431365
transform -1 0 31920 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0974_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0975_
timestamp 1698431365
transform -1 0 12320 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0976_
timestamp 1698431365
transform 1 0 7728 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0977_
timestamp 1698431365
transform -1 0 12320 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0978_
timestamp 1698431365
transform -1 0 12208 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0979_
timestamp 1698431365
transform -1 0 10864 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0980_
timestamp 1698431365
transform -1 0 10080 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0981_
timestamp 1698431365
transform -1 0 8848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0982_
timestamp 1698431365
transform 1 0 7392 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0983_
timestamp 1698431365
transform 1 0 8848 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0984_
timestamp 1698431365
transform 1 0 10192 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0985_
timestamp 1698431365
transform -1 0 11648 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0986_
timestamp 1698431365
transform 1 0 6944 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0987_
timestamp 1698431365
transform 1 0 9744 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0988_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0989_
timestamp 1698431365
transform 1 0 8736 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0990_
timestamp 1698431365
transform 1 0 10752 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0991_
timestamp 1698431365
transform 1 0 9968 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0992_
timestamp 1698431365
transform 1 0 8960 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0993_
timestamp 1698431365
transform 1 0 5936 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0994_
timestamp 1698431365
transform 1 0 8064 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0995_
timestamp 1698431365
transform 1 0 10192 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0996_
timestamp 1698431365
transform -1 0 12544 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0997_
timestamp 1698431365
transform 1 0 7616 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0998_
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0999_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1000_
timestamp 1698431365
transform 1 0 10976 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1001_
timestamp 1698431365
transform -1 0 14784 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1002_
timestamp 1698431365
transform -1 0 14224 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1003_
timestamp 1698431365
transform -1 0 14560 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1004_
timestamp 1698431365
transform -1 0 29568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1005_
timestamp 1698431365
transform 1 0 28112 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1006_
timestamp 1698431365
transform -1 0 30688 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1007_
timestamp 1698431365
transform 1 0 31024 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1008_
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1009_
timestamp 1698431365
transform -1 0 14336 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1010_
timestamp 1698431365
transform 1 0 15568 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1011_
timestamp 1698431365
transform -1 0 26544 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1012_
timestamp 1698431365
transform 1 0 24864 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1013_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1014_
timestamp 1698431365
transform 1 0 26432 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1015_
timestamp 1698431365
transform 1 0 31136 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1016_
timestamp 1698431365
transform 1 0 30688 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1017_
timestamp 1698431365
transform -1 0 32704 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1018_
timestamp 1698431365
transform 1 0 25760 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1019_
timestamp 1698431365
transform -1 0 32032 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1020_
timestamp 1698431365
transform -1 0 30576 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1021_
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1022_
timestamp 1698431365
transform -1 0 28784 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1023_
timestamp 1698431365
transform -1 0 27776 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1024_
timestamp 1698431365
transform 1 0 27104 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1025_
timestamp 1698431365
transform 1 0 26992 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1026_
timestamp 1698431365
transform 1 0 27888 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1027_
timestamp 1698431365
transform -1 0 27552 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1028_
timestamp 1698431365
transform 1 0 26320 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1029_
timestamp 1698431365
transform 1 0 25088 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1030_
timestamp 1698431365
transform -1 0 27664 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1031_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1032_
timestamp 1698431365
transform 1 0 28000 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1033_
timestamp 1698431365
transform 1 0 29568 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1034_
timestamp 1698431365
transform 1 0 29568 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1035_
timestamp 1698431365
transform 1 0 27664 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1036_
timestamp 1698431365
transform 1 0 28784 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1037_
timestamp 1698431365
transform -1 0 29344 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1038_
timestamp 1698431365
transform 1 0 26544 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1039_
timestamp 1698431365
transform -1 0 27888 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1040_
timestamp 1698431365
transform -1 0 4592 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1041_
timestamp 1698431365
transform -1 0 11872 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1042_
timestamp 1698431365
transform -1 0 3696 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1043_
timestamp 1698431365
transform 1 0 2688 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1044_
timestamp 1698431365
transform -1 0 4256 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1045_
timestamp 1698431365
transform -1 0 2912 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1046_
timestamp 1698431365
transform 1 0 16240 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1047_
timestamp 1698431365
transform -1 0 4592 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1048_
timestamp 1698431365
transform 1 0 4592 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1049_
timestamp 1698431365
transform -1 0 4144 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1050_
timestamp 1698431365
transform -1 0 7840 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1051_
timestamp 1698431365
transform 1 0 3808 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1052_
timestamp 1698431365
transform -1 0 3472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1053_
timestamp 1698431365
transform -1 0 6384 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1054_
timestamp 1698431365
transform 1 0 4032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1055_
timestamp 1698431365
transform -1 0 4256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1056_
timestamp 1698431365
transform -1 0 4256 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1057_
timestamp 1698431365
transform -1 0 3360 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1058_
timestamp 1698431365
transform 1 0 8176 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1059_
timestamp 1698431365
transform -1 0 6832 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1060_
timestamp 1698431365
transform 1 0 7728 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1061_
timestamp 1698431365
transform -1 0 5488 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1062_
timestamp 1698431365
transform -1 0 6160 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1063_
timestamp 1698431365
transform -1 0 5040 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1064_
timestamp 1698431365
transform -1 0 4144 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1065_
timestamp 1698431365
transform -1 0 2688 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1066_
timestamp 1698431365
transform 1 0 3584 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1067_
timestamp 1698431365
transform -1 0 5488 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1068_
timestamp 1698431365
transform -1 0 3696 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1069_
timestamp 1698431365
transform 1 0 37968 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1070_
timestamp 1698431365
transform -1 0 38192 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1071_
timestamp 1698431365
transform -1 0 37408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1072_
timestamp 1698431365
transform -1 0 38192 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1073_
timestamp 1698431365
transform -1 0 36512 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1074_
timestamp 1698431365
transform -1 0 34160 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1075_
timestamp 1698431365
transform -1 0 32368 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1076_
timestamp 1698431365
transform 1 0 15344 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1077_
timestamp 1698431365
transform -1 0 14784 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1078_
timestamp 1698431365
transform -1 0 18592 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1079_
timestamp 1698431365
transform -1 0 19600 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1080_
timestamp 1698431365
transform -1 0 18144 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1081_
timestamp 1698431365
transform 1 0 16912 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1082_
timestamp 1698431365
transform -1 0 19600 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1083_
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1084_
timestamp 1698431365
transform 1 0 17584 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1085_
timestamp 1698431365
transform 1 0 18480 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1086_
timestamp 1698431365
transform -1 0 18480 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1087_
timestamp 1698431365
transform -1 0 20160 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1088_
timestamp 1698431365
transform -1 0 20048 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1089_
timestamp 1698431365
transform -1 0 19488 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1090_
timestamp 1698431365
transform -1 0 19264 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1091_
timestamp 1698431365
transform -1 0 19040 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1092_
timestamp 1698431365
transform -1 0 19376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1093_
timestamp 1698431365
transform -1 0 18704 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1094_
timestamp 1698431365
transform -1 0 18368 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1095_
timestamp 1698431365
transform -1 0 14784 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1096_
timestamp 1698431365
transform -1 0 18592 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1097_
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1098_
timestamp 1698431365
transform -1 0 19824 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1099_
timestamp 1698431365
transform -1 0 18592 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1100_
timestamp 1698431365
transform 1 0 19264 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1101_
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1102_
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1103_
timestamp 1698431365
transform 1 0 19600 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1104_
timestamp 1698431365
transform -1 0 20384 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1105_
timestamp 1698431365
transform 1 0 22288 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1106_
timestamp 1698431365
transform 1 0 23072 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1107_
timestamp 1698431365
transform 1 0 23744 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1108_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1109_
timestamp 1698431365
transform -1 0 22288 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1110_
timestamp 1698431365
transform -1 0 24192 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1111_
timestamp 1698431365
transform 1 0 23072 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1112_
timestamp 1698431365
transform 1 0 24192 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1113_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22736 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1114_
timestamp 1698431365
transform -1 0 17248 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1115_
timestamp 1698431365
transform 1 0 9408 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1116_
timestamp 1698431365
transform 1 0 1680 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1117_
timestamp 1698431365
transform -1 0 8736 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1118_
timestamp 1698431365
transform 1 0 20944 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1119_
timestamp 1698431365
transform -1 0 32368 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1120_
timestamp 1698431365
transform 1 0 25312 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1121_
timestamp 1698431365
transform 1 0 23744 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1122_
timestamp 1698431365
transform 1 0 22624 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1123_
timestamp 1698431365
transform 1 0 32480 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1124_
timestamp 1698431365
transform -1 0 34720 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1125_
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1126_
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1127_
timestamp 1698431365
transform 1 0 32704 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1128_
timestamp 1698431365
transform 1 0 36512 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1129_
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1130_
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1131_
timestamp 1698431365
transform -1 0 37520 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1132_
timestamp 1698431365
transform 1 0 28000 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1133_
timestamp 1698431365
transform -1 0 34944 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1134_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1135_
timestamp 1698431365
transform 1 0 20384 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1136_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28560 0 -1 37632
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1137_
timestamp 1698431365
transform -1 0 24416 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1138_
timestamp 1698431365
transform 1 0 15568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1139_
timestamp 1698431365
transform 1 0 5936 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1140_
timestamp 1698431365
transform -1 0 23296 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1141_
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1142_
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1143_
timestamp 1698431365
transform 1 0 2688 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1144_
timestamp 1698431365
transform 1 0 15904 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1145_
timestamp 1698431365
transform -1 0 16576 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1146_
timestamp 1698431365
transform 1 0 32144 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1147_
timestamp 1698431365
transform 1 0 15792 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1148_
timestamp 1698431365
transform 1 0 26880 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1149_
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1150_
timestamp 1698431365
transform 1 0 1792 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1151_
timestamp 1698431365
transform 1 0 2128 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1152_
timestamp 1698431365
transform 1 0 1680 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1153_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1154_
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1155_
timestamp 1698431365
transform 1 0 8176 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1156_
timestamp 1698431365
transform 1 0 3696 0 -1 28224
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1157_
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1158_
timestamp 1698431365
transform 1 0 1680 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1159_
timestamp 1698431365
transform -1 0 15568 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1160_
timestamp 1698431365
transform 1 0 17696 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1161_
timestamp 1698431365
transform -1 0 19600 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1162_
timestamp 1698431365
transform -1 0 16800 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1163_
timestamp 1698431365
transform -1 0 15792 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1164_
timestamp 1698431365
transform 1 0 16016 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1165_
timestamp 1698431365
transform 1 0 17696 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1166_
timestamp 1698431365
transform 1 0 19824 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1167_
timestamp 1698431365
transform 1 0 22624 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1168_
timestamp 1698431365
transform 1 0 21504 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1169_
timestamp 1698431365
transform 1 0 26544 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1175_
timestamp 1698431365
transform 1 0 4480 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0554__A2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0570__A1
timestamp 1698431365
transform 1 0 15904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0574__A1
timestamp 1698431365
transform 1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0576__A1
timestamp 1698431365
transform 1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0584__I
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0585__A1
timestamp 1698431365
transform -1 0 20048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0589__A1
timestamp 1698431365
transform 1 0 19824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0615__A1
timestamp 1698431365
transform 1 0 20720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0626__A1
timestamp 1698431365
transform 1 0 15792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0649__A1
timestamp 1698431365
transform 1 0 12544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0673__I
timestamp 1698431365
transform 1 0 10528 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0688__I
timestamp 1698431365
transform -1 0 12768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0690__I
timestamp 1698431365
transform -1 0 20832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0696__A2
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0700__A1
timestamp 1698431365
transform -1 0 27888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A2
timestamp 1698431365
transform 1 0 22848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0703__A1
timestamp 1698431365
transform 1 0 22064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0705__A1
timestamp 1698431365
transform -1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0706__I
timestamp 1698431365
transform -1 0 22848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0708__A2
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0709__A3
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0710__A1
timestamp 1698431365
transform 1 0 18368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0714__B
timestamp 1698431365
transform 1 0 11648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0718__A1
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0721__A1
timestamp 1698431365
transform -1 0 9632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0730__A1
timestamp 1698431365
transform 1 0 23632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0730__B
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0734__A1
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0734__B
timestamp 1698431365
transform 1 0 31696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0736__B
timestamp 1698431365
transform 1 0 29232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0747__C
timestamp 1698431365
transform 1 0 30128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0749__A2
timestamp 1698431365
transform 1 0 26320 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0750__A1
timestamp 1698431365
transform 1 0 25648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0752__I
timestamp 1698431365
transform 1 0 30912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0753__A1
timestamp 1698431365
transform 1 0 30576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0764__B2
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__A1
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0772__A1
timestamp 1698431365
transform 1 0 23744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__I
timestamp 1698431365
transform 1 0 33040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__B2
timestamp 1698431365
transform 1 0 31248 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0787__A1
timestamp 1698431365
transform 1 0 33824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0798__B
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0800__A1
timestamp 1698431365
transform 1 0 31584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0810__I
timestamp 1698431365
transform 1 0 19264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0811__I
timestamp 1698431365
transform 1 0 34608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0812__B2
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0813__A1
timestamp 1698431365
transform -1 0 33488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0823__B2
timestamp 1698431365
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0824__A1
timestamp 1698431365
transform 1 0 39312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__A2
timestamp 1698431365
transform 1 0 30912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__B
timestamp 1698431365
transform 1 0 30352 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__A2
timestamp 1698431365
transform 1 0 31360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A1
timestamp 1698431365
transform 1 0 24864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__A2
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__B2
timestamp 1698431365
transform 1 0 35952 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0834__A1
timestamp 1698431365
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0835__I
timestamp 1698431365
transform -1 0 33488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__A2
timestamp 1698431365
transform 1 0 35168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__B2
timestamp 1698431365
transform -1 0 35616 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__I
timestamp 1698431365
transform 1 0 33040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__A1
timestamp 1698431365
transform -1 0 28224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__A2
timestamp 1698431365
transform 1 0 29456 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__A1
timestamp 1698431365
transform -1 0 29456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__B
timestamp 1698431365
transform 1 0 30576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__I
timestamp 1698431365
transform -1 0 20272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0884__A1
timestamp 1698431365
transform 1 0 23856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0884__A2
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0884__B
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__A1
timestamp 1698431365
transform 1 0 22624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__A2
timestamp 1698431365
transform 1 0 23072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__A2
timestamp 1698431365
transform 1 0 23184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__A1
timestamp 1698431365
transform -1 0 23632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A1
timestamp 1698431365
transform 1 0 26208 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A2
timestamp 1698431365
transform 1 0 22176 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0898__A1
timestamp 1698431365
transform 1 0 23072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__A2
timestamp 1698431365
transform 1 0 20384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__A2
timestamp 1698431365
transform -1 0 18704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A1
timestamp 1698431365
transform 1 0 19040 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A2
timestamp 1698431365
transform 1 0 17696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__B
timestamp 1698431365
transform -1 0 16800 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0922__B
timestamp 1698431365
transform 1 0 18256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__A2
timestamp 1698431365
transform -1 0 19376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0926__B
timestamp 1698431365
transform 1 0 20944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0927__I
timestamp 1698431365
transform 1 0 15344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__B
timestamp 1698431365
transform 1 0 14336 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__A1
timestamp 1698431365
transform -1 0 11760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__A1
timestamp 1698431365
transform 1 0 12544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0944__A2
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__A1
timestamp 1698431365
transform 1 0 18928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__B
timestamp 1698431365
transform 1 0 16688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__A1
timestamp 1698431365
transform -1 0 17920 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0965__A1
timestamp 1698431365
transform -1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__B
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__C
timestamp 1698431365
transform -1 0 19600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__A1
timestamp 1698431365
transform 1 0 12544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A2
timestamp 1698431365
transform -1 0 10528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0982__A2
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A2
timestamp 1698431365
transform 1 0 11648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__A2
timestamp 1698431365
transform -1 0 10528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__C
timestamp 1698431365
transform 1 0 14784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__A1
timestamp 1698431365
transform 1 0 30800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__A1
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A1
timestamp 1698431365
transform 1 0 30464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A1
timestamp 1698431365
transform -1 0 29792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A1
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1024__A1
timestamp 1698431365
transform 1 0 28224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1028__A1
timestamp 1698431365
transform -1 0 26320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A1
timestamp 1698431365
transform -1 0 26992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__A2
timestamp 1698431365
transform -1 0 11312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A1
timestamp 1698431365
transform -1 0 4592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A1
timestamp 1698431365
transform 1 0 3472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A1
timestamp 1698431365
transform 1 0 4256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A1
timestamp 1698431365
transform 1 0 34384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__A2
timestamp 1698431365
transform -1 0 16688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__B
timestamp 1698431365
transform 1 0 16912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698431365
transform 1 0 15568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__A1
timestamp 1698431365
transform 1 0 17920 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A2
timestamp 1698431365
transform -1 0 19824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__I
timestamp 1698431365
transform 1 0 17584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A3
timestamp 1698431365
transform -1 0 20272 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__B
timestamp 1698431365
transform 1 0 17360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A1
timestamp 1698431365
transform 1 0 18144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A1
timestamp 1698431365
transform -1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__A1
timestamp 1698431365
transform 1 0 15680 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__A1
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A1
timestamp 1698431365
transform 1 0 19264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__C
timestamp 1698431365
transform 1 0 18816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__B
timestamp 1698431365
transform 1 0 20384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__A1
timestamp 1698431365
transform 1 0 19264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__A1
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1110__C
timestamp 1698431365
transform 1 0 25088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1111__A1
timestamp 1698431365
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1113__CLK
timestamp 1698431365
transform 1 0 22960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__CLK
timestamp 1698431365
transform -1 0 17696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__CLK
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__CLK
timestamp 1698431365
transform 1 0 4928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__CLK
timestamp 1698431365
transform 1 0 8848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__CLK
timestamp 1698431365
transform -1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__CLK
timestamp 1698431365
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__CLK
timestamp 1698431365
transform -1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__CLK
timestamp 1698431365
transform 1 0 27216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__CLK
timestamp 1698431365
transform 1 0 26096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__CLK
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__CLK
timestamp 1698431365
transform 1 0 31248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__CLK
timestamp 1698431365
transform 1 0 35280 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__CLK
timestamp 1698431365
transform 1 0 36288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__CLK
timestamp 1698431365
transform -1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1128__CLK
timestamp 1698431365
transform -1 0 36512 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__CLK
timestamp 1698431365
transform 1 0 35840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1130__CLK
timestamp 1698431365
transform 1 0 36288 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__CLK
timestamp 1698431365
transform 1 0 34048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1132__CLK
timestamp 1698431365
transform 1 0 31472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__CLK
timestamp 1698431365
transform 1 0 31472 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__CLK
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__CLK
timestamp 1698431365
transform -1 0 24080 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__CLK
timestamp 1698431365
transform 1 0 28784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__CLK
timestamp 1698431365
transform 1 0 24640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__CLK
timestamp 1698431365
transform 1 0 15344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1140__CLK
timestamp 1698431365
transform 1 0 23520 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__CLK
timestamp 1698431365
transform 1 0 13552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1142__CLK
timestamp 1698431365
transform 1 0 9632 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__CLK
timestamp 1698431365
transform 1 0 5936 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__CLK
timestamp 1698431365
transform 1 0 15680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1145__CLK
timestamp 1698431365
transform 1 0 16800 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__CLK
timestamp 1698431365
transform 1 0 31920 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__CLK
timestamp 1698431365
transform 1 0 15568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__CLK
timestamp 1698431365
transform -1 0 30576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__CLK
timestamp 1698431365
transform 1 0 5264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__CLK
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__CLK
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__CLK
timestamp 1698431365
transform 1 0 11872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__CLK
timestamp 1698431365
transform 1 0 7168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__CLK
timestamp 1698431365
transform 1 0 5040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__CLK
timestamp 1698431365
transform 1 0 15232 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__CLK
timestamp 1698431365
transform 1 0 16352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1161__CLK
timestamp 1698431365
transform 1 0 19824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__CLK
timestamp 1698431365
transform 1 0 17024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__CLK
timestamp 1698431365
transform 1 0 16016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__CLK
timestamp 1698431365
transform 1 0 15792 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__CLK
timestamp 1698431365
transform 1 0 17472 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__CLK
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1167__CLK
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1168__CLK
timestamp 1698431365
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1169__CLK
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 18816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_clk_I
timestamp 1698431365
transform 1 0 16912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_clk_I
timestamp 1698431365
transform 1 0 16240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_clk_I
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_clk_I
timestamp 1698431365
transform 1 0 25984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_clk_I
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_clk_I
timestamp 1698431365
transform 1 0 15904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_clk_I
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_clk_I
timestamp 1698431365
transform -1 0 28896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold2_I
timestamp 1698431365
transform 1 0 33264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold12_I
timestamp 1698431365
transform -1 0 32032 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold13_I
timestamp 1698431365
transform -1 0 31136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold18_I
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold20_I
timestamp 1698431365
transform 1 0 38528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold21_I
timestamp 1698431365
transform -1 0 31584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 3248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output9_I
timestamp 1698431365
transform 1 0 9296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output14_I
timestamp 1698431365
transform 1 0 13216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1698431365
transform 1 0 11424 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1698431365
transform 1 0 10416 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1698431365
transform 1 0 25200 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1698431365
transform 1 0 11424 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1698431365
transform -1 0 15680 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1698431365
transform 1 0 27104 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_10 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_14 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2912 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_23
timestamp 1698431365
transform 1 0 3920 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_31
timestamp 1698431365
transform 1 0 4816 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_74
timestamp 1698431365
transform 1 0 9632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_108
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_168
timestamp 1698431365
transform 1 0 20160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_177
timestamp 1698431365
transform 1 0 21168 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_189
timestamp 1698431365
transform 1 0 22512 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_197
timestamp 1698431365
transform 1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_242
timestamp 1698431365
transform 1 0 28448 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_245 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28784 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_261
timestamp 1698431365
transform 1 0 30576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_263
timestamp 1698431365
transform 1 0 30800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_20
timestamp 1698431365
transform 1 0 3584 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_25
timestamp 1698431365
transform 1 0 4144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_27
timestamp 1698431365
transform 1 0 4368 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_34
timestamp 1698431365
transform 1 0 5152 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_74
timestamp 1698431365
transform 1 0 9632 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_127
timestamp 1698431365
transform 1 0 15568 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_135
timestamp 1698431365
transform 1 0 16464 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_146
timestamp 1698431365
transform 1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_148
timestamp 1698431365
transform 1 0 17920 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_153
timestamp 1698431365
transform 1 0 18480 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_161
timestamp 1698431365
transform 1 0 19376 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_191
timestamp 1698431365
transform 1 0 22736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195
timestamp 1698431365
transform 1 0 23184 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_243
timestamp 1698431365
transform 1 0 28560 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_254
timestamp 1698431365
transform 1 0 29792 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_262
timestamp 1698431365
transform 1 0 30688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_266
timestamp 1698431365
transform 1 0 31136 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_270
timestamp 1698431365
transform 1 0 31584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_142
timestamp 1698431365
transform 1 0 17248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_146
timestamp 1698431365
transform 1 0 17696 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_162
timestamp 1698431365
transform 1 0 19488 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_170
timestamp 1698431365
transform 1 0 20384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_183
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_187
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_195
timestamp 1698431365
transform 1 0 23184 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_199
timestamp 1698431365
transform 1 0 23632 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_229
timestamp 1698431365
transform 1 0 26992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_233
timestamp 1698431365
transform 1 0 27440 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_277
timestamp 1698431365
transform 1 0 32368 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_313
timestamp 1698431365
transform 1 0 36400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_342
timestamp 1698431365
transform 1 0 39648 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_18
timestamp 1698431365
transform 1 0 3360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_26
timestamp 1698431365
transform 1 0 4256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_30
timestamp 1698431365
transform 1 0 4704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_34
timestamp 1698431365
transform 1 0 5152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_67
timestamp 1698431365
transform 1 0 8848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_87
timestamp 1698431365
transform 1 0 11088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_95
timestamp 1698431365
transform 1 0 11984 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_99
timestamp 1698431365
transform 1 0 12432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_110
timestamp 1698431365
transform 1 0 13664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_118
timestamp 1698431365
transform 1 0 14560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_154
timestamp 1698431365
transform 1 0 18592 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_170
timestamp 1698431365
transform 1 0 20384 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_190
timestamp 1698431365
transform 1 0 22624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_194
timestamp 1698431365
transform 1 0 23072 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_202
timestamp 1698431365
transform 1 0 23968 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_218
timestamp 1698431365
transform 1 0 25760 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_234
timestamp 1698431365
transform 1 0 27552 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_238
timestamp 1698431365
transform 1 0 28000 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_251
timestamp 1698431365
transform 1 0 29456 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_267
timestamp 1698431365
transform 1 0 31248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_278
timestamp 1698431365
transform 1 0 32480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_284
timestamp 1698431365
transform 1 0 33152 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_342
timestamp 1698431365
transform 1 0 39648 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_45
timestamp 1698431365
transform 1 0 6384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_65
timestamp 1698431365
transform 1 0 8624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_73
timestamp 1698431365
transform 1 0 9520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_75
timestamp 1698431365
transform 1 0 9744 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_90
timestamp 1698431365
transform 1 0 11424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_94
timestamp 1698431365
transform 1 0 11872 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_98
timestamp 1698431365
transform 1 0 12320 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_100
timestamp 1698431365
transform 1 0 12544 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_129
timestamp 1698431365
transform 1 0 15792 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_133
timestamp 1698431365
transform 1 0 16240 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_189
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_219
timestamp 1698431365
transform 1 0 25872 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_223
timestamp 1698431365
transform 1 0 26320 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_231
timestamp 1698431365
transform 1 0 27216 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_235
timestamp 1698431365
transform 1 0 27664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_243
timestamp 1698431365
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_254
timestamp 1698431365
transform 1 0 29792 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_270
timestamp 1698431365
transform 1 0 31584 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_278
timestamp 1698431365
transform 1 0 32480 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_282
timestamp 1698431365
transform 1 0 32928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_290
timestamp 1698431365
transform 1 0 33824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_292
timestamp 1698431365
transform 1 0 34048 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_323
timestamp 1698431365
transform 1 0 37520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_33
timestamp 1698431365
transform 1 0 5040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_37
timestamp 1698431365
transform 1 0 5488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_45
timestamp 1698431365
transform 1 0 6384 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_50
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_63
timestamp 1698431365
transform 1 0 8400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_67
timestamp 1698431365
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_85
timestamp 1698431365
transform 1 0 10864 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_101
timestamp 1698431365
transform 1 0 12656 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_105
timestamp 1698431365
transform 1 0 13104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_119
timestamp 1698431365
transform 1 0 14672 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_127
timestamp 1698431365
transform 1 0 15568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_131
timestamp 1698431365
transform 1 0 16016 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_148
timestamp 1698431365
transform 1 0 17920 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_164
timestamp 1698431365
transform 1 0 19712 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_192
timestamp 1698431365
transform 1 0 22848 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_208
timestamp 1698431365
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_255
timestamp 1698431365
transform 1 0 29904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_259
timestamp 1698431365
transform 1 0 30352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_261
timestamp 1698431365
transform 1 0 30576 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_274
timestamp 1698431365
transform 1 0 32032 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_292
timestamp 1698431365
transform 1 0 34048 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_300
timestamp 1698431365
transform 1 0 34944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_302
timestamp 1698431365
transform 1 0 35168 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_6
timestamp 1698431365
transform 1 0 2016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_26
timestamp 1698431365
transform 1 0 4256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_30
timestamp 1698431365
transform 1 0 4704 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_43
timestamp 1698431365
transform 1 0 6160 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_59
timestamp 1698431365
transform 1 0 7952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_63
timestamp 1698431365
transform 1 0 8400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_65
timestamp 1698431365
transform 1 0 8624 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_70
timestamp 1698431365
transform 1 0 9184 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_86
timestamp 1698431365
transform 1 0 10976 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_94
timestamp 1698431365
transform 1 0 11872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_96
timestamp 1698431365
transform 1 0 12096 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_163
timestamp 1698431365
transform 1 0 19600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_167
timestamp 1698431365
transform 1 0 20048 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_217
timestamp 1698431365
transform 1 0 25648 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_227
timestamp 1698431365
transform 1 0 26768 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_268
timestamp 1698431365
transform 1 0 31360 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_280
timestamp 1698431365
transform 1 0 32704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_282
timestamp 1698431365
transform 1 0 32928 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_299
timestamp 1698431365
transform 1 0 34832 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_307
timestamp 1698431365
transform 1 0 35728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_309
timestamp 1698431365
transform 1 0 35952 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_330
timestamp 1698431365
transform 1 0 38304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_31
timestamp 1698431365
transform 1 0 4816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_35
timestamp 1698431365
transform 1 0 5264 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_80
timestamp 1698431365
transform 1 0 10304 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_88
timestamp 1698431365
transform 1 0 11200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_90
timestamp 1698431365
transform 1 0 11424 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_114
timestamp 1698431365
transform 1 0 14112 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_130
timestamp 1698431365
transform 1 0 15904 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698431365
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_263
timestamp 1698431365
transform 1 0 30800 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_273
timestamp 1698431365
transform 1 0 31920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_277
timestamp 1698431365
transform 1 0 32368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_298
timestamp 1698431365
transform 1 0 34720 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_315
timestamp 1698431365
transform 1 0 36624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_341
timestamp 1698431365
transform 1 0 39536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_10
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_18
timestamp 1698431365
transform 1 0 3360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_22
timestamp 1698431365
transform 1 0 3808 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_29
timestamp 1698431365
transform 1 0 4592 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_33
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_55
timestamp 1698431365
transform 1 0 7504 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_79
timestamp 1698431365
transform 1 0 10192 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_95
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_103
timestamp 1698431365
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_124
timestamp 1698431365
transform 1 0 15232 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_132
timestamp 1698431365
transform 1 0 16128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_136
timestamp 1698431365
transform 1 0 16576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_138
timestamp 1698431365
transform 1 0 16800 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_141
timestamp 1698431365
transform 1 0 17136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_145
timestamp 1698431365
transform 1 0 17584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_147
timestamp 1698431365
transform 1 0 17808 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_160
timestamp 1698431365
transform 1 0 19264 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_168
timestamp 1698431365
transform 1 0 20160 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_172
timestamp 1698431365
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_185
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_190
timestamp 1698431365
transform 1 0 22624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_204
timestamp 1698431365
transform 1 0 24192 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_220
timestamp 1698431365
transform 1 0 25984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_222
timestamp 1698431365
transform 1 0 26208 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_264
timestamp 1698431365
transform 1 0 30912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_266
timestamp 1698431365
transform 1 0 31136 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_283
timestamp 1698431365
transform 1 0 33040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_312
timestamp 1698431365
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_332
timestamp 1698431365
transform 1 0 38528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_334
timestamp 1698431365
transform 1 0 38752 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_340
timestamp 1698431365
transform 1 0 39424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_342
timestamp 1698431365
transform 1 0 39648 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_42
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_46
timestamp 1698431365
transform 1 0 6496 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_48
timestamp 1698431365
transform 1 0 6720 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_62
timestamp 1698431365
transform 1 0 8288 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_144
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_160
timestamp 1698431365
transform 1 0 19264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_162
timestamp 1698431365
transform 1 0 19488 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_165
timestamp 1698431365
transform 1 0 19824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_169
timestamp 1698431365
transform 1 0 20272 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_173
timestamp 1698431365
transform 1 0 20720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_204
timestamp 1698431365
transform 1 0 24192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_208
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_259
timestamp 1698431365
transform 1 0 30352 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_267
timestamp 1698431365
transform 1 0 31248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_271
timestamp 1698431365
transform 1 0 31696 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_292
timestamp 1698431365
transform 1 0 34048 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_296
timestamp 1698431365
transform 1 0 34496 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_298
timestamp 1698431365
transform 1 0 34720 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_339
timestamp 1698431365
transform 1 0 39312 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_79
timestamp 1698431365
transform 1 0 10192 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_87
timestamp 1698431365
transform 1 0 11088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1698431365
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_138
timestamp 1698431365
transform 1 0 16800 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_142
timestamp 1698431365
transform 1 0 17248 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_144
timestamp 1698431365
transform 1 0 17472 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_168
timestamp 1698431365
transform 1 0 20160 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_179
timestamp 1698431365
transform 1 0 21392 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_197
timestamp 1698431365
transform 1 0 23408 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_201
timestamp 1698431365
transform 1 0 23856 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_209
timestamp 1698431365
transform 1 0 24752 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_236
timestamp 1698431365
transform 1 0 27776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_238
timestamp 1698431365
transform 1 0 28000 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_267
timestamp 1698431365
transform 1 0 31248 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_269
timestamp 1698431365
transform 1 0 31472 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_281
timestamp 1698431365
transform 1 0 32816 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_297
timestamp 1698431365
transform 1 0 34608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_301
timestamp 1698431365
transform 1 0 35056 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_303
timestamp 1698431365
transform 1 0 35280 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_310
timestamp 1698431365
transform 1 0 36064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_312
timestamp 1698431365
transform 1 0 36288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_336
timestamp 1698431365
transform 1 0 38976 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_340
timestamp 1698431365
transform 1 0 39424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_342
timestamp 1698431365
transform 1 0 39648 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_6
timestamp 1698431365
transform 1 0 2016 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_36
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_40
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_42
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_49
timestamp 1698431365
transform 1 0 6832 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_53
timestamp 1698431365
transform 1 0 7280 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_55
timestamp 1698431365
transform 1 0 7504 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_84
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_92
timestamp 1698431365
transform 1 0 11648 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_102
timestamp 1698431365
transform 1 0 12768 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_134
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_167
timestamp 1698431365
transform 1 0 20048 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_175
timestamp 1698431365
transform 1 0 20944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_177
timestamp 1698431365
transform 1 0 21168 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_184
timestamp 1698431365
transform 1 0 21952 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_188
timestamp 1698431365
transform 1 0 22400 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_204
timestamp 1698431365
transform 1 0 24192 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_261
timestamp 1698431365
transform 1 0 30576 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_277
timestamp 1698431365
transform 1 0 32368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_296
timestamp 1698431365
transform 1 0 34496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_304
timestamp 1698431365
transform 1 0 35392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_306
timestamp 1698431365
transform 1 0 35616 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_313
timestamp 1698431365
transform 1 0 36400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_327
timestamp 1698431365
transform 1 0 37968 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_45
timestamp 1698431365
transform 1 0 6384 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_49
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_55
timestamp 1698431365
transform 1 0 7504 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_64
timestamp 1698431365
transform 1 0 8512 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_80
timestamp 1698431365
transform 1 0 10304 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_147
timestamp 1698431365
transform 1 0 17808 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_151
timestamp 1698431365
transform 1 0 18256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_167
timestamp 1698431365
transform 1 0 20048 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_203
timestamp 1698431365
transform 1 0 24080 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_259
timestamp 1698431365
transform 1 0 30352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_303
timestamp 1698431365
transform 1 0 35280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_334
timestamp 1698431365
transform 1 0 38752 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_342
timestamp 1698431365
transform 1 0 39648 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_32
timestamp 1698431365
transform 1 0 4928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_36
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_131
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_135
timestamp 1698431365
transform 1 0 16464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_146
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_155
timestamp 1698431365
transform 1 0 18704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_163
timestamp 1698431365
transform 1 0 19600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_167
timestamp 1698431365
transform 1 0 20048 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_183
timestamp 1698431365
transform 1 0 21840 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_187
timestamp 1698431365
transform 1 0 22288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_193
timestamp 1698431365
transform 1 0 22960 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_272
timestamp 1698431365
transform 1 0 31808 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_288
timestamp 1698431365
transform 1 0 33600 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_316
timestamp 1698431365
transform 1 0 36736 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_337
timestamp 1698431365
transform 1 0 39088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_341
timestamp 1698431365
transform 1 0 39536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_10
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_14
timestamp 1698431365
transform 1 0 2912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_16
timestamp 1698431365
transform 1 0 3136 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_25
timestamp 1698431365
transform 1 0 4144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_51
timestamp 1698431365
transform 1 0 7056 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_83
timestamp 1698431365
transform 1 0 10640 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_87
timestamp 1698431365
transform 1 0 11088 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_125
timestamp 1698431365
transform 1 0 15344 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_141
timestamp 1698431365
transform 1 0 17136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_170
timestamp 1698431365
transform 1 0 20384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_187
timestamp 1698431365
transform 1 0 22288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_194
timestamp 1698431365
transform 1 0 23072 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_198
timestamp 1698431365
transform 1 0 23520 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_203
timestamp 1698431365
transform 1 0 24080 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_219
timestamp 1698431365
transform 1 0 25872 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_222
timestamp 1698431365
transform 1 0 26208 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_238
timestamp 1698431365
transform 1 0 28000 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_242
timestamp 1698431365
transform 1 0 28448 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_269
timestamp 1698431365
transform 1 0 31472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_273
timestamp 1698431365
transform 1 0 31920 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_305
timestamp 1698431365
transform 1 0 35504 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_313
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_10
timestamp 1698431365
transform 1 0 2464 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_46
timestamp 1698431365
transform 1 0 6496 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_76
timestamp 1698431365
transform 1 0 9856 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_129
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_171
timestamp 1698431365
transform 1 0 20496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_175
timestamp 1698431365
transform 1 0 20944 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_191
timestamp 1698431365
transform 1 0 22736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698431365
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_244
timestamp 1698431365
transform 1 0 28672 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_248
timestamp 1698431365
transform 1 0 29120 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_250
timestamp 1698431365
transform 1 0 29344 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_257
timestamp 1698431365
transform 1 0 30128 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_263
timestamp 1698431365
transform 1 0 30800 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_269
timestamp 1698431365
transform 1 0 31472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_271
timestamp 1698431365
transform 1 0 31696 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_307
timestamp 1698431365
transform 1 0 35728 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_311
timestamp 1698431365
transform 1 0 36176 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_18
timestamp 1698431365
transform 1 0 3360 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_21
timestamp 1698431365
transform 1 0 3696 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_49
timestamp 1698431365
transform 1 0 6832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_58
timestamp 1698431365
transform 1 0 7840 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_78
timestamp 1698431365
transform 1 0 10080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_82
timestamp 1698431365
transform 1 0 10528 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_98
timestamp 1698431365
transform 1 0 12320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_102
timestamp 1698431365
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_113
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_126
timestamp 1698431365
transform 1 0 15456 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_130
timestamp 1698431365
transform 1 0 15904 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_146
timestamp 1698431365
transform 1 0 17696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_163
timestamp 1698431365
transform 1 0 19600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_167
timestamp 1698431365
transform 1 0 20048 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_199
timestamp 1698431365
transform 1 0 23632 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_218
timestamp 1698431365
transform 1 0 25760 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_233
timestamp 1698431365
transform 1 0 27440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_251
timestamp 1698431365
transform 1 0 29456 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_253
timestamp 1698431365
transform 1 0 29680 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_267
timestamp 1698431365
transform 1 0 31248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_310
timestamp 1698431365
transform 1 0 36064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_335
timestamp 1698431365
transform 1 0 38864 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_34
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_50
timestamp 1698431365
transform 1 0 6944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_58
timestamp 1698431365
transform 1 0 7840 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_90
timestamp 1698431365
transform 1 0 11424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_94
timestamp 1698431365
transform 1 0 11872 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_126
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_134
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_154
timestamp 1698431365
transform 1 0 18592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_158
timestamp 1698431365
transform 1 0 19040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_162
timestamp 1698431365
transform 1 0 19488 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_178
timestamp 1698431365
transform 1 0 21280 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_186
timestamp 1698431365
transform 1 0 22176 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_190
timestamp 1698431365
transform 1 0 22624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_218
timestamp 1698431365
transform 1 0 25760 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_222
timestamp 1698431365
transform 1 0 26208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_224
timestamp 1698431365
transform 1 0 26432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_258
timestamp 1698431365
transform 1 0 30240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_262
timestamp 1698431365
transform 1 0 30688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_307
timestamp 1698431365
transform 1 0 35728 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_311
timestamp 1698431365
transform 1 0 36176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_313
timestamp 1698431365
transform 1 0 36400 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_322
timestamp 1698431365
transform 1 0 37408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_338
timestamp 1698431365
transform 1 0 39200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_342
timestamp 1698431365
transform 1 0 39648 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_43
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_59
timestamp 1698431365
transform 1 0 7952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_61
timestamp 1698431365
transform 1 0 8176 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_67
timestamp 1698431365
transform 1 0 8848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_99
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_123
timestamp 1698431365
transform 1 0 15120 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_127
timestamp 1698431365
transform 1 0 15568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698431365
transform 1 0 20384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_187
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_210
timestamp 1698431365
transform 1 0 24864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_214
timestamp 1698431365
transform 1 0 25312 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_230
timestamp 1698431365
transform 1 0 27104 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_238
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_263
timestamp 1698431365
transform 1 0 30800 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_267
timestamp 1698431365
transform 1 0 31248 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_269
timestamp 1698431365
transform 1 0 31472 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_272
timestamp 1698431365
transform 1 0 31808 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_276
timestamp 1698431365
transform 1 0 32256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_302
timestamp 1698431365
transform 1 0 35168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_310
timestamp 1698431365
transform 1 0 36064 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_329
timestamp 1698431365
transform 1 0 38192 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_337
timestamp 1698431365
transform 1 0 39088 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_341
timestamp 1698431365
transform 1 0 39536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_22
timestamp 1698431365
transform 1 0 3808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_30
timestamp 1698431365
transform 1 0 4704 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_62
timestamp 1698431365
transform 1 0 8288 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_104
timestamp 1698431365
transform 1 0 12992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_106
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_121
timestamp 1698431365
transform 1 0 14896 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698431365
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_148
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_154
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_158
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_167
timestamp 1698431365
transform 1 0 20048 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_199
timestamp 1698431365
transform 1 0 23632 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_226
timestamp 1698431365
transform 1 0 26656 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_258
timestamp 1698431365
transform 1 0 30240 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_266
timestamp 1698431365
transform 1 0 31136 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698431365
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_293
timestamp 1698431365
transform 1 0 34160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_297
timestamp 1698431365
transform 1 0 34608 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_301
timestamp 1698431365
transform 1 0 35056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_303
timestamp 1698431365
transform 1 0 35280 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_333
timestamp 1698431365
transform 1 0 38640 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_341
timestamp 1698431365
transform 1 0 39536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_28
timestamp 1698431365
transform 1 0 4480 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_45
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_61
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_65
timestamp 1698431365
transform 1 0 8624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_67
timestamp 1698431365
transform 1 0 8848 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_128
timestamp 1698431365
transform 1 0 15680 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_132
timestamp 1698431365
transform 1 0 16128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_136
timestamp 1698431365
transform 1 0 16576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_138
timestamp 1698431365
transform 1 0 16800 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_145
timestamp 1698431365
transform 1 0 17584 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_153
timestamp 1698431365
transform 1 0 18480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_157
timestamp 1698431365
transform 1 0 18928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_165
timestamp 1698431365
transform 1 0 19824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_187
timestamp 1698431365
transform 1 0 22288 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_191
timestamp 1698431365
transform 1 0 22736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_193
timestamp 1698431365
transform 1 0 22960 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_200
timestamp 1698431365
transform 1 0 23744 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_216
timestamp 1698431365
transform 1 0 25536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_220
timestamp 1698431365
transform 1 0 25984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_222
timestamp 1698431365
transform 1 0 26208 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_233
timestamp 1698431365
transform 1 0 27440 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_237
timestamp 1698431365
transform 1 0 27888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_263
timestamp 1698431365
transform 1 0 30800 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_291
timestamp 1698431365
transform 1 0 33936 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_307
timestamp 1698431365
transform 1 0 35728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_309
timestamp 1698431365
transform 1 0 35952 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_341
timestamp 1698431365
transform 1 0 39536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_10
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_18
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_28
timestamp 1698431365
transform 1 0 4480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_36
timestamp 1698431365
transform 1 0 5376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_38
timestamp 1698431365
transform 1 0 5600 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_49
timestamp 1698431365
transform 1 0 6832 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_57
timestamp 1698431365
transform 1 0 7728 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_86
timestamp 1698431365
transform 1 0 10976 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_94
timestamp 1698431365
transform 1 0 11872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_96
timestamp 1698431365
transform 1 0 12096 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_154
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_173
timestamp 1698431365
transform 1 0 20720 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_241
timestamp 1698431365
transform 1 0 28336 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_245
timestamp 1698431365
transform 1 0 28784 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_298
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_302
timestamp 1698431365
transform 1 0 35168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_304
timestamp 1698431365
transform 1 0 35392 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_311
timestamp 1698431365
transform 1 0 36176 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_45
timestamp 1698431365
transform 1 0 6384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_49
timestamp 1698431365
transform 1 0 6832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_83
timestamp 1698431365
transform 1 0 10640 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_94
timestamp 1698431365
transform 1 0 11872 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_102
timestamp 1698431365
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_115
timestamp 1698431365
transform 1 0 14224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_117
timestamp 1698431365
transform 1 0 14448 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_124
timestamp 1698431365
transform 1 0 15232 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_158
timestamp 1698431365
transform 1 0 19040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_170
timestamp 1698431365
transform 1 0 20384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_183
timestamp 1698431365
transform 1 0 21840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_187
timestamp 1698431365
transform 1 0 22288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_189
timestamp 1698431365
transform 1 0 22512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_225
timestamp 1698431365
transform 1 0 26544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_229
timestamp 1698431365
transform 1 0 26992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_238
timestamp 1698431365
transform 1 0 28000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_255
timestamp 1698431365
transform 1 0 29904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_259
timestamp 1698431365
transform 1 0 30352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_262
timestamp 1698431365
transform 1 0 30688 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_278
timestamp 1698431365
transform 1 0 32480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_282
timestamp 1698431365
transform 1 0 32928 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_291
timestamp 1698431365
transform 1 0 33936 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_307
timestamp 1698431365
transform 1 0 35728 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_327
timestamp 1698431365
transform 1 0 37968 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_10
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_26
timestamp 1698431365
transform 1 0 4256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_30
timestamp 1698431365
transform 1 0 4704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_38
timestamp 1698431365
transform 1 0 5600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_42
timestamp 1698431365
transform 1 0 6048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_78
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_94
timestamp 1698431365
transform 1 0 11872 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_102
timestamp 1698431365
transform 1 0 12768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_125
timestamp 1698431365
transform 1 0 15344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_129
timestamp 1698431365
transform 1 0 15792 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698431365
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_221
timestamp 1698431365
transform 1 0 26096 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_257
timestamp 1698431365
transform 1 0 30128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_261
timestamp 1698431365
transform 1 0 30576 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698431365
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_298
timestamp 1698431365
transform 1 0 34720 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_306
timestamp 1698431365
transform 1 0 35616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_310
timestamp 1698431365
transform 1 0 36064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698431365
transform 1 0 9072 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_73
timestamp 1698431365
transform 1 0 9520 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_85
timestamp 1698431365
transform 1 0 10864 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_120
timestamp 1698431365
transform 1 0 14784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_122
timestamp 1698431365
transform 1 0 15008 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_133
timestamp 1698431365
transform 1 0 16240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_137
timestamp 1698431365
transform 1 0 16688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_141
timestamp 1698431365
transform 1 0 17136 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_145
timestamp 1698431365
transform 1 0 17584 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_209
timestamp 1698431365
transform 1 0 24752 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_225
timestamp 1698431365
transform 1 0 26544 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_233
timestamp 1698431365
transform 1 0 27440 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698431365
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_262
timestamp 1698431365
transform 1 0 30688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_266
timestamp 1698431365
transform 1 0 31136 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_337
timestamp 1698431365
transform 1 0 39088 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_341
timestamp 1698431365
transform 1 0 39536 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_10
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_14
timestamp 1698431365
transform 1 0 2912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_21
timestamp 1698431365
transform 1 0 3696 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_37
timestamp 1698431365
transform 1 0 5488 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_45
timestamp 1698431365
transform 1 0 6384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_47
timestamp 1698431365
transform 1 0 6608 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_54
timestamp 1698431365
transform 1 0 7392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_56
timestamp 1698431365
transform 1 0 7616 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_65
timestamp 1698431365
transform 1 0 8624 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698431365
transform 1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_96
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_134
timestamp 1698431365
transform 1 0 16352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_168
timestamp 1698431365
transform 1 0 20160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_172
timestamp 1698431365
transform 1 0 20608 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_180
timestamp 1698431365
transform 1 0 21504 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_184
timestamp 1698431365
transform 1 0 21952 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_195
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_199
timestamp 1698431365
transform 1 0 23632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_224
timestamp 1698431365
transform 1 0 26432 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_226
timestamp 1698431365
transform 1 0 26656 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_237
timestamp 1698431365
transform 1 0 27888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_245
timestamp 1698431365
transform 1 0 28784 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_253
timestamp 1698431365
transform 1 0 29680 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_257
timestamp 1698431365
transform 1 0 30128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_261
timestamp 1698431365
transform 1 0 30576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_307
timestamp 1698431365
transform 1 0 35728 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_315
timestamp 1698431365
transform 1 0 36624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_317
timestamp 1698431365
transform 1 0 36848 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_339
timestamp 1698431365
transform 1 0 39312 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_18
timestamp 1698431365
transform 1 0 3360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_33
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_51
timestamp 1698431365
transform 1 0 7056 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_92
timestamp 1698431365
transform 1 0 11648 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_96
timestamp 1698431365
transform 1 0 12096 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_100
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_116
timestamp 1698431365
transform 1 0 14336 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_126
timestamp 1698431365
transform 1 0 15456 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_159
timestamp 1698431365
transform 1 0 19152 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_163
timestamp 1698431365
transform 1 0 19600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_179
timestamp 1698431365
transform 1 0 21392 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_209
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_213
timestamp 1698431365
transform 1 0 25200 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_221
timestamp 1698431365
transform 1 0 26096 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_223
timestamp 1698431365
transform 1 0 26320 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_229
timestamp 1698431365
transform 1 0 26992 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_263
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_267
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_270
timestamp 1698431365
transform 1 0 31584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_272
timestamp 1698431365
transform 1 0 31808 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_304
timestamp 1698431365
transform 1 0 35392 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_308
timestamp 1698431365
transform 1 0 35840 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_326
timestamp 1698431365
transform 1 0 37856 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_342
timestamp 1698431365
transform 1 0 39648 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_43
timestamp 1698431365
transform 1 0 6160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_51
timestamp 1698431365
transform 1 0 7056 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_67
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_158
timestamp 1698431365
transform 1 0 19040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_162
timestamp 1698431365
transform 1 0 19488 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_178
timestamp 1698431365
transform 1 0 21280 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_182
timestamp 1698431365
transform 1 0 21728 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_198
timestamp 1698431365
transform 1 0 23520 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_224
timestamp 1698431365
transform 1 0 26432 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_258
timestamp 1698431365
transform 1 0 30240 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_298
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_326
timestamp 1698431365
transform 1 0 37856 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_342
timestamp 1698431365
transform 1 0 39648 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_10
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_14
timestamp 1698431365
transform 1 0 2912 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_21
timestamp 1698431365
transform 1 0 3696 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_29
timestamp 1698431365
transform 1 0 4592 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_33
timestamp 1698431365
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_64
timestamp 1698431365
transform 1 0 8512 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_96
timestamp 1698431365
transform 1 0 12096 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_136
timestamp 1698431365
transform 1 0 16576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_140
timestamp 1698431365
transform 1 0 17024 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_189
timestamp 1698431365
transform 1 0 22512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_192
timestamp 1698431365
transform 1 0 22848 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_208
timestamp 1698431365
transform 1 0 24640 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_224
timestamp 1698431365
transform 1 0 26432 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698431365
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_261
timestamp 1698431365
transform 1 0 30576 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_293
timestamp 1698431365
transform 1 0 34160 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_333
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_341
timestamp 1698431365
transform 1 0 39536 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_34
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_42
timestamp 1698431365
transform 1 0 6048 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_49
timestamp 1698431365
transform 1 0 6832 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_65
timestamp 1698431365
transform 1 0 8624 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_88
timestamp 1698431365
transform 1 0 11200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_162
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_164
timestamp 1698431365
transform 1 0 19712 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_194
timestamp 1698431365
transform 1 0 23072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_198
timestamp 1698431365
transform 1 0 23520 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_250
timestamp 1698431365
transform 1 0 29344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_254
timestamp 1698431365
transform 1 0 29792 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_258
timestamp 1698431365
transform 1 0 30240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_260
timestamp 1698431365
transform 1 0 30464 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_290
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_294
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_296
timestamp 1698431365
transform 1 0 34496 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_305
timestamp 1698431365
transform 1 0 35504 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_307
timestamp 1698431365
transform 1 0 35728 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_31
timestamp 1698431365
transform 1 0 4816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_49
timestamp 1698431365
transform 1 0 6832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_51
timestamp 1698431365
transform 1 0 7056 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_54
timestamp 1698431365
transform 1 0 7392 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_62
timestamp 1698431365
transform 1 0 8288 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_78
timestamp 1698431365
transform 1 0 10080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_82
timestamp 1698431365
transform 1 0 10528 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_98
timestamp 1698431365
transform 1 0 12320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_102
timestamp 1698431365
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_113
timestamp 1698431365
transform 1 0 14000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_117
timestamp 1698431365
transform 1 0 14448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_125
timestamp 1698431365
transform 1 0 15344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_158
timestamp 1698431365
transform 1 0 19040 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_209
timestamp 1698431365
transform 1 0 24752 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_235
timestamp 1698431365
transform 1 0 27664 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_259
timestamp 1698431365
transform 1 0 30352 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_267
timestamp 1698431365
transform 1 0 31248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_300
timestamp 1698431365
transform 1 0 34944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_304
timestamp 1698431365
transform 1 0 35392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_341
timestamp 1698431365
transform 1 0 39536 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_20
timestamp 1698431365
transform 1 0 3584 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_52
timestamp 1698431365
transform 1 0 7168 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_76
timestamp 1698431365
transform 1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_78
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_90
timestamp 1698431365
transform 1 0 11424 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_122
timestamp 1698431365
transform 1 0 15008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_124
timestamp 1698431365
transform 1 0 15232 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_127
timestamp 1698431365
transform 1 0 15568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_135
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_174
timestamp 1698431365
transform 1 0 20832 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_178
timestamp 1698431365
transform 1 0 21280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_188
timestamp 1698431365
transform 1 0 22400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_192
timestamp 1698431365
transform 1 0 22848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_196
timestamp 1698431365
transform 1 0 23296 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698431365
transform 1 0 24192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_223
timestamp 1698431365
transform 1 0 26320 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_227
timestamp 1698431365
transform 1 0 26768 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_290
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_298
timestamp 1698431365
transform 1 0 34720 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_302
timestamp 1698431365
transform 1 0 35168 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_306
timestamp 1698431365
transform 1 0 35616 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_314
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_318
timestamp 1698431365
transform 1 0 36960 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_331
timestamp 1698431365
transform 1 0 38416 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_339
timestamp 1698431365
transform 1 0 39312 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_53
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_57
timestamp 1698431365
transform 1 0 7728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_77
timestamp 1698431365
transform 1 0 9968 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_88
timestamp 1698431365
transform 1 0 11200 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_100
timestamp 1698431365
transform 1 0 12544 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_118
timestamp 1698431365
transform 1 0 14560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_122
timestamp 1698431365
transform 1 0 15008 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_154
timestamp 1698431365
transform 1 0 18592 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_162
timestamp 1698431365
transform 1 0 19488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_166
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_189
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_206
timestamp 1698431365
transform 1 0 24416 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_222
timestamp 1698431365
transform 1 0 26208 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_226
timestamp 1698431365
transform 1 0 26656 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_234
timestamp 1698431365
transform 1 0 27552 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_251
timestamp 1698431365
transform 1 0 29456 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_257
timestamp 1698431365
transform 1 0 30128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_283
timestamp 1698431365
transform 1 0 33040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_287
timestamp 1698431365
transform 1 0 33488 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_303
timestamp 1698431365
transform 1 0 35280 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_333
timestamp 1698431365
transform 1 0 38640 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_341
timestamp 1698431365
transform 1 0 39536 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_32
timestamp 1698431365
transform 1 0 4928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_36
timestamp 1698431365
transform 1 0 5376 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_76
timestamp 1698431365
transform 1 0 9856 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_93
timestamp 1698431365
transform 1 0 11760 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_109
timestamp 1698431365
transform 1 0 13552 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_120
timestamp 1698431365
transform 1 0 14784 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_148
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_152
timestamp 1698431365
transform 1 0 18368 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_156
timestamp 1698431365
transform 1 0 18816 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_162
timestamp 1698431365
transform 1 0 19488 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_199
timestamp 1698431365
transform 1 0 23632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_203
timestamp 1698431365
transform 1 0 24080 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_207
timestamp 1698431365
transform 1 0 24528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_218
timestamp 1698431365
transform 1 0 25760 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_245
timestamp 1698431365
transform 1 0 28784 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_271
timestamp 1698431365
transform 1 0 31696 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_314
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_329
timestamp 1698431365
transform 1 0 38192 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_337
timestamp 1698431365
transform 1 0 39088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_341
timestamp 1698431365
transform 1 0 39536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_43
timestamp 1698431365
transform 1 0 6160 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_50
timestamp 1698431365
transform 1 0 6944 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_54
timestamp 1698431365
transform 1 0 7392 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_68
timestamp 1698431365
transform 1 0 8960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_76
timestamp 1698431365
transform 1 0 9856 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_78
timestamp 1698431365
transform 1 0 10080 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_86
timestamp 1698431365
transform 1 0 10976 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_97
timestamp 1698431365
transform 1 0 12208 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_122
timestamp 1698431365
transform 1 0 15008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_130
timestamp 1698431365
transform 1 0 15904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_134
timestamp 1698431365
transform 1 0 16352 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_136
timestamp 1698431365
transform 1 0 16576 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_147
timestamp 1698431365
transform 1 0 17808 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_157
timestamp 1698431365
transform 1 0 18928 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_173
timestamp 1698431365
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_193
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_197
timestamp 1698431365
transform 1 0 23408 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_208
timestamp 1698431365
transform 1 0 24640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_212
timestamp 1698431365
transform 1 0 25088 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_216
timestamp 1698431365
transform 1 0 25536 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_239
timestamp 1698431365
transform 1 0 28112 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_243
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_251
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_259
timestamp 1698431365
transform 1 0 30352 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_280
timestamp 1698431365
transform 1 0 32704 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_296
timestamp 1698431365
transform 1 0 34496 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_304
timestamp 1698431365
transform 1 0 35392 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_306
timestamp 1698431365
transform 1 0 35616 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_341
timestamp 1698431365
transform 1 0 39536 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_10
timestamp 1698431365
transform 1 0 2464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_54
timestamp 1698431365
transform 1 0 7392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_56
timestamp 1698431365
transform 1 0 7616 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_83
timestamp 1698431365
transform 1 0 10640 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_99
timestamp 1698431365
transform 1 0 12432 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_107
timestamp 1698431365
transform 1 0 13328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_115
timestamp 1698431365
transform 1 0 14224 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_123
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_127
timestamp 1698431365
transform 1 0 15568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_129
timestamp 1698431365
transform 1 0 15792 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_158
timestamp 1698431365
transform 1 0 19040 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_174
timestamp 1698431365
transform 1 0 20832 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_182
timestamp 1698431365
transform 1 0 21728 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_186
timestamp 1698431365
transform 1 0 22176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_188
timestamp 1698431365
transform 1 0 22400 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_205
timestamp 1698431365
transform 1 0 24304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_244
timestamp 1698431365
transform 1 0 28672 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_248
timestamp 1698431365
transform 1 0 29120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_250
timestamp 1698431365
transform 1 0 29344 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_261
timestamp 1698431365
transform 1 0 30576 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_269
timestamp 1698431365
transform 1 0 31472 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_289
timestamp 1698431365
transform 1 0 33712 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_327
timestamp 1698431365
transform 1 0 37968 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_53
timestamp 1698431365
transform 1 0 7280 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_57
timestamp 1698431365
transform 1 0 7728 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_59
timestamp 1698431365
transform 1 0 7952 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_85
timestamp 1698431365
transform 1 0 10864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_98
timestamp 1698431365
transform 1 0 12320 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_151
timestamp 1698431365
transform 1 0 18256 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_155
timestamp 1698431365
transform 1 0 18704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_159
timestamp 1698431365
transform 1 0 19152 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_167
timestamp 1698431365
transform 1 0 20048 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_187
timestamp 1698431365
transform 1 0 22288 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_219
timestamp 1698431365
transform 1 0 25872 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_235
timestamp 1698431365
transform 1 0 27664 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_275
timestamp 1698431365
transform 1 0 32144 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_291
timestamp 1698431365
transform 1 0 33936 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_293
timestamp 1698431365
transform 1 0 34160 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_309
timestamp 1698431365
transform 1 0 35952 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_323
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_339
timestamp 1698431365
transform 1 0 39312 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_76
timestamp 1698431365
transform 1 0 9856 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_128
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_132
timestamp 1698431365
transform 1 0 16128 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_152
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_156
timestamp 1698431365
transform 1 0 18816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_158
timestamp 1698431365
transform 1 0 19040 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_196
timestamp 1698431365
transform 1 0 23296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_200
timestamp 1698431365
transform 1 0 23744 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_208
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_218
timestamp 1698431365
transform 1 0 25760 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_249
timestamp 1698431365
transform 1 0 29232 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_287
timestamp 1698431365
transform 1 0 33488 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_291
timestamp 1698431365
transform 1 0 33936 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_309
timestamp 1698431365
transform 1 0 35952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_311
timestamp 1698431365
transform 1 0 36176 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_49
timestamp 1698431365
transform 1 0 6832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_63
timestamp 1698431365
transform 1 0 8400 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_67
timestamp 1698431365
transform 1 0 8848 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_92
timestamp 1698431365
transform 1 0 11648 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_96
timestamp 1698431365
transform 1 0 12096 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_98
timestamp 1698431365
transform 1 0 12320 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_134
timestamp 1698431365
transform 1 0 16352 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_146
timestamp 1698431365
transform 1 0 17696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_201
timestamp 1698431365
transform 1 0 23856 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_209
timestamp 1698431365
transform 1 0 24752 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_228
timestamp 1698431365
transform 1 0 26880 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_236
timestamp 1698431365
transform 1 0 27776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_309
timestamp 1698431365
transform 1 0 35952 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_333
timestamp 1698431365
transform 1 0 38640 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_341
timestamp 1698431365
transform 1 0 39536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_84
timestamp 1698431365
transform 1 0 10752 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_92
timestamp 1698431365
transform 1 0 11648 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_96
timestamp 1698431365
transform 1 0 12096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_116
timestamp 1698431365
transform 1 0 14336 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_135
timestamp 1698431365
transform 1 0 16464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_149
timestamp 1698431365
transform 1 0 18032 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_167
timestamp 1698431365
transform 1 0 20048 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_177
timestamp 1698431365
transform 1 0 21168 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698431365
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_241
timestamp 1698431365
transform 1 0 28336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_243
timestamp 1698431365
transform 1 0 28560 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_277
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_290
timestamp 1698431365
transform 1 0 33824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_323
timestamp 1698431365
transform 1 0 37520 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_339
timestamp 1698431365
transform 1 0 39312 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_72
timestamp 1698431365
transform 1 0 9408 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_76
timestamp 1698431365
transform 1 0 9856 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_84
timestamp 1698431365
transform 1 0 10752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_86
timestamp 1698431365
transform 1 0 10976 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_123
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_131
timestamp 1698431365
transform 1 0 16016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_135
timestamp 1698431365
transform 1 0 16464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_137
timestamp 1698431365
transform 1 0 16688 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_155
timestamp 1698431365
transform 1 0 18704 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_189
timestamp 1698431365
transform 1 0 22512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_198
timestamp 1698431365
transform 1 0 23520 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_230
timestamp 1698431365
transform 1 0 27104 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_238
timestamp 1698431365
transform 1 0 28000 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_240
timestamp 1698431365
transform 1 0 28224 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_283
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_309
timestamp 1698431365
transform 1 0 35952 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_333
timestamp 1698431365
transform 1 0 38640 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_341
timestamp 1698431365
transform 1 0 39536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_34
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_38
timestamp 1698431365
transform 1 0 5600 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_40
timestamp 1698431365
transform 1 0 5824 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_76
timestamp 1698431365
transform 1 0 9856 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_92
timestamp 1698431365
transform 1 0 11648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_121
timestamp 1698431365
transform 1 0 14896 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_137
timestamp 1698431365
transform 1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_158
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_160
timestamp 1698431365
transform 1 0 19264 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_167
timestamp 1698431365
transform 1 0 20048 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_175
timestamp 1698431365
transform 1 0 20944 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_179
timestamp 1698431365
transform 1 0 21392 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_193
timestamp 1698431365
transform 1 0 22960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_197
timestamp 1698431365
transform 1 0 23408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_201
timestamp 1698431365
transform 1 0 23856 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_228
timestamp 1698431365
transform 1 0 26880 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_236
timestamp 1698431365
transform 1 0 27776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_267
timestamp 1698431365
transform 1 0 31248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_271
timestamp 1698431365
transform 1 0 31696 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_314
timestamp 1698431365
transform 1 0 36512 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_330
timestamp 1698431365
transform 1 0 38304 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_338
timestamp 1698431365
transform 1 0 39200 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_342
timestamp 1698431365
transform 1 0 39648 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_69
timestamp 1698431365
transform 1 0 9072 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_85
timestamp 1698431365
transform 1 0 10864 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_93
timestamp 1698431365
transform 1 0 11760 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_97
timestamp 1698431365
transform 1 0 12208 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_99
timestamp 1698431365
transform 1 0 12432 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_102
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_115
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_131
timestamp 1698431365
transform 1 0 16016 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_139
timestamp 1698431365
transform 1 0 16912 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_143
timestamp 1698431365
transform 1 0 17360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_145
timestamp 1698431365
transform 1 0 17584 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_148
timestamp 1698431365
transform 1 0 17920 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_164
timestamp 1698431365
transform 1 0 19712 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_220
timestamp 1698431365
transform 1 0 25984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_224
timestamp 1698431365
transform 1 0 26432 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_279
timestamp 1698431365
transform 1 0 32592 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_291
timestamp 1698431365
transform 1 0 33936 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_307
timestamp 1698431365
transform 1 0 35728 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698431365
transform 1 0 38640 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_341
timestamp 1698431365
transform 1 0 39536 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_104
timestamp 1698431365
transform 1 0 12992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_114
timestamp 1698431365
transform 1 0 14112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_118
timestamp 1698431365
transform 1 0 14560 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_156
timestamp 1698431365
transform 1 0 18816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_160
timestamp 1698431365
transform 1 0 19264 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_168
timestamp 1698431365
transform 1 0 20160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_172
timestamp 1698431365
transform 1 0 20608 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_180
timestamp 1698431365
transform 1 0 21504 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_184
timestamp 1698431365
transform 1 0 21952 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_188
timestamp 1698431365
transform 1 0 22400 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_196
timestamp 1698431365
transform 1 0 23296 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_199
timestamp 1698431365
transform 1 0 23632 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_203
timestamp 1698431365
transform 1 0 24080 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_243
timestamp 1698431365
transform 1 0 28560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_247
timestamp 1698431365
transform 1 0 29008 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_314
timestamp 1698431365
transform 1 0 36512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_330
timestamp 1698431365
transform 1 0 38304 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_338
timestamp 1698431365
transform 1 0 39200 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_342
timestamp 1698431365
transform 1 0 39648 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_69
timestamp 1698431365
transform 1 0 9072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_71
timestamp 1698431365
transform 1 0 9296 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_80
timestamp 1698431365
transform 1 0 10304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_84
timestamp 1698431365
transform 1 0 10752 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_86
timestamp 1698431365
transform 1 0 10976 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_93
timestamp 1698431365
transform 1 0 11760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_95
timestamp 1698431365
transform 1 0 11984 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_116
timestamp 1698431365
transform 1 0 14336 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_124
timestamp 1698431365
transform 1 0 15232 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_128
timestamp 1698431365
transform 1 0 15680 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_138
timestamp 1698431365
transform 1 0 16800 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698431365
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_192
timestamp 1698431365
transform 1 0 22848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_196
timestamp 1698431365
transform 1 0 23296 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_228
timestamp 1698431365
transform 1 0 26880 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_341
timestamp 1698431365
transform 1 0 39536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_88
timestamp 1698431365
transform 1 0 11200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_90
timestamp 1698431365
transform 1 0 11424 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_111
timestamp 1698431365
transform 1 0 13776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_115
timestamp 1698431365
transform 1 0 14224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_156
timestamp 1698431365
transform 1 0 18816 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_160
timestamp 1698431365
transform 1 0 19264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_194
timestamp 1698431365
transform 1 0 23072 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_314
timestamp 1698431365
transform 1 0 36512 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_330
timestamp 1698431365
transform 1 0 38304 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_338
timestamp 1698431365
transform 1 0 39200 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_342
timestamp 1698431365
transform 1 0 39648 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_69
timestamp 1698431365
transform 1 0 9072 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_73
timestamp 1698431365
transform 1 0 9520 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_75
timestamp 1698431365
transform 1 0 9744 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_119
timestamp 1698431365
transform 1 0 14672 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_123
timestamp 1698431365
transform 1 0 15120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_156
timestamp 1698431365
transform 1 0 18816 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_172
timestamp 1698431365
transform 1 0 20608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_206
timestamp 1698431365
transform 1 0 24416 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_210
timestamp 1698431365
transform 1 0 24864 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_333
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_341
timestamp 1698431365
transform 1 0 39536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_314
timestamp 1698431365
transform 1 0 36512 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_330
timestamp 1698431365
transform 1 0 38304 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_338
timestamp 1698431365
transform 1 0 39200 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_342
timestamp 1698431365
transform 1 0 39648 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_36
timestamp 1698431365
transform 1 0 5376 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_70
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_138
timestamp 1698431365
transform 1 0 16800 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_206
timestamp 1698431365
transform 1 0 24416 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_240
timestamp 1698431365
transform 1 0 28224 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_274
timestamp 1698431365
transform 1 0 32032 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_308
timestamp 1698431365
transform 1 0 35840 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_342
timestamp 1698431365
transform 1 0 39648 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39760 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36288 0 1 9408
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  hold3
timestamp 1698431365
transform -1 0 28448 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 24416 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 39760 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform -1 0 35728 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform 1 0 34720 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform -1 0 37968 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  hold10
timestamp 1698431365
transform -1 0 36064 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 36176 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold13
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold14
timestamp 1698431365
transform -1 0 36512 0 -1 14112
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold15
timestamp 1698431365
transform -1 0 35728 0 -1 15680
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold16
timestamp 1698431365
transform -1 0 35728 0 -1 17248
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold17
timestamp 1698431365
transform 1 0 32368 0 1 17248
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold18
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold19
timestamp 1698431365
transform 1 0 36960 0 1 14112
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold20
timestamp 1698431365
transform -1 0 38976 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold21
timestamp 1698431365
transform 1 0 32816 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 6048 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 38192 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 38864 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 32816 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 31136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 32032 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 3248 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698431365
transform -1 0 9184 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698431365
transform 1 0 5936 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698431365
transform 1 0 13664 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform -1 0 15568 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform -1 0 12656 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_49 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 39984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 39984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 39984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 39984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 39984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 39984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 39984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 39984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 39984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 39984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 39984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 39984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 39984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 39984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 39984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 39984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 39984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 39984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 39984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 39984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 39984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 39984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 39984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 39984 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 39984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 39984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 39984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 39984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 39984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 39984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 39984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 39984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 39984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 39984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 39984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 39984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 39984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 39984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 39984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 39984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 39984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 39984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 39984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 39984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 39984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 39984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 39984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 39984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 39984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_108
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_109
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_110
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_112
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_113
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_114
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_115
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_117
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_118
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_119
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_120
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_121
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_122
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_123
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_124
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_125
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_126
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_127
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_128
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_129
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_130
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_131
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_132
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_133
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_134
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_135
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_136
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_137
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_138
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_139
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_140
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_141
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_142
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_143
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_144
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_145
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_146
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_147
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_148
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_149
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_150
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_151
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_152
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_153
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_154
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_155
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_156
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_157
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_158
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_159
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_160
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_161
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_162
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_163
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_164
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_165
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_166
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_167
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_168
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_169
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_170
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_171
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_172
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_173
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_174
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_175
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_176
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_177
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_178
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_179
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_180
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_181
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_182
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_183
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_184
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_185
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_186
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_187
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_188
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_189
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_190
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_191
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_192
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_193
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_194
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_195
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_196
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_197
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_198
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_199
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_200
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_201
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_202
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_203
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_204
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_205
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_206
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_207
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_208
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_209
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_210
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_211
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_212
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_213
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_214
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_215
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_216
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_217
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_218
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_219
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_220
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_221
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_222
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_223
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_224
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_225
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_226
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_227
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_228
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_229
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_230
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_231
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_232
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_233
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_234
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_235
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_236
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_237
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_238
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_239
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_240
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_241
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_242
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_243
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_244
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_245
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_246
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_247
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_248
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_249
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_250
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_251
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_252
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_253
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_254
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_255
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_256
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_257
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_258
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_259
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_260
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_261
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_262
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_263
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_264
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_265
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_266
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_267
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_268
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_269
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_270
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_271
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_272
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_273
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_274
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_275
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_276
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_277
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_278
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_279
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_280
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_281
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_282
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_283
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_284
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_285
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_286
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_287
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_288
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_289
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_290
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_291
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_292
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_293
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_294
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_295
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_296
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_297
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_298
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_299
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_300
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_303
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_304
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_305
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_306
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_307
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_308
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_309
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_310
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_311
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_312
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_313
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_314
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_315
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_316
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_317
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_318
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_319
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_320
timestamp 1698431365
transform 1 0 8960 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_321
timestamp 1698431365
transform 1 0 12768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_322
timestamp 1698431365
transform 1 0 16576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_323
timestamp 1698431365
transform 1 0 20384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_324
timestamp 1698431365
transform 1 0 24192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_325
timestamp 1698431365
transform 1 0 28000 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_326
timestamp 1698431365
transform 1 0 31808 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_327
timestamp 1698431365
transform 1 0 35616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_328
timestamp 1698431365
transform 1 0 39424 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_solo_squash_16 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_solo_squash_17
timestamp 1698431365
transform -1 0 21168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_solo_squash_18
timestamp 1698431365
transform -1 0 20160 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_solo_squash_19
timestamp 1698431365
transform -1 0 18480 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_solo_squash_20
timestamp 1698431365
transform -1 0 17696 0 -1 4704
box -86 -86 534 870
<< labels >>
flabel metal2 s 1792 0 1904 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 4480 0 4592 800 0 FreeSans 448 90 0 0 gpio_ready
port 1 nsew signal input
flabel metal2 s 39424 0 39536 800 0 FreeSans 448 90 0 0 io_in[0]
port 2 nsew signal input
flabel metal2 s 25984 0 26096 800 0 FreeSans 448 90 0 0 io_in[10]
port 3 nsew signal input
flabel metal2 s 24640 0 24752 800 0 FreeSans 448 90 0 0 io_in[11]
port 4 nsew signal input
flabel metal2 s 23296 0 23408 800 0 FreeSans 448 90 0 0 io_in[12]
port 5 nsew signal input
flabel metal2 s 38080 0 38192 800 0 FreeSans 448 90 0 0 io_in[1]
port 6 nsew signal input
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 io_in[2]
port 7 nsew signal input
flabel metal2 s 35392 0 35504 800 0 FreeSans 448 90 0 0 io_in[3]
port 8 nsew signal input
flabel metal2 s 34048 0 34160 800 0 FreeSans 448 90 0 0 io_in[4]
port 9 nsew signal input
flabel metal2 s 32704 0 32816 800 0 FreeSans 448 90 0 0 io_in[5]
port 10 nsew signal input
flabel metal2 s 31360 0 31472 800 0 FreeSans 448 90 0 0 io_in[6]
port 11 nsew signal input
flabel metal2 s 30016 0 30128 800 0 FreeSans 448 90 0 0 io_in[7]
port 12 nsew signal input
flabel metal2 s 28672 0 28784 800 0 FreeSans 448 90 0 0 io_in[8]
port 13 nsew signal input
flabel metal2 s 27328 0 27440 800 0 FreeSans 448 90 0 0 io_in[9]
port 14 nsew signal input
flabel metal2 s 21952 0 22064 800 0 FreeSans 448 90 0 0 io_out[0]
port 15 nsew signal tristate
flabel metal2 s 8512 0 8624 800 0 FreeSans 448 90 0 0 io_out[10]
port 16 nsew signal tristate
flabel metal2 s 7168 0 7280 800 0 FreeSans 448 90 0 0 io_out[11]
port 17 nsew signal tristate
flabel metal2 s 5824 0 5936 800 0 FreeSans 448 90 0 0 io_out[12]
port 18 nsew signal tristate
flabel metal2 s 20608 0 20720 800 0 FreeSans 448 90 0 0 io_out[1]
port 19 nsew signal tristate
flabel metal2 s 19264 0 19376 800 0 FreeSans 448 90 0 0 io_out[2]
port 20 nsew signal tristate
flabel metal2 s 17920 0 18032 800 0 FreeSans 448 90 0 0 io_out[3]
port 21 nsew signal tristate
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 io_out[4]
port 22 nsew signal tristate
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 io_out[5]
port 23 nsew signal tristate
flabel metal2 s 13888 0 14000 800 0 FreeSans 448 90 0 0 io_out[6]
port 24 nsew signal tristate
flabel metal2 s 12544 0 12656 800 0 FreeSans 448 90 0 0 io_out[7]
port 25 nsew signal tristate
flabel metal2 s 11200 0 11312 800 0 FreeSans 448 90 0 0 io_out[8]
port 26 nsew signal tristate
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 io_out[9]
port 27 nsew signal tristate
flabel metal2 s 3136 0 3248 800 0 FreeSans 448 90 0 0 rst
port 28 nsew signal input
flabel metal4 s 4448 3076 4768 41612 0 FreeSans 1280 90 0 0 vdd
port 29 nsew power bidirectional
flabel metal4 s 35168 3076 35488 41612 0 FreeSans 1280 90 0 0 vdd
port 29 nsew power bidirectional
flabel metal4 s 19808 3076 20128 41612 0 FreeSans 1280 90 0 0 vss
port 30 nsew ground bidirectional
rlabel metal1 20664 41552 20664 41552 0 vdd
rlabel metal1 20664 40768 20664 40768 0 vss
rlabel metal2 21784 4480 21784 4480 0 _0000_
rlabel metal3 17136 5208 17136 5208 0 _0001_
rlabel metal2 10360 5264 10360 5264 0 _0002_
rlabel metal2 5992 4760 5992 4760 0 _0003_
rlabel metal3 8400 5208 8400 5208 0 _0004_
rlabel metal2 22344 10248 22344 10248 0 _0005_
rlabel metal2 31416 8960 31416 8960 0 _0006_
rlabel metal2 26152 4424 26152 4424 0 _0007_
rlabel metal2 24752 5208 24752 5208 0 _0008_
rlabel metal2 23576 6832 23576 6832 0 _0009_
rlabel metal2 33376 5208 33376 5208 0 _0010_
rlabel metal2 32032 16632 32032 16632 0 _0011_
rlabel metal2 38920 3920 38920 3920 0 _0012_
rlabel metal2 37744 14728 37744 14728 0 _0013_
rlabel metal2 31864 22680 31864 22680 0 _0014_
rlabel metal2 37576 21168 37576 21168 0 _0015_
rlabel metal2 38416 26824 38416 26824 0 _0016_
rlabel metal2 37408 31976 37408 31976 0 _0017_
rlabel metal2 36568 34608 36568 34608 0 _0018_
rlabel metal2 28952 34944 28952 34944 0 _0019_
rlabel metal2 33992 27776 33992 27776 0 _0020_
rlabel metal2 25592 33712 25592 33712 0 _0021_
rlabel metal2 21784 28280 21784 28280 0 _0022_
rlabel metal3 26096 37128 26096 37128 0 _0023_
rlabel metal2 23072 39480 23072 39480 0 _0024_
rlabel metal2 16632 39480 16632 39480 0 _0025_
rlabel metal2 6888 34496 6888 34496 0 _0026_
rlabel metal2 22344 32872 22344 32872 0 _0027_
rlabel metal2 12152 39256 12152 39256 0 _0028_
rlabel metal3 9240 35000 9240 35000 0 _0029_
rlabel metal3 16156 29960 16156 29960 0 _0030_
rlabel metal2 16856 23576 16856 23576 0 _0031_
rlabel metal3 14840 25592 14840 25592 0 _0032_
rlabel metal2 31528 23576 31528 23576 0 _0033_
rlabel metal2 16352 23352 16352 23352 0 _0034_
rlabel metal2 27832 21896 27832 21896 0 _0035_
rlabel metal2 2520 9184 2520 9184 0 _0036_
rlabel metal2 2688 7560 2688 7560 0 _0037_
rlabel metal2 3080 13328 3080 13328 0 _0038_
rlabel metal2 2744 14448 2744 14448 0 _0039_
rlabel metal2 2520 18424 2520 18424 0 _0040_
rlabel metal2 2520 20412 2520 20412 0 _0041_
rlabel metal2 8512 23240 8512 23240 0 _0042_
rlabel metal2 4760 23912 4760 23912 0 _0043_
rlabel metal2 2464 24920 2464 24920 0 _0044_
rlabel metal2 3192 26488 3192 26488 0 _0045_
rlabel metal2 14504 22736 14504 22736 0 _0046_
rlabel metal2 18648 7168 18648 7168 0 _0047_
rlabel metal2 18648 8680 18648 8680 0 _0048_
rlabel metal2 15848 11928 15848 11928 0 _0049_
rlabel metal2 14840 15456 14840 15456 0 _0050_
rlabel metal2 16968 17304 16968 17304 0 _0051_
rlabel metal2 18648 24360 18648 24360 0 _0052_
rlabel metal2 19656 21504 19656 21504 0 _0053_
rlabel metal2 23464 19992 23464 19992 0 _0054_
rlabel metal2 21560 21952 21560 21952 0 _0055_
rlabel metal2 27496 17192 27496 17192 0 _0056_
rlabel metal3 7280 4536 7280 4536 0 _0057_
rlabel metal2 15176 18648 15176 18648 0 _0058_
rlabel metal2 14504 19320 14504 19320 0 _0059_
rlabel metal2 15960 20048 15960 20048 0 _0060_
rlabel metal2 25144 19264 25144 19264 0 _0061_
rlabel metal2 19992 19880 19992 19880 0 _0062_
rlabel metal3 25592 19992 25592 19992 0 _0063_
rlabel metal2 26712 21112 26712 21112 0 _0064_
rlabel metal2 21560 18872 21560 18872 0 _0065_
rlabel metal2 19320 15456 19320 15456 0 _0066_
rlabel metal2 8008 22456 8008 22456 0 _0067_
rlabel metal2 5320 23408 5320 23408 0 _0068_
rlabel metal2 7672 23184 7672 23184 0 _0069_
rlabel metal2 3696 23688 3696 23688 0 _0070_
rlabel metal3 5488 24808 5488 24808 0 _0071_
rlabel metal2 14168 19208 14168 19208 0 _0072_
rlabel metal2 13496 19264 13496 19264 0 _0073_
rlabel metal3 6776 20552 6776 20552 0 _0074_
rlabel metal2 14728 21952 14728 21952 0 _0075_
rlabel metal2 20776 16016 20776 16016 0 _0076_
rlabel metal2 14952 21392 14952 21392 0 _0077_
rlabel metal2 25480 18144 25480 18144 0 _0078_
rlabel metal2 15176 21336 15176 21336 0 _0079_
rlabel metal3 14056 21560 14056 21560 0 _0080_
rlabel metal3 23352 16744 23352 16744 0 _0081_
rlabel metal3 12600 14280 12600 14280 0 _0082_
rlabel metal2 30072 25200 30072 25200 0 _0083_
rlabel metal2 21784 11648 21784 11648 0 _0084_
rlabel metal2 21448 12992 21448 12992 0 _0085_
rlabel metal2 21952 11368 21952 11368 0 _0086_
rlabel metal2 19656 14280 19656 14280 0 _0087_
rlabel metal2 19880 15008 19880 15008 0 _0088_
rlabel metal2 24360 16184 24360 16184 0 _0089_
rlabel metal3 25144 24696 25144 24696 0 _0090_
rlabel metal2 19432 15904 19432 15904 0 _0091_
rlabel metal2 19096 15568 19096 15568 0 _0092_
rlabel metal2 23912 13720 23912 13720 0 _0093_
rlabel metal3 26152 11368 26152 11368 0 _0094_
rlabel metal2 19768 11144 19768 11144 0 _0095_
rlabel metal3 19880 15288 19880 15288 0 _0096_
rlabel metal2 18536 15848 18536 15848 0 _0097_
rlabel metal3 8064 15288 8064 15288 0 _0098_
rlabel metal2 5656 15680 5656 15680 0 _0099_
rlabel metal2 10192 16856 10192 16856 0 _0100_
rlabel metal2 5320 15232 5320 15232 0 _0101_
rlabel metal3 6552 16296 6552 16296 0 _0102_
rlabel metal2 5096 19600 5096 19600 0 _0103_
rlabel metal3 6832 15848 6832 15848 0 _0104_
rlabel metal2 6944 16072 6944 16072 0 _0105_
rlabel metal2 7784 16520 7784 16520 0 _0106_
rlabel metal3 4424 21560 4424 21560 0 _0107_
rlabel metal3 9688 21000 9688 21000 0 _0108_
rlabel metal2 9912 21672 9912 21672 0 _0109_
rlabel metal2 10360 22680 10360 22680 0 _0110_
rlabel metal2 13440 22344 13440 22344 0 _0111_
rlabel metal2 13720 19656 13720 19656 0 _0112_
rlabel metal2 14168 18984 14168 18984 0 _0113_
rlabel metal3 13328 24024 13328 24024 0 _0114_
rlabel metal2 13944 17136 13944 17136 0 _0115_
rlabel metal3 17304 15176 17304 15176 0 _0116_
rlabel metal2 9072 22232 9072 22232 0 _0117_
rlabel metal2 7784 21224 7784 21224 0 _0118_
rlabel metal2 6440 21840 6440 21840 0 _0119_
rlabel metal2 7896 21112 7896 21112 0 _0120_
rlabel metal2 8456 6720 8456 6720 0 _0121_
rlabel metal3 10248 7560 10248 7560 0 _0122_
rlabel metal2 10584 7896 10584 7896 0 _0123_
rlabel metal3 19824 11256 19824 11256 0 _0124_
rlabel metal2 15400 6440 15400 6440 0 _0125_
rlabel metal3 10248 11144 10248 11144 0 _0126_
rlabel metal2 11480 11480 11480 11480 0 _0127_
rlabel metal2 12600 11704 12600 11704 0 _0128_
rlabel metal2 11928 11368 11928 11368 0 _0129_
rlabel metal2 12600 13552 12600 13552 0 _0130_
rlabel metal2 12264 10248 12264 10248 0 _0131_
rlabel metal3 11032 13944 11032 13944 0 _0132_
rlabel metal2 12320 14504 12320 14504 0 _0133_
rlabel metal2 11592 14952 11592 14952 0 _0134_
rlabel metal2 7448 12152 7448 12152 0 _0135_
rlabel metal2 8176 12152 8176 12152 0 _0136_
rlabel metal3 6944 10808 6944 10808 0 _0137_
rlabel metal2 4984 7840 4984 7840 0 _0138_
rlabel metal2 10024 7168 10024 7168 0 _0139_
rlabel metal2 15848 6440 15848 6440 0 _0140_
rlabel metal2 10080 9016 10080 9016 0 _0141_
rlabel metal2 8680 10304 8680 10304 0 _0142_
rlabel metal2 7112 10976 7112 10976 0 _0143_
rlabel metal2 8344 10920 8344 10920 0 _0144_
rlabel metal2 7336 11704 7336 11704 0 _0145_
rlabel metal2 8120 15148 8120 15148 0 _0146_
rlabel metal3 9688 15400 9688 15400 0 _0147_
rlabel metal3 10976 15176 10976 15176 0 _0148_
rlabel metal2 8792 12544 8792 12544 0 _0149_
rlabel metal2 8568 10976 8568 10976 0 _0150_
rlabel metal2 9576 11704 9576 11704 0 _0151_
rlabel metal2 9576 10472 9576 10472 0 _0152_
rlabel metal2 10024 9632 10024 9632 0 _0153_
rlabel metal2 13944 9408 13944 9408 0 _0154_
rlabel metal2 20048 12152 20048 12152 0 _0155_
rlabel metal2 14504 7840 14504 7840 0 _0156_
rlabel metal2 14616 7000 14616 7000 0 _0157_
rlabel metal3 14616 8232 14616 8232 0 _0158_
rlabel metal2 13608 9128 13608 9128 0 _0159_
rlabel metal2 13608 6104 13608 6104 0 _0160_
rlabel metal3 19768 22232 19768 22232 0 _0161_
rlabel metal3 27384 29400 27384 29400 0 _0162_
rlabel metal2 27384 29512 27384 29512 0 _0163_
rlabel metal2 27720 30128 27720 30128 0 _0164_
rlabel metal3 27776 28392 27776 28392 0 _0165_
rlabel metal2 28392 29848 28392 29848 0 _0166_
rlabel metal3 22960 29512 22960 29512 0 _0167_
rlabel metal2 17640 29288 17640 29288 0 _0168_
rlabel metal3 18312 30128 18312 30128 0 _0169_
rlabel metal2 17192 38192 17192 38192 0 _0170_
rlabel metal2 16184 38080 16184 38080 0 _0171_
rlabel metal2 15400 31976 15400 31976 0 _0172_
rlabel metal2 17416 32200 17416 32200 0 _0173_
rlabel metal2 13832 29624 13832 29624 0 _0174_
rlabel metal2 11592 37968 11592 37968 0 _0175_
rlabel metal2 14280 35336 14280 35336 0 _0176_
rlabel metal3 13832 31752 13832 31752 0 _0177_
rlabel metal2 18144 30072 18144 30072 0 _0178_
rlabel metal2 31416 32256 31416 32256 0 _0179_
rlabel metal3 29848 30968 29848 30968 0 _0180_
rlabel metal3 23072 30072 23072 30072 0 _0181_
rlabel metal2 19096 29736 19096 29736 0 _0182_
rlabel metal2 19768 23352 19768 23352 0 _0183_
rlabel metal2 20104 22232 20104 22232 0 _0184_
rlabel metal3 17052 22120 17052 22120 0 _0185_
rlabel metal3 21448 19880 21448 19880 0 _0186_
rlabel metal2 21336 5208 21336 5208 0 _0187_
rlabel metal2 7672 17248 7672 17248 0 _0188_
rlabel metal2 9128 19264 9128 19264 0 _0189_
rlabel metal3 8736 19096 8736 19096 0 _0190_
rlabel metal2 19656 17976 19656 17976 0 _0191_
rlabel metal2 26376 20832 26376 20832 0 _0192_
rlabel metal3 23352 11928 23352 11928 0 _0193_
rlabel metal2 23912 16296 23912 16296 0 _0194_
rlabel metal2 23128 15904 23128 15904 0 _0195_
rlabel metal3 22680 15512 22680 15512 0 _0196_
rlabel metal3 27720 15848 27720 15848 0 _0197_
rlabel metal2 30968 29344 30968 29344 0 _0198_
rlabel metal2 21672 5544 21672 5544 0 _0199_
rlabel metal2 17752 19880 17752 19880 0 _0200_
rlabel metal2 22568 24696 22568 24696 0 _0201_
rlabel metal2 22904 25088 22904 25088 0 _0202_
rlabel metal2 28168 32984 28168 32984 0 _0203_
rlabel metal3 16968 5768 16968 5768 0 _0204_
rlabel metal2 17528 6160 17528 6160 0 _0205_
rlabel metal2 7672 6608 7672 6608 0 _0206_
rlabel metal2 18984 19488 18984 19488 0 _0207_
rlabel metal2 15176 22400 15176 22400 0 _0208_
rlabel metal2 10248 5656 10248 5656 0 _0209_
rlabel metal2 5880 5152 5880 5152 0 _0210_
rlabel metal3 6160 6776 6160 6776 0 _0211_
rlabel metal2 6160 4088 6160 4088 0 _0212_
rlabel metal2 8848 5320 8848 5320 0 _0213_
rlabel metal2 18144 22120 18144 22120 0 _0214_
rlabel metal2 34888 6608 34888 6608 0 _0215_
rlabel metal2 39256 8680 39256 8680 0 _0216_
rlabel metal2 35896 5880 35896 5880 0 _0217_
rlabel metal2 36960 6776 36960 6776 0 _0218_
rlabel metal2 37128 7280 37128 7280 0 _0219_
rlabel metal2 29848 15204 29848 15204 0 _0220_
rlabel metal2 23240 11424 23240 11424 0 _0221_
rlabel metal2 22456 10696 22456 10696 0 _0222_
rlabel metal3 25928 12936 25928 12936 0 _0223_
rlabel metal3 30464 12936 30464 12936 0 _0224_
rlabel metal3 31696 15512 31696 15512 0 _0225_
rlabel metal2 22568 23072 22568 23072 0 _0226_
rlabel metal3 30408 12824 30408 12824 0 _0227_
rlabel metal2 26712 10640 26712 10640 0 _0228_
rlabel metal3 28392 7448 28392 7448 0 _0229_
rlabel metal2 39032 7504 39032 7504 0 _0230_
rlabel metal2 38920 8316 38920 8316 0 _0231_
rlabel metal2 36344 8176 36344 8176 0 _0232_
rlabel metal3 36792 9128 36792 9128 0 _0233_
rlabel metal2 29792 8120 29792 8120 0 _0234_
rlabel metal3 33376 7560 33376 7560 0 _0235_
rlabel metal3 29120 7336 29120 7336 0 _0236_
rlabel metal2 26376 7560 26376 7560 0 _0237_
rlabel metal3 29456 10584 29456 10584 0 _0238_
rlabel metal2 26712 7448 26712 7448 0 _0239_
rlabel metal2 28504 10584 28504 10584 0 _0240_
rlabel metal2 24584 30184 24584 30184 0 _0241_
rlabel metal2 37128 14112 37128 14112 0 _0242_
rlabel metal2 37016 9968 37016 9968 0 _0243_
rlabel metal3 31192 7448 31192 7448 0 _0244_
rlabel metal3 29848 10024 29848 10024 0 _0245_
rlabel metal2 29512 8512 29512 8512 0 _0246_
rlabel metal2 39032 9352 39032 9352 0 _0247_
rlabel metal2 31976 7504 31976 7504 0 _0248_
rlabel metal2 31136 9128 31136 9128 0 _0249_
rlabel metal2 30184 8400 30184 8400 0 _0250_
rlabel metal2 29624 8960 29624 8960 0 _0251_
rlabel metal2 23464 22512 23464 22512 0 _0252_
rlabel metal2 25592 7056 25592 7056 0 _0253_
rlabel metal2 30968 7896 30968 7896 0 _0254_
rlabel metal2 31640 8512 31640 8512 0 _0255_
rlabel metal3 31752 7672 31752 7672 0 _0256_
rlabel metal2 31192 8064 31192 8064 0 _0257_
rlabel metal2 30800 7560 30800 7560 0 _0258_
rlabel metal2 24472 7728 24472 7728 0 _0259_
rlabel metal2 33432 28280 33432 28280 0 _0260_
rlabel metal2 38920 5880 38920 5880 0 _0261_
rlabel metal3 27832 9800 27832 9800 0 _0262_
rlabel metal3 28392 9688 28392 9688 0 _0263_
rlabel metal3 35000 10472 35000 10472 0 _0264_
rlabel metal2 31640 12432 31640 12432 0 _0265_
rlabel metal2 33600 9240 33600 9240 0 _0266_
rlabel metal3 33152 10584 33152 10584 0 _0267_
rlabel metal2 31864 9856 31864 9856 0 _0268_
rlabel metal2 31752 10640 31752 10640 0 _0269_
rlabel metal2 33208 11368 33208 11368 0 _0270_
rlabel metal2 33096 11032 33096 11032 0 _0271_
rlabel metal2 32424 10024 32424 10024 0 _0272_
rlabel metal2 33320 7644 33320 7644 0 _0273_
rlabel metal2 29176 34496 29176 34496 0 _0274_
rlabel metal2 35896 16352 35896 16352 0 _0275_
rlabel metal3 34160 15960 34160 15960 0 _0276_
rlabel metal2 34272 11928 34272 11928 0 _0277_
rlabel metal2 33432 12544 33432 12544 0 _0278_
rlabel metal2 33768 12600 33768 12600 0 _0279_
rlabel metal2 34440 13440 34440 13440 0 _0280_
rlabel metal2 33992 12208 33992 12208 0 _0281_
rlabel metal2 32088 12824 32088 12824 0 _0282_
rlabel metal3 32760 12712 32760 12712 0 _0283_
rlabel metal2 33152 13048 33152 13048 0 _0284_
rlabel metal2 32144 15512 32144 15512 0 _0285_
rlabel metal2 38696 11368 38696 11368 0 _0286_
rlabel metal3 36848 10808 36848 10808 0 _0287_
rlabel metal3 35448 9016 35448 9016 0 _0288_
rlabel metal2 39144 10360 39144 10360 0 _0289_
rlabel metal2 38584 11032 38584 11032 0 _0290_
rlabel metal2 39088 9688 39088 9688 0 _0291_
rlabel metal2 37968 10584 37968 10584 0 _0292_
rlabel metal2 38248 10136 38248 10136 0 _0293_
rlabel metal3 38192 9576 38192 9576 0 _0294_
rlabel metal2 34496 31416 34496 31416 0 _0295_
rlabel metal2 36456 26908 36456 26908 0 _0296_
rlabel metal2 38808 4368 38808 4368 0 _0297_
rlabel metal2 38360 16856 38360 16856 0 _0298_
rlabel metal2 37016 10752 37016 10752 0 _0299_
rlabel metal3 37744 18536 37744 18536 0 _0300_
rlabel metal3 36456 11144 36456 11144 0 _0301_
rlabel metal2 37128 11760 37128 11760 0 _0302_
rlabel metal2 38696 13608 38696 13608 0 _0303_
rlabel metal2 37464 12600 37464 12600 0 _0304_
rlabel metal2 37352 13216 37352 13216 0 _0305_
rlabel metal3 38024 13832 38024 13832 0 _0306_
rlabel metal2 37352 14168 37352 14168 0 _0307_
rlabel metal2 36120 22288 36120 22288 0 _0308_
rlabel metal2 30072 16352 30072 16352 0 _0309_
rlabel metal3 33712 22120 33712 22120 0 _0310_
rlabel metal2 24360 35728 24360 35728 0 _0311_
rlabel metal2 35168 27160 35168 27160 0 _0312_
rlabel metal2 37352 22792 37352 22792 0 _0313_
rlabel metal2 37016 23016 37016 23016 0 _0314_
rlabel metal2 37408 21000 37408 21000 0 _0315_
rlabel metal3 36120 27944 36120 27944 0 _0316_
rlabel metal2 36008 27160 36008 27160 0 _0317_
rlabel metal2 31360 27496 31360 27496 0 _0318_
rlabel metal2 37016 29848 37016 29848 0 _0319_
rlabel metal2 38416 23128 38416 23128 0 _0320_
rlabel metal2 36792 29008 36792 29008 0 _0321_
rlabel metal3 36624 26936 36624 26936 0 _0322_
rlabel metal3 37240 27048 37240 27048 0 _0323_
rlabel metal3 34832 31640 34832 31640 0 _0324_
rlabel metal2 30968 30744 30968 30744 0 _0325_
rlabel metal2 31752 34496 31752 34496 0 _0326_
rlabel metal3 32760 30968 32760 30968 0 _0327_
rlabel metal3 29232 31192 29232 31192 0 _0328_
rlabel metal2 37464 29680 37464 29680 0 _0329_
rlabel metal3 36344 29624 36344 29624 0 _0330_
rlabel metal2 35896 31248 35896 31248 0 _0331_
rlabel metal2 33432 36008 33432 36008 0 _0332_
rlabel metal3 36288 31864 36288 31864 0 _0333_
rlabel metal2 37632 29288 37632 29288 0 _0334_
rlabel metal2 36344 30240 36344 30240 0 _0335_
rlabel metal2 37352 31024 37352 31024 0 _0336_
rlabel metal2 34888 32928 34888 32928 0 _0337_
rlabel metal2 35336 32816 35336 32816 0 _0338_
rlabel metal2 35336 32536 35336 32536 0 _0339_
rlabel metal2 30856 31528 30856 31528 0 _0340_
rlabel metal2 31080 31752 31080 31752 0 _0341_
rlabel metal2 31528 31976 31528 31976 0 _0342_
rlabel metal2 30184 33096 30184 33096 0 _0343_
rlabel metal2 28616 32592 28616 32592 0 _0344_
rlabel metal2 29848 32816 29848 32816 0 _0345_
rlabel metal3 29848 32760 29848 32760 0 _0346_
rlabel metal2 31192 29120 31192 29120 0 _0347_
rlabel metal2 32424 31640 32424 31640 0 _0348_
rlabel metal2 31640 29904 31640 29904 0 _0349_
rlabel metal3 30912 30184 30912 30184 0 _0350_
rlabel metal2 31472 29624 31472 29624 0 _0351_
rlabel metal2 31304 29568 31304 29568 0 _0352_
rlabel metal2 25480 32760 25480 32760 0 _0353_
rlabel metal2 30128 31080 30128 31080 0 _0354_
rlabel metal3 28896 30744 28896 30744 0 _0355_
rlabel metal2 26824 32704 26824 32704 0 _0356_
rlabel metal2 25928 33432 25928 33432 0 _0357_
rlabel metal3 22400 23128 22400 23128 0 _0358_
rlabel metal2 22960 23352 22960 23352 0 _0359_
rlabel metal3 21896 37968 21896 37968 0 _0360_
rlabel metal2 20664 38304 20664 38304 0 _0361_
rlabel metal2 23688 36456 23688 36456 0 _0362_
rlabel metal3 25200 36344 25200 36344 0 _0363_
rlabel metal2 25200 36568 25200 36568 0 _0364_
rlabel metal2 18312 35896 18312 35896 0 _0365_
rlabel metal2 20272 38808 20272 38808 0 _0366_
rlabel metal2 22176 36456 22176 36456 0 _0367_
rlabel metal2 18088 38724 18088 38724 0 _0368_
rlabel metal2 20776 38696 20776 38696 0 _0369_
rlabel metal2 17864 34048 17864 34048 0 _0370_
rlabel metal2 22120 38136 22120 38136 0 _0371_
rlabel metal3 20104 37800 20104 37800 0 _0372_
rlabel metal2 16520 35280 16520 35280 0 _0373_
rlabel metal2 16856 37912 16856 37912 0 _0374_
rlabel metal2 19320 38808 19320 38808 0 _0375_
rlabel metal2 16632 38864 16632 38864 0 _0376_
rlabel metal2 16464 39032 16464 39032 0 _0377_
rlabel metal2 17416 37576 17416 37576 0 _0378_
rlabel metal2 17752 31976 17752 31976 0 _0379_
rlabel metal2 17640 38668 17640 38668 0 _0380_
rlabel metal2 18200 37688 18200 37688 0 _0381_
rlabel metal2 18424 35280 18424 35280 0 _0382_
rlabel metal2 18648 34384 18648 34384 0 _0383_
rlabel metal3 13888 34776 13888 34776 0 _0384_
rlabel metal3 17640 34888 17640 34888 0 _0385_
rlabel metal2 16184 34440 16184 34440 0 _0386_
rlabel metal2 17304 34384 17304 34384 0 _0387_
rlabel metal2 17528 33600 17528 33600 0 _0388_
rlabel metal3 17640 34104 17640 34104 0 _0389_
rlabel metal2 17920 32760 17920 32760 0 _0390_
rlabel metal3 19488 33208 19488 33208 0 _0391_
rlabel metal2 20104 33824 20104 33824 0 _0392_
rlabel metal2 21448 33320 21448 33320 0 _0393_
rlabel metal2 19880 32368 19880 32368 0 _0394_
rlabel metal3 20496 32760 20496 32760 0 _0395_
rlabel metal3 11872 38696 11872 38696 0 _0396_
rlabel metal2 12824 37744 12824 37744 0 _0397_
rlabel metal2 14280 32536 14280 32536 0 _0398_
rlabel metal2 14056 34944 14056 34944 0 _0399_
rlabel metal3 13384 37800 13384 37800 0 _0400_
rlabel metal3 12880 37464 12880 37464 0 _0401_
rlabel metal3 12936 37912 12936 37912 0 _0402_
rlabel metal2 13832 38360 13832 38360 0 _0403_
rlabel metal2 13720 25340 13720 25340 0 _0404_
rlabel metal2 10584 33712 10584 33712 0 _0405_
rlabel metal2 11592 35728 11592 35728 0 _0406_
rlabel metal2 13272 35840 13272 35840 0 _0407_
rlabel metal2 13496 34720 13496 34720 0 _0408_
rlabel metal2 13720 35728 13720 35728 0 _0409_
rlabel metal3 13384 35560 13384 35560 0 _0410_
rlabel metal2 17416 29848 17416 29848 0 _0411_
rlabel metal3 14392 34104 14392 34104 0 _0412_
rlabel metal2 16408 32200 16408 32200 0 _0413_
rlabel metal2 16240 30968 16240 30968 0 _0414_
rlabel metal2 16576 30968 16576 30968 0 _0415_
rlabel metal3 16800 31528 16800 31528 0 _0416_
rlabel metal2 16968 31472 16968 31472 0 _0417_
rlabel metal2 17136 30184 17136 30184 0 _0418_
rlabel metal2 17864 22344 17864 22344 0 _0419_
rlabel metal2 15960 22960 15960 22960 0 _0420_
rlabel metal2 19208 13776 19208 13776 0 _0421_
rlabel metal2 26040 12264 26040 12264 0 _0422_
rlabel metal2 27496 12488 27496 12488 0 _0423_
rlabel metal2 25480 12656 25480 12656 0 _0424_
rlabel metal2 28112 12152 28112 12152 0 _0425_
rlabel metal2 24080 9912 24080 9912 0 _0426_
rlabel metal2 25928 12488 25928 12488 0 _0427_
rlabel metal2 25760 12152 25760 12152 0 _0428_
rlabel metal2 25816 13048 25816 13048 0 _0429_
rlabel metal2 26544 12264 26544 12264 0 _0430_
rlabel metal2 31640 18536 31640 18536 0 _0431_
rlabel metal3 32760 19208 32760 19208 0 _0432_
rlabel metal2 37240 18144 37240 18144 0 _0433_
rlabel metal2 37240 17752 37240 17752 0 _0434_
rlabel metal2 24248 19936 24248 19936 0 _0435_
rlabel metal2 37016 18312 37016 18312 0 _0436_
rlabel metal2 33264 18200 33264 18200 0 _0437_
rlabel metal3 32480 19432 32480 19432 0 _0438_
rlabel metal2 19544 23632 19544 23632 0 _0439_
rlabel metal2 10472 29120 10472 29120 0 _0440_
rlabel metal2 9016 29736 9016 29736 0 _0441_
rlabel metal2 11816 30912 11816 30912 0 _0442_
rlabel metal2 10136 29344 10136 29344 0 _0443_
rlabel metal3 9520 29400 9520 29400 0 _0444_
rlabel metal2 8008 28728 8008 28728 0 _0445_
rlabel metal3 9016 28728 9016 28728 0 _0446_
rlabel metal3 9184 28616 9184 28616 0 _0447_
rlabel metal2 10304 27944 10304 27944 0 _0448_
rlabel metal2 11256 28392 11256 28392 0 _0449_
rlabel metal2 10472 33152 10472 33152 0 _0450_
rlabel metal2 10024 33264 10024 33264 0 _0451_
rlabel metal2 11816 29400 11816 29400 0 _0452_
rlabel metal2 10864 16968 10864 16968 0 _0453_
rlabel metal2 9912 16408 9912 16408 0 _0454_
rlabel metal2 11200 20328 11200 20328 0 _0455_
rlabel metal2 10472 29904 10472 29904 0 _0456_
rlabel metal2 8904 32592 8904 32592 0 _0457_
rlabel metal2 8456 31472 8456 31472 0 _0458_
rlabel metal3 9800 30184 9800 30184 0 _0459_
rlabel metal2 11592 28784 11592 28784 0 _0460_
rlabel metal3 12768 28616 12768 28616 0 _0461_
rlabel metal2 8792 30240 8792 30240 0 _0462_
rlabel metal3 11032 29624 11032 29624 0 _0463_
rlabel metal2 11032 29120 11032 29120 0 _0464_
rlabel metal2 13720 28952 13720 28952 0 _0465_
rlabel metal2 14168 29400 14168 29400 0 _0466_
rlabel metal2 14056 28896 14056 28896 0 _0467_
rlabel metal2 30072 23520 30072 23520 0 _0468_
rlabel metal2 30296 22736 30296 22736 0 _0469_
rlabel metal2 29960 22736 29960 22736 0 _0470_
rlabel metal3 13440 23688 13440 23688 0 _0471_
rlabel metal2 15624 23184 15624 23184 0 _0472_
rlabel metal2 18872 18872 18872 18872 0 _0473_
rlabel metal2 26600 25872 26600 25872 0 _0474_
rlabel metal2 26152 24696 26152 24696 0 _0475_
rlabel metal3 27048 23800 27048 23800 0 _0476_
rlabel metal2 32312 21504 32312 21504 0 _0477_
rlabel metal2 31864 21784 31864 21784 0 _0478_
rlabel metal2 29176 25648 29176 25648 0 _0479_
rlabel metal2 28504 29456 28504 29456 0 _0480_
rlabel metal3 28896 25816 28896 25816 0 _0481_
rlabel metal2 29400 25088 29400 25088 0 _0482_
rlabel metal3 29176 24696 29176 24696 0 _0483_
rlabel metal2 27608 24752 27608 24752 0 _0484_
rlabel metal2 27328 20776 27328 20776 0 _0485_
rlabel metal2 27496 21728 27496 21728 0 _0486_
rlabel metal2 28168 27888 28168 27888 0 _0487_
rlabel metal2 28336 28056 28336 28056 0 _0488_
rlabel metal2 26712 27776 26712 27776 0 _0489_
rlabel metal2 27552 26936 27552 26936 0 _0490_
rlabel metal2 26264 25928 26264 25928 0 _0491_
rlabel metal2 27272 25816 27272 25816 0 _0492_
rlabel metal2 30184 27440 30184 27440 0 _0493_
rlabel metal3 29232 28504 29232 28504 0 _0494_
rlabel metal2 29120 27272 29120 27272 0 _0495_
rlabel metal2 29848 24528 29848 24528 0 _0496_
rlabel metal2 28952 24920 28952 24920 0 _0497_
rlabel metal2 28728 25648 28728 25648 0 _0498_
rlabel metal3 26712 25984 26712 25984 0 _0499_
rlabel metal2 27720 23576 27720 23576 0 _0500_
rlabel metal2 3192 9744 3192 9744 0 _0501_
rlabel metal2 3304 24416 3304 24416 0 _0502_
rlabel metal2 3192 22960 3192 22960 0 _0503_
rlabel metal2 2912 8120 2912 8120 0 _0504_
rlabel metal2 16744 19488 16744 19488 0 _0505_
rlabel metal2 3640 15736 3640 15736 0 _0506_
rlabel metal2 4424 15512 4424 15512 0 _0507_
rlabel metal2 3080 16016 3080 16016 0 _0508_
rlabel metal2 3304 15568 3304 15568 0 _0509_
rlabel metal2 3976 20776 3976 20776 0 _0510_
rlabel metal2 4312 18928 4312 18928 0 _0511_
rlabel metal2 3080 20804 3080 20804 0 _0512_
rlabel metal2 8456 22008 8456 22008 0 _0513_
rlabel metal2 5096 22512 5096 22512 0 _0514_
rlabel metal2 3696 23912 3696 23912 0 _0515_
rlabel metal2 5656 23968 5656 23968 0 _0516_
rlabel metal2 2688 24696 2688 24696 0 _0517_
rlabel metal2 4088 24192 4088 24192 0 _0518_
rlabel metal2 4312 25088 4312 25088 0 _0519_
rlabel metal3 37296 18424 37296 18424 0 _0520_
rlabel metal2 37016 16408 37016 16408 0 _0521_
rlabel metal2 36680 17304 36680 17304 0 _0522_
rlabel metal3 36736 17416 36736 17416 0 _0523_
rlabel metal3 35000 18312 35000 18312 0 _0524_
rlabel metal2 33096 18536 33096 18536 0 _0525_
rlabel metal2 16632 20104 16632 20104 0 _0526_
rlabel metal3 15120 22232 15120 22232 0 _0527_
rlabel metal3 18368 11368 18368 11368 0 _0528_
rlabel metal2 19096 13216 19096 13216 0 _0529_
rlabel metal3 18368 11592 18368 11592 0 _0530_
rlabel metal2 17416 18312 17416 18312 0 _0531_
rlabel metal2 17640 15204 17640 15204 0 _0532_
rlabel metal2 17920 10696 17920 10696 0 _0533_
rlabel metal2 18424 10472 18424 10472 0 _0534_
rlabel metal2 19656 11536 19656 11536 0 _0535_
rlabel metal2 18816 15512 18816 15512 0 _0536_
rlabel metal2 18648 12600 18648 12600 0 _0537_
rlabel metal2 19768 17696 19768 17696 0 _0538_
rlabel metal3 18312 14728 18312 14728 0 _0539_
rlabel metal2 18200 14616 18200 14616 0 _0540_
rlabel metal2 17864 15736 17864 15736 0 _0541_
rlabel metal2 18368 16968 18368 16968 0 _0542_
rlabel metal3 20664 19096 20664 19096 0 _0543_
rlabel metal2 19320 18704 19320 18704 0 _0544_
rlabel metal2 19096 23296 19096 23296 0 _0545_
rlabel metal2 19992 21224 19992 21224 0 _0546_
rlabel metal2 20552 20132 20552 20132 0 _0547_
rlabel metal2 23240 19600 23240 19600 0 _0548_
rlabel metal3 22960 19880 22960 19880 0 _0549_
rlabel metal2 22120 19712 22120 19712 0 _0550_
rlabel metal2 23688 17136 23688 17136 0 _0551_
rlabel metal2 23464 17304 23464 17304 0 _0552_
rlabel metal2 18872 20944 18872 20944 0 clk
rlabel metal3 28728 27832 28728 27832 0 clknet_0_clk
rlabel metal2 1904 7448 1904 7448 0 clknet_3_0__leaf_clk
rlabel metal2 1848 19208 1848 19208 0 clknet_3_1__leaf_clk
rlabel via2 22904 10584 22904 10584 0 clknet_3_2__leaf_clk
rlabel metal3 24864 20776 24864 20776 0 clknet_3_3__leaf_clk
rlabel metal2 1848 26992 1848 26992 0 clknet_3_4__leaf_clk
rlabel metal2 2856 30184 2856 30184 0 clknet_3_5__leaf_clk
rlabel metal2 34776 26992 34776 26992 0 clknet_3_6__leaf_clk
rlabel metal2 24472 39592 24472 39592 0 clknet_3_7__leaf_clk
rlabel metal2 4760 2184 4760 2184 0 gpio_ready
rlabel metal2 39480 2086 39480 2086 0 io_in[0]
rlabel metal2 38136 2058 38136 2058 0 io_in[1]
rlabel metal3 35168 4424 35168 4424 0 io_in[2]
rlabel metal3 33264 3416 33264 3416 0 io_in[3]
rlabel metal3 35616 4984 35616 4984 0 io_in[4]
rlabel metal3 8176 3640 8176 3640 0 io_out[10]
rlabel metal2 7224 2478 7224 2478 0 io_out[11]
rlabel metal2 5992 4312 5992 4312 0 io_out[12]
rlabel metal3 16912 3416 16912 3416 0 io_out[5]
rlabel metal3 14392 3416 14392 3416 0 io_out[6]
rlabel metal2 12600 2058 12600 2058 0 io_out[7]
rlabel metal2 11256 2198 11256 2198 0 io_out[8]
rlabel metal2 9912 2058 9912 2058 0 io_out[9]
rlabel metal2 5544 3864 5544 3864 0 net1
rlabel metal2 4984 5208 4984 5208 0 net10
rlabel metal2 14392 4592 14392 4592 0 net11
rlabel metal2 14112 17640 14112 17640 0 net12
rlabel metal2 13832 4592 13832 4592 0 net13
rlabel metal3 6944 20664 6944 20664 0 net14
rlabel metal2 10920 6272 10920 6272 0 net15
rlabel metal2 22008 2030 22008 2030 0 net16
rlabel metal2 20664 2030 20664 2030 0 net17
rlabel metal2 19320 2030 19320 2030 0 net18
rlabel metal2 17976 2058 17976 2058 0 net19
rlabel metal2 13160 5992 13160 5992 0 net2
rlabel metal3 17024 4424 17024 4424 0 net20
rlabel metal2 32648 4088 32648 4088 0 net21
rlabel metal2 31080 15624 31080 15624 0 net22
rlabel metal2 30464 29960 30464 29960 0 net23
rlabel metal2 21336 29008 21336 29008 0 net24
rlabel metal2 38024 9072 38024 9072 0 net25
rlabel metal2 32312 23072 32312 23072 0 net26
rlabel metal2 33656 21840 33656 21840 0 net27
rlabel metal2 38528 9016 38528 9016 0 net28
rlabel metal2 32200 4648 32200 4648 0 net29
rlabel metal3 22904 15960 22904 15960 0 net3
rlabel metal3 30184 14392 30184 14392 0 net30
rlabel metal2 31304 4312 31304 4312 0 net31
rlabel metal2 39144 5096 39144 5096 0 net32
rlabel metal2 35784 4872 35784 4872 0 net33
rlabel metal2 33320 13216 33320 13216 0 net34
rlabel metal2 32816 15288 32816 15288 0 net35
rlabel metal2 32592 16856 32592 16856 0 net36
rlabel metal2 33768 16968 33768 16968 0 net37
rlabel metal2 37688 6384 37688 6384 0 net38
rlabel metal2 38360 14056 38360 14056 0 net39
rlabel metal3 32144 16968 32144 16968 0 net4
rlabel metal2 35224 4760 35224 4760 0 net40
rlabel metal2 39032 5936 39032 5936 0 net41
rlabel metal3 32984 6552 32984 6552 0 net5
rlabel metal3 34832 5768 34832 5768 0 net6
rlabel metal2 3808 3416 3808 3416 0 net7
rlabel metal2 8680 4424 8680 4424 0 net8
rlabel metal2 15456 20104 15456 20104 0 net9
rlabel metal2 3192 2086 3192 2086 0 rst
rlabel metal2 18872 32704 18872 32704 0 solo_squash.ballDirX
rlabel metal2 36120 24360 36120 24360 0 solo_squash.ballDirY
rlabel metal2 23408 34664 23408 34664 0 solo_squash.ballX\[0\]
rlabel metal3 21560 35560 21560 35560 0 solo_squash.ballX\[1\]
rlabel metal2 21336 39200 21336 39200 0 solo_squash.ballX\[2\]
rlabel metal2 17752 39312 17752 39312 0 solo_squash.ballX\[3\]
rlabel metal2 12152 35056 12152 35056 0 solo_squash.ballX\[4\]
rlabel metal2 20216 32872 20216 32872 0 solo_squash.ballX\[5\]
rlabel metal3 12040 38808 12040 38808 0 solo_squash.ballX\[6\]
rlabel metal2 8456 35000 8456 35000 0 solo_squash.ballX\[7\]
rlabel metal2 6440 30520 6440 30520 0 solo_squash.ballX\[8\]
rlabel metal2 36456 22792 36456 22792 0 solo_squash.ballY\[0\]
rlabel metal2 38920 23464 38920 23464 0 solo_squash.ballY\[1\]
rlabel metal2 39256 27384 39256 27384 0 solo_squash.ballY\[2\]
rlabel metal2 36456 29736 36456 29736 0 solo_squash.ballY\[3\]
rlabel metal2 34440 34496 34440 34496 0 solo_squash.ballY\[4\]
rlabel metal2 31304 33264 31304 33264 0 solo_squash.ballY\[5\]
rlabel metal2 31640 27160 31640 27160 0 solo_squash.ballY\[6\]
rlabel metal2 28112 33992 28112 33992 0 solo_squash.ballY\[7\]
rlabel metal2 8904 8064 8904 8064 0 solo_squash.h\[0\]
rlabel metal3 5376 8120 5376 8120 0 solo_squash.h\[1\]
rlabel metal2 6328 12040 6328 12040 0 solo_squash.h\[2\]
rlabel metal2 7224 13272 7224 13272 0 solo_squash.h\[3\]
rlabel metal2 8568 18480 8568 18480 0 solo_squash.h\[4\]
rlabel metal2 7672 21112 7672 21112 0 solo_squash.h\[5\]
rlabel metal2 11424 24024 11424 24024 0 solo_squash.h\[6\]
rlabel metal2 8456 19600 8456 19600 0 solo_squash.h\[7\]
rlabel metal2 6440 25872 6440 25872 0 solo_squash.h\[8\]
rlabel metal2 7728 25368 7728 25368 0 solo_squash.h\[9\]
rlabel metal2 18984 23184 18984 23184 0 solo_squash.hit
rlabel metal3 12208 28392 12208 28392 0 solo_squash.inBallX
rlabel metal2 14392 21728 14392 21728 0 solo_squash.inBallY
rlabel metal2 12488 22680 12488 22680 0 solo_squash.inPaddle
rlabel metal2 19656 5040 19656 5040 0 solo_squash.offset\[0\]
rlabel metal2 15400 6048 15400 6048 0 solo_squash.offset\[1\]
rlabel metal3 13440 5992 13440 5992 0 solo_squash.offset\[2\]
rlabel metal2 5600 5992 5600 5992 0 solo_squash.offset\[3\]
rlabel metal2 8120 5992 8120 5992 0 solo_squash.offset\[4\]
rlabel metal2 23128 10360 23128 10360 0 solo_squash.paddle\[0\]
rlabel metal2 29288 4760 29288 4760 0 solo_squash.paddle\[1\]
rlabel metal2 29064 5096 29064 5096 0 solo_squash.paddle\[2\]
rlabel metal3 26852 5208 26852 5208 0 solo_squash.paddle\[3\]
rlabel metal2 26152 8232 26152 8232 0 solo_squash.paddle\[4\]
rlabel metal3 33992 8232 33992 8232 0 solo_squash.paddle\[5\]
rlabel metal2 31752 16184 31752 16184 0 solo_squash.paddle\[6\]
rlabel metal2 39368 5992 39368 5992 0 solo_squash.paddle\[7\]
rlabel metal2 38584 15624 38584 15624 0 solo_squash.paddle\[8\]
rlabel metal3 21560 7448 21560 7448 0 solo_squash.v\[0\]
rlabel metal3 17640 8344 17640 8344 0 solo_squash.v\[1\]
rlabel metal3 14224 11480 14224 11480 0 solo_squash.v\[2\]
rlabel metal2 12712 15512 12712 15512 0 solo_squash.v\[3\]
rlabel metal2 19544 17248 19544 17248 0 solo_squash.v\[4\]
rlabel metal2 25928 20160 25928 20160 0 solo_squash.v\[5\]
rlabel metal3 24080 26152 24080 26152 0 solo_squash.v\[6\]
rlabel metal2 25704 20944 25704 20944 0 solo_squash.v\[7\]
rlabel metal2 24584 24080 24584 24080 0 solo_squash.v\[8\]
rlabel metal2 25592 16800 25592 16800 0 solo_squash.v\[9\]
<< properties >>
string FIXED_BBOX 0 0 41437 45021
<< end >>
