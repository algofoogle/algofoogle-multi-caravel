VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_cpu
  CLASS BLOCK ;
  FOREIGN user_proj_cpu ;
  ORIGIN 0.000 0.000 ;
  SIZE 1162.320 BY 1180.240 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 1176.240 782.320 1180.240 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 893.760 1176.240 894.320 1180.240 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 904.960 1176.240 905.520 1180.240 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 916.160 1176.240 916.720 1180.240 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 1176.240 927.920 1180.240 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 938.560 1176.240 939.120 1180.240 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 949.760 1176.240 950.320 1180.240 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 1176.240 961.520 1180.240 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 972.160 1176.240 972.720 1180.240 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 1176.240 983.920 1180.240 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 1176.240 995.120 1180.240 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 792.960 1176.240 793.520 1180.240 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1005.760 1176.240 1006.320 1180.240 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1016.960 1176.240 1017.520 1180.240 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1028.160 1176.240 1028.720 1180.240 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1039.360 1176.240 1039.920 1180.240 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1050.560 1176.240 1051.120 1180.240 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1061.760 1176.240 1062.320 1180.240 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1072.960 1176.240 1073.520 1180.240 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1084.160 1176.240 1084.720 1180.240 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1095.360 1176.240 1095.920 1180.240 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1106.560 1176.240 1107.120 1180.240 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 804.160 1176.240 804.720 1180.240 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1117.760 1176.240 1118.320 1180.240 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1128.960 1176.240 1129.520 1180.240 ;
    END
  END io_in[31]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 815.360 1176.240 815.920 1180.240 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 826.560 1176.240 827.120 1180.240 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 1176.240 838.320 1180.240 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 848.960 1176.240 849.520 1180.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 860.160 1176.240 860.720 1180.240 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 871.360 1176.240 871.920 1180.240 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 882.560 1176.240 883.120 1180.240 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 1176.240 423.920 1180.240 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 1176.240 535.920 1180.240 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 546.560 1176.240 547.120 1180.240 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 1176.240 558.320 1180.240 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 568.960 1176.240 569.520 1180.240 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 1176.240 580.720 1180.240 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 1176.240 591.920 1180.240 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 1176.240 603.120 1180.240 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 613.760 1176.240 614.320 1180.240 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 1176.240 625.520 1180.240 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 636.160 1176.240 636.720 1180.240 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 1176.240 435.120 1180.240 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 647.360 1176.240 647.920 1180.240 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 1176.240 659.120 1180.240 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 669.760 1176.240 670.320 1180.240 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 1176.240 681.520 1180.240 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 1176.240 692.720 1180.240 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 703.360 1176.240 703.920 1180.240 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 714.560 1176.240 715.120 1180.240 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 1176.240 726.320 1180.240 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 736.960 1176.240 737.520 1180.240 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 748.160 1176.240 748.720 1180.240 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 1176.240 446.320 1180.240 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 1176.240 759.920 1180.240 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 770.560 1176.240 771.120 1180.240 ;
    END
  END io_oeb[31]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 1176.240 457.520 1180.240 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 1176.240 468.720 1180.240 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 479.360 1176.240 479.920 1180.240 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 1176.240 491.120 1180.240 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 501.760 1176.240 502.320 1180.240 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 512.960 1176.240 513.520 1180.240 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 1176.240 524.720 1180.240 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 1176.240 65.520 1180.240 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 1176.240 177.520 1180.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 1176.240 188.720 1180.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 1176.240 199.920 1180.240 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 1176.240 211.120 1180.240 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1176.240 222.320 1180.240 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 232.960 1176.240 233.520 1180.240 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 1176.240 244.720 1180.240 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 1176.240 255.920 1180.240 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 1176.240 267.120 1180.240 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 1176.240 278.320 1180.240 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 1176.240 76.720 1180.240 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 1176.240 289.520 1180.240 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 300.160 1176.240 300.720 1180.240 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 1176.240 311.920 1180.240 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 1176.240 323.120 1180.240 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 1176.240 334.320 1180.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 344.960 1176.240 345.520 1180.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 1176.240 356.720 1180.240 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 1176.240 367.920 1180.240 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 1176.240 379.120 1180.240 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 1176.240 390.320 1180.240 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 1176.240 87.920 1180.240 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 1176.240 401.520 1180.240 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 412.160 1176.240 412.720 1180.240 ;
    END
  END io_out[31]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 1176.240 99.120 1180.240 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 1176.240 110.320 1180.240 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 1176.240 121.520 1180.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 1176.240 132.720 1180.240 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 1176.240 143.920 1180.240 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 1176.240 155.120 1180.240 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 1176.240 166.320 1180.240 ;
    END
  END io_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1164.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1164.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1164.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 1176.240 31.920 1180.240 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 1162.205 1155.710 1164.670 ;
        RECT 6.290 1162.080 718.305 1162.205 ;
      LAYER Pwell ;
        RECT 6.290 1158.560 1155.710 1162.080 ;
      LAYER Nwell ;
        RECT 6.290 1158.435 96.705 1158.560 ;
        RECT 6.290 1154.365 1155.710 1158.435 ;
        RECT 6.290 1154.240 202.545 1154.365 ;
      LAYER Pwell ;
        RECT 6.290 1150.720 1155.710 1154.240 ;
      LAYER Nwell ;
        RECT 6.290 1150.595 223.265 1150.720 ;
        RECT 6.290 1146.525 1155.710 1150.595 ;
        RECT 6.290 1146.400 87.745 1146.525 ;
      LAYER Pwell ;
        RECT 6.290 1142.880 1155.710 1146.400 ;
      LAYER Nwell ;
        RECT 6.290 1142.755 342.760 1142.880 ;
        RECT 6.290 1138.685 1155.710 1142.755 ;
        RECT 6.290 1138.560 116.305 1138.685 ;
      LAYER Pwell ;
        RECT 6.290 1135.040 1155.710 1138.560 ;
      LAYER Nwell ;
        RECT 6.290 1134.915 137.025 1135.040 ;
        RECT 6.290 1130.845 1155.710 1134.915 ;
        RECT 6.290 1130.720 86.065 1130.845 ;
      LAYER Pwell ;
        RECT 6.290 1127.200 1155.710 1130.720 ;
      LAYER Nwell ;
        RECT 6.290 1127.075 68.145 1127.200 ;
        RECT 6.290 1123.005 1155.710 1127.075 ;
        RECT 6.290 1122.880 110.705 1123.005 ;
      LAYER Pwell ;
        RECT 6.290 1119.360 1155.710 1122.880 ;
      LAYER Nwell ;
        RECT 6.290 1119.235 141.505 1119.360 ;
        RECT 6.290 1115.165 1155.710 1119.235 ;
        RECT 6.290 1115.040 171.745 1115.165 ;
      LAYER Pwell ;
        RECT 6.290 1111.520 1155.710 1115.040 ;
      LAYER Nwell ;
        RECT 6.290 1111.395 69.825 1111.520 ;
        RECT 6.290 1107.335 1155.710 1111.395 ;
        RECT 6.290 1107.325 399.360 1107.335 ;
        RECT 6.290 1107.200 115.960 1107.325 ;
      LAYER Pwell ;
        RECT 6.290 1103.680 1155.710 1107.200 ;
      LAYER Nwell ;
        RECT 6.290 1103.555 217.105 1103.680 ;
        RECT 6.290 1103.545 462.080 1103.555 ;
        RECT 6.290 1099.485 1155.710 1103.545 ;
        RECT 6.290 1099.360 132.545 1099.485 ;
      LAYER Pwell ;
        RECT 6.290 1095.840 1155.710 1099.360 ;
      LAYER Nwell ;
        RECT 6.290 1095.715 177.345 1095.840 ;
        RECT 6.290 1095.705 418.400 1095.715 ;
        RECT 6.290 1091.655 1155.710 1095.705 ;
        RECT 6.290 1091.645 446.960 1091.655 ;
        RECT 6.290 1091.520 78.225 1091.645 ;
      LAYER Pwell ;
        RECT 6.290 1088.000 1155.710 1091.520 ;
      LAYER Nwell ;
        RECT 6.290 1087.875 60.305 1088.000 ;
        RECT 6.290 1087.865 420.640 1087.875 ;
        RECT 6.290 1083.815 1155.710 1087.865 ;
        RECT 6.290 1083.805 394.320 1083.815 ;
        RECT 6.290 1083.680 177.000 1083.805 ;
      LAYER Pwell ;
        RECT 6.290 1080.160 1155.710 1083.680 ;
      LAYER Nwell ;
        RECT 6.290 1080.035 146.200 1080.160 ;
        RECT 6.290 1080.025 452.000 1080.035 ;
        RECT 6.290 1075.975 1155.710 1080.025 ;
        RECT 6.290 1075.965 436.320 1075.975 ;
        RECT 6.290 1075.840 87.185 1075.965 ;
      LAYER Pwell ;
        RECT 6.290 1072.320 1155.710 1075.840 ;
      LAYER Nwell ;
        RECT 6.290 1072.195 68.145 1072.320 ;
        RECT 6.290 1072.185 384.240 1072.195 ;
        RECT 6.290 1068.125 1155.710 1072.185 ;
        RECT 6.290 1068.000 126.385 1068.125 ;
      LAYER Pwell ;
        RECT 6.290 1064.480 1155.710 1068.000 ;
      LAYER Nwell ;
        RECT 6.290 1064.355 148.225 1064.480 ;
        RECT 6.290 1060.295 1155.710 1064.355 ;
        RECT 6.290 1060.285 389.840 1060.295 ;
        RECT 6.290 1060.160 189.105 1060.285 ;
      LAYER Pwell ;
        RECT 6.290 1056.640 1155.710 1060.160 ;
      LAYER Nwell ;
        RECT 6.290 1056.515 67.240 1056.640 ;
        RECT 6.290 1056.505 409.440 1056.515 ;
        RECT 6.290 1052.445 1155.710 1056.505 ;
        RECT 6.290 1052.320 81.025 1052.445 ;
      LAYER Pwell ;
        RECT 6.290 1048.800 1155.710 1052.320 ;
      LAYER Nwell ;
        RECT 6.290 1048.675 146.760 1048.800 ;
        RECT 6.290 1048.665 389.280 1048.675 ;
        RECT 6.290 1044.605 1155.710 1048.665 ;
        RECT 6.290 1044.480 203.105 1044.605 ;
      LAYER Pwell ;
        RECT 6.290 1040.960 1155.710 1044.480 ;
      LAYER Nwell ;
        RECT 6.290 1040.835 70.945 1040.960 ;
        RECT 6.290 1040.825 384.800 1040.835 ;
        RECT 6.290 1036.765 1155.710 1040.825 ;
        RECT 6.290 1036.640 91.105 1036.765 ;
      LAYER Pwell ;
        RECT 6.290 1033.120 1155.710 1036.640 ;
      LAYER Nwell ;
        RECT 6.290 1032.995 137.025 1033.120 ;
        RECT 6.290 1028.925 1155.710 1032.995 ;
        RECT 6.290 1028.800 256.010 1028.925 ;
      LAYER Pwell ;
        RECT 6.290 1025.280 1155.710 1028.800 ;
      LAYER Nwell ;
        RECT 6.290 1025.155 419.265 1025.280 ;
        RECT 6.290 1021.085 1155.710 1025.155 ;
        RECT 6.290 1020.960 83.825 1021.085 ;
      LAYER Pwell ;
        RECT 6.290 1017.440 1155.710 1020.960 ;
      LAYER Nwell ;
        RECT 6.290 1017.315 64.225 1017.440 ;
        RECT 6.290 1013.245 1155.710 1017.315 ;
        RECT 6.290 1013.120 236.705 1013.245 ;
      LAYER Pwell ;
        RECT 6.290 1009.600 1155.710 1013.120 ;
      LAYER Nwell ;
        RECT 6.290 1009.475 61.080 1009.600 ;
        RECT 6.290 1005.405 1155.710 1009.475 ;
        RECT 6.290 1005.280 114.065 1005.405 ;
      LAYER Pwell ;
        RECT 6.290 1001.760 1155.710 1005.280 ;
      LAYER Nwell ;
        RECT 6.290 1001.635 73.185 1001.760 ;
        RECT 6.290 997.565 1155.710 1001.635 ;
        RECT 6.290 997.440 333.800 997.565 ;
      LAYER Pwell ;
        RECT 6.290 993.920 1155.710 997.440 ;
      LAYER Nwell ;
        RECT 6.290 993.795 73.745 993.920 ;
        RECT 6.290 989.725 1155.710 993.795 ;
        RECT 6.290 989.600 239.505 989.725 ;
      LAYER Pwell ;
        RECT 6.290 986.080 1155.710 989.600 ;
      LAYER Nwell ;
        RECT 6.290 985.955 140.040 986.080 ;
        RECT 6.290 981.885 1155.710 985.955 ;
        RECT 6.290 981.760 82.360 981.885 ;
      LAYER Pwell ;
        RECT 6.290 978.240 1155.710 981.760 ;
      LAYER Nwell ;
        RECT 6.290 978.115 269.745 978.240 ;
        RECT 6.290 974.045 1155.710 978.115 ;
        RECT 6.290 973.920 463.505 974.045 ;
      LAYER Pwell ;
        RECT 6.290 970.400 1155.710 973.920 ;
      LAYER Nwell ;
        RECT 6.290 970.275 99.505 970.400 ;
        RECT 6.290 966.205 1155.710 970.275 ;
        RECT 6.290 966.080 120.225 966.205 ;
      LAYER Pwell ;
        RECT 6.290 962.560 1155.710 966.080 ;
      LAYER Nwell ;
        RECT 6.290 962.435 143.745 962.560 ;
        RECT 6.290 958.365 1155.710 962.435 ;
        RECT 6.290 958.240 235.585 958.365 ;
      LAYER Pwell ;
        RECT 6.290 954.720 1155.710 958.240 ;
      LAYER Nwell ;
        RECT 6.290 954.595 216.545 954.720 ;
        RECT 6.290 950.525 1155.710 954.595 ;
        RECT 6.290 950.400 119.105 950.525 ;
      LAYER Pwell ;
        RECT 6.290 946.880 1155.710 950.400 ;
      LAYER Nwell ;
        RECT 6.290 946.755 101.185 946.880 ;
        RECT 6.290 942.685 1155.710 946.755 ;
        RECT 6.290 942.560 249.025 942.685 ;
      LAYER Pwell ;
        RECT 6.290 939.040 1155.710 942.560 ;
      LAYER Nwell ;
        RECT 6.290 938.915 287.105 939.040 ;
        RECT 6.290 934.845 1155.710 938.915 ;
        RECT 6.290 934.720 114.625 934.845 ;
      LAYER Pwell ;
        RECT 6.290 931.200 1155.710 934.720 ;
      LAYER Nwell ;
        RECT 6.290 931.075 218.785 931.200 ;
        RECT 6.290 927.005 1155.710 931.075 ;
        RECT 6.290 926.880 241.960 927.005 ;
      LAYER Pwell ;
        RECT 6.290 923.360 1155.710 926.880 ;
      LAYER Nwell ;
        RECT 6.290 923.235 257.640 923.360 ;
        RECT 6.290 919.165 1155.710 923.235 ;
        RECT 6.290 919.040 193.585 919.165 ;
      LAYER Pwell ;
        RECT 6.290 915.520 1155.710 919.040 ;
      LAYER Nwell ;
        RECT 6.290 915.395 296.625 915.520 ;
        RECT 6.290 911.325 1155.710 915.395 ;
        RECT 6.290 911.200 210.945 911.325 ;
      LAYER Pwell ;
        RECT 6.290 907.680 1155.710 911.200 ;
      LAYER Nwell ;
        RECT 6.290 907.555 370.125 907.680 ;
        RECT 6.290 903.485 1155.710 907.555 ;
        RECT 6.290 903.360 189.105 903.485 ;
      LAYER Pwell ;
        RECT 6.290 899.840 1155.710 903.360 ;
      LAYER Nwell ;
        RECT 6.290 899.715 261.905 899.840 ;
        RECT 6.290 895.645 1155.710 899.715 ;
        RECT 6.290 895.520 369.565 895.645 ;
      LAYER Pwell ;
        RECT 6.290 892.000 1155.710 895.520 ;
      LAYER Nwell ;
        RECT 6.290 891.875 210.945 892.000 ;
        RECT 6.290 887.805 1155.710 891.875 ;
        RECT 6.290 887.680 195.265 887.805 ;
      LAYER Pwell ;
        RECT 6.290 884.160 1155.710 887.680 ;
      LAYER Nwell ;
        RECT 6.290 884.035 180.360 884.160 ;
        RECT 6.290 879.965 1155.710 884.035 ;
        RECT 6.290 879.840 319.585 879.965 ;
      LAYER Pwell ;
        RECT 6.290 876.320 1155.710 879.840 ;
      LAYER Nwell ;
        RECT 6.290 876.195 226.280 876.320 ;
        RECT 6.290 872.125 1155.710 876.195 ;
        RECT 6.290 872.000 243.080 872.125 ;
      LAYER Pwell ;
        RECT 6.290 868.480 1155.710 872.000 ;
      LAYER Nwell ;
        RECT 6.290 868.355 177.345 868.480 ;
        RECT 6.290 864.285 1155.710 868.355 ;
        RECT 6.290 864.160 199.745 864.285 ;
      LAYER Pwell ;
        RECT 6.290 860.640 1155.710 864.160 ;
      LAYER Nwell ;
        RECT 6.290 860.515 176.225 860.640 ;
        RECT 6.290 856.445 1155.710 860.515 ;
        RECT 6.290 856.320 241.745 856.445 ;
      LAYER Pwell ;
        RECT 6.290 852.800 1155.710 856.320 ;
      LAYER Nwell ;
        RECT 6.290 852.675 228.520 852.800 ;
        RECT 6.290 848.605 1155.710 852.675 ;
        RECT 6.290 848.480 276.465 848.605 ;
      LAYER Pwell ;
        RECT 6.290 844.960 1155.710 848.480 ;
      LAYER Nwell ;
        RECT 6.290 844.835 178.465 844.960 ;
        RECT 6.290 840.765 1155.710 844.835 ;
        RECT 6.290 840.640 168.600 840.765 ;
      LAYER Pwell ;
        RECT 6.290 837.120 1155.710 840.640 ;
      LAYER Nwell ;
        RECT 6.290 836.995 235.800 837.120 ;
        RECT 6.290 832.925 1155.710 836.995 ;
        RECT 6.290 832.800 199.185 832.925 ;
      LAYER Pwell ;
        RECT 6.290 829.280 1155.710 832.800 ;
      LAYER Nwell ;
        RECT 6.290 829.155 218.225 829.280 ;
        RECT 6.290 825.085 1155.710 829.155 ;
        RECT 6.290 824.960 201.005 825.085 ;
      LAYER Pwell ;
        RECT 6.290 821.440 1155.710 824.960 ;
      LAYER Nwell ;
        RECT 6.290 821.315 152.145 821.440 ;
        RECT 6.290 817.245 1155.710 821.315 ;
        RECT 6.290 817.120 255.400 817.245 ;
      LAYER Pwell ;
        RECT 6.290 813.600 1155.710 817.120 ;
      LAYER Nwell ;
        RECT 6.290 813.475 193.725 813.600 ;
        RECT 6.290 809.405 1155.710 813.475 ;
        RECT 6.290 809.280 201.005 809.405 ;
      LAYER Pwell ;
        RECT 6.290 805.760 1155.710 809.280 ;
      LAYER Nwell ;
        RECT 6.290 805.635 98.945 805.760 ;
        RECT 6.290 801.565 1155.710 805.635 ;
        RECT 6.290 801.440 523.640 801.565 ;
      LAYER Pwell ;
        RECT 6.290 797.920 1155.710 801.440 ;
      LAYER Nwell ;
        RECT 6.290 797.795 218.415 797.920 ;
        RECT 6.290 793.725 1155.710 797.795 ;
        RECT 6.290 793.600 117.425 793.725 ;
      LAYER Pwell ;
        RECT 6.290 790.080 1155.710 793.600 ;
      LAYER Nwell ;
        RECT 6.290 789.955 96.145 790.080 ;
        RECT 6.290 785.885 1155.710 789.955 ;
        RECT 6.290 785.760 247.485 785.885 ;
      LAYER Pwell ;
        RECT 6.290 782.240 1155.710 785.760 ;
      LAYER Nwell ;
        RECT 6.290 782.115 268.625 782.240 ;
        RECT 6.290 778.045 1155.710 782.115 ;
        RECT 6.290 777.920 72.625 778.045 ;
      LAYER Pwell ;
        RECT 6.290 774.400 1155.710 777.920 ;
      LAYER Nwell ;
        RECT 6.290 774.275 169.505 774.400 ;
        RECT 6.290 770.205 1155.710 774.275 ;
        RECT 6.290 770.080 92.785 770.205 ;
      LAYER Pwell ;
        RECT 6.290 766.560 1155.710 770.080 ;
      LAYER Nwell ;
        RECT 6.290 766.435 68.705 766.560 ;
        RECT 6.290 762.365 1155.710 766.435 ;
        RECT 6.290 762.240 44.625 762.365 ;
      LAYER Pwell ;
        RECT 6.290 758.720 1155.710 762.240 ;
      LAYER Nwell ;
        RECT 6.290 758.595 411.985 758.720 ;
        RECT 6.290 754.525 1155.710 758.595 ;
        RECT 6.290 754.400 149.905 754.525 ;
      LAYER Pwell ;
        RECT 6.290 750.880 1155.710 754.400 ;
      LAYER Nwell ;
        RECT 6.290 750.755 24.465 750.880 ;
        RECT 6.290 746.685 1155.710 750.755 ;
        RECT 6.290 746.560 345.905 746.685 ;
      LAYER Pwell ;
        RECT 6.290 743.040 1155.710 746.560 ;
      LAYER Nwell ;
        RECT 6.290 742.915 179.800 743.040 ;
        RECT 6.290 738.845 1155.710 742.915 ;
        RECT 6.290 738.720 12.705 738.845 ;
      LAYER Pwell ;
        RECT 6.290 735.200 1155.710 738.720 ;
      LAYER Nwell ;
        RECT 6.290 735.075 98.385 735.200 ;
        RECT 6.290 731.005 1155.710 735.075 ;
        RECT 6.290 730.880 310.220 731.005 ;
      LAYER Pwell ;
        RECT 6.290 727.360 1155.710 730.880 ;
      LAYER Nwell ;
        RECT 6.290 727.235 348.920 727.360 ;
        RECT 6.290 723.165 1155.710 727.235 ;
        RECT 6.290 723.040 12.705 723.165 ;
      LAYER Pwell ;
        RECT 6.290 719.520 1155.710 723.040 ;
      LAYER Nwell ;
        RECT 6.290 719.395 107.905 719.520 ;
        RECT 6.290 715.325 1155.710 719.395 ;
        RECT 6.290 715.200 162.225 715.325 ;
      LAYER Pwell ;
        RECT 6.290 711.680 1155.710 715.200 ;
      LAYER Nwell ;
        RECT 6.290 711.555 265.825 711.680 ;
        RECT 6.290 707.485 1155.710 711.555 ;
        RECT 6.290 707.360 12.705 707.485 ;
      LAYER Pwell ;
        RECT 6.290 703.840 1155.710 707.360 ;
      LAYER Nwell ;
        RECT 6.290 703.715 64.785 703.840 ;
        RECT 6.290 699.645 1155.710 703.715 ;
        RECT 6.290 699.520 233.905 699.645 ;
      LAYER Pwell ;
        RECT 6.290 696.000 1155.710 699.520 ;
      LAYER Nwell ;
        RECT 6.290 695.875 223.480 696.000 ;
        RECT 6.290 691.805 1155.710 695.875 ;
        RECT 6.290 691.680 12.705 691.805 ;
      LAYER Pwell ;
        RECT 6.290 688.160 1155.710 691.680 ;
      LAYER Nwell ;
        RECT 6.290 688.035 184.625 688.160 ;
        RECT 6.290 683.965 1155.710 688.035 ;
        RECT 6.290 683.840 90.545 683.965 ;
      LAYER Pwell ;
        RECT 6.290 680.320 1155.710 683.840 ;
      LAYER Nwell ;
        RECT 6.290 680.195 54.145 680.320 ;
        RECT 6.290 676.125 1155.710 680.195 ;
        RECT 6.290 676.000 12.705 676.125 ;
      LAYER Pwell ;
        RECT 6.290 672.480 1155.710 676.000 ;
      LAYER Nwell ;
        RECT 6.290 672.355 31.745 672.480 ;
        RECT 6.290 668.285 1155.710 672.355 ;
        RECT 6.290 668.160 54.145 668.285 ;
      LAYER Pwell ;
        RECT 6.290 664.640 1155.710 668.160 ;
      LAYER Nwell ;
        RECT 6.290 664.515 100.625 664.640 ;
        RECT 6.290 660.445 1155.710 664.515 ;
        RECT 6.290 660.320 12.705 660.445 ;
      LAYER Pwell ;
        RECT 6.290 656.800 1155.710 660.320 ;
      LAYER Nwell ;
        RECT 6.290 656.675 184.130 656.800 ;
        RECT 6.290 652.605 1155.710 656.675 ;
        RECT 6.290 652.480 39.025 652.605 ;
      LAYER Pwell ;
        RECT 6.290 648.960 1155.710 652.480 ;
      LAYER Nwell ;
        RECT 6.290 648.835 100.625 648.960 ;
        RECT 6.290 644.765 1155.710 648.835 ;
        RECT 6.290 644.640 12.705 644.765 ;
      LAYER Pwell ;
        RECT 6.290 641.120 1155.710 644.640 ;
      LAYER Nwell ;
        RECT 6.290 640.995 28.385 641.120 ;
        RECT 6.290 636.925 1155.710 640.995 ;
        RECT 6.290 636.800 50.225 636.925 ;
      LAYER Pwell ;
        RECT 6.290 633.280 1155.710 636.800 ;
      LAYER Nwell ;
        RECT 6.290 633.155 66.465 633.280 ;
        RECT 6.290 629.085 1155.710 633.155 ;
        RECT 6.290 628.960 12.705 629.085 ;
      LAYER Pwell ;
        RECT 6.290 625.440 1155.710 628.960 ;
      LAYER Nwell ;
        RECT 6.290 625.315 32.865 625.440 ;
        RECT 6.290 621.245 1155.710 625.315 ;
        RECT 6.290 621.120 194.330 621.245 ;
      LAYER Pwell ;
        RECT 6.290 617.600 1155.710 621.120 ;
      LAYER Nwell ;
        RECT 6.290 617.475 52.655 617.600 ;
        RECT 6.290 613.405 1155.710 617.475 ;
        RECT 6.290 613.280 12.705 613.405 ;
      LAYER Pwell ;
        RECT 6.290 609.760 1155.710 613.280 ;
      LAYER Nwell ;
        RECT 6.290 609.635 50.975 609.760 ;
        RECT 6.290 605.565 1155.710 609.635 ;
        RECT 6.290 605.440 40.360 605.565 ;
      LAYER Pwell ;
        RECT 6.290 601.920 1155.710 605.440 ;
      LAYER Nwell ;
        RECT 6.290 601.795 99.505 601.920 ;
        RECT 6.290 597.725 1155.710 601.795 ;
        RECT 6.290 597.600 12.705 597.725 ;
      LAYER Pwell ;
        RECT 6.290 594.080 1155.710 597.600 ;
      LAYER Nwell ;
        RECT 6.290 593.955 60.865 594.080 ;
        RECT 6.290 589.885 1155.710 593.955 ;
        RECT 6.290 589.760 129.185 589.885 ;
      LAYER Pwell ;
        RECT 6.290 586.240 1155.710 589.760 ;
      LAYER Nwell ;
        RECT 6.290 586.115 12.705 586.240 ;
        RECT 6.290 582.045 1155.710 586.115 ;
        RECT 6.290 581.920 345.905 582.045 ;
      LAYER Pwell ;
        RECT 6.290 578.400 1155.710 581.920 ;
      LAYER Nwell ;
        RECT 6.290 578.275 62.545 578.400 ;
        RECT 6.290 574.205 1155.710 578.275 ;
        RECT 6.290 574.080 282.065 574.205 ;
      LAYER Pwell ;
        RECT 6.290 570.560 1155.710 574.080 ;
      LAYER Nwell ;
        RECT 6.290 570.435 12.705 570.560 ;
        RECT 6.290 566.365 1155.710 570.435 ;
        RECT 6.290 566.240 53.800 566.365 ;
      LAYER Pwell ;
        RECT 6.290 562.720 1155.710 566.240 ;
      LAYER Nwell ;
        RECT 6.290 562.595 64.785 562.720 ;
        RECT 6.290 558.525 1155.710 562.595 ;
        RECT 6.290 558.400 82.145 558.525 ;
      LAYER Pwell ;
        RECT 6.290 554.880 1155.710 558.400 ;
      LAYER Nwell ;
        RECT 6.290 554.755 27.265 554.880 ;
        RECT 6.290 550.685 1155.710 554.755 ;
        RECT 6.290 550.560 12.705 550.685 ;
      LAYER Pwell ;
        RECT 6.290 547.040 1155.710 550.560 ;
      LAYER Nwell ;
        RECT 6.290 546.915 64.225 547.040 ;
        RECT 6.290 542.845 1155.710 546.915 ;
        RECT 6.290 542.720 95.715 542.845 ;
      LAYER Pwell ;
        RECT 6.290 539.200 1155.710 542.720 ;
      LAYER Nwell ;
        RECT 6.290 539.075 215.640 539.200 ;
        RECT 6.290 535.005 1155.710 539.075 ;
        RECT 6.290 534.880 12.705 535.005 ;
      LAYER Pwell ;
        RECT 6.290 531.360 1155.710 534.880 ;
      LAYER Nwell ;
        RECT 6.290 531.235 53.025 531.360 ;
        RECT 6.290 527.165 1155.710 531.235 ;
        RECT 6.290 527.040 75.555 527.165 ;
      LAYER Pwell ;
        RECT 6.290 523.520 1155.710 527.040 ;
      LAYER Nwell ;
        RECT 6.290 523.395 34.545 523.520 ;
        RECT 6.290 519.325 1155.710 523.395 ;
        RECT 6.290 519.200 12.705 519.325 ;
      LAYER Pwell ;
        RECT 6.290 515.680 1155.710 519.200 ;
      LAYER Nwell ;
        RECT 6.290 515.555 287.105 515.680 ;
        RECT 6.290 511.485 1155.710 515.555 ;
        RECT 6.290 511.360 71.505 511.485 ;
      LAYER Pwell ;
        RECT 6.290 507.840 1155.710 511.360 ;
      LAYER Nwell ;
        RECT 6.290 507.715 34.545 507.840 ;
        RECT 6.290 503.645 1155.710 507.715 ;
        RECT 6.290 503.520 150.465 503.645 ;
      LAYER Pwell ;
        RECT 6.290 500.000 1155.710 503.520 ;
      LAYER Nwell ;
        RECT 6.290 499.875 12.705 500.000 ;
        RECT 6.290 495.805 1155.710 499.875 ;
        RECT 6.290 495.680 404.370 495.805 ;
      LAYER Pwell ;
        RECT 6.290 492.160 1155.710 495.680 ;
      LAYER Nwell ;
        RECT 6.290 492.035 54.145 492.160 ;
        RECT 6.290 487.965 1155.710 492.035 ;
        RECT 6.290 487.840 35.105 487.965 ;
      LAYER Pwell ;
        RECT 6.290 484.320 1155.710 487.840 ;
      LAYER Nwell ;
        RECT 6.290 484.195 12.705 484.320 ;
        RECT 6.290 480.125 1155.710 484.195 ;
        RECT 6.290 480.000 131.985 480.125 ;
      LAYER Pwell ;
        RECT 6.290 476.480 1155.710 480.000 ;
      LAYER Nwell ;
        RECT 6.290 476.355 63.105 476.480 ;
        RECT 6.290 472.285 1155.710 476.355 ;
        RECT 6.290 472.160 45.745 472.285 ;
      LAYER Pwell ;
        RECT 6.290 468.640 1155.710 472.160 ;
      LAYER Nwell ;
        RECT 6.290 468.515 24.465 468.640 ;
        RECT 6.290 464.445 1155.710 468.515 ;
        RECT 6.290 464.320 128.065 464.445 ;
      LAYER Pwell ;
        RECT 6.290 460.800 1155.710 464.320 ;
      LAYER Nwell ;
        RECT 6.290 460.675 62.545 460.800 ;
        RECT 6.290 456.605 1155.710 460.675 ;
        RECT 6.290 456.480 33.425 456.605 ;
      LAYER Pwell ;
        RECT 6.290 452.960 1155.710 456.480 ;
      LAYER Nwell ;
        RECT 6.290 452.835 14.385 452.960 ;
        RECT 6.290 448.765 1155.710 452.835 ;
        RECT 6.290 448.640 79.905 448.765 ;
      LAYER Pwell ;
        RECT 6.290 445.120 1155.710 448.640 ;
      LAYER Nwell ;
        RECT 6.290 444.995 51.905 445.120 ;
        RECT 6.290 440.925 1155.710 444.995 ;
        RECT 6.290 440.800 32.305 440.925 ;
      LAYER Pwell ;
        RECT 6.290 437.280 1155.710 440.800 ;
      LAYER Nwell ;
        RECT 6.290 437.155 171.185 437.280 ;
        RECT 6.290 433.085 1155.710 437.155 ;
        RECT 6.290 432.960 570.505 433.085 ;
      LAYER Pwell ;
        RECT 6.290 429.440 1155.710 432.960 ;
      LAYER Nwell ;
        RECT 6.290 429.315 12.705 429.440 ;
        RECT 6.290 425.245 1155.710 429.315 ;
        RECT 6.290 425.120 308.385 425.245 ;
      LAYER Pwell ;
        RECT 6.290 421.600 1155.710 425.120 ;
      LAYER Nwell ;
        RECT 6.290 421.475 31.185 421.600 ;
        RECT 6.290 417.405 1155.710 421.475 ;
        RECT 6.290 417.280 71.505 417.405 ;
      LAYER Pwell ;
        RECT 6.290 413.760 1155.710 417.280 ;
      LAYER Nwell ;
        RECT 6.290 413.635 12.705 413.760 ;
        RECT 6.290 409.565 1155.710 413.635 ;
        RECT 6.290 409.440 56.600 409.565 ;
      LAYER Pwell ;
        RECT 6.290 405.920 1155.710 409.440 ;
      LAYER Nwell ;
        RECT 6.290 405.795 247.905 405.920 ;
        RECT 6.290 401.725 1155.710 405.795 ;
        RECT 6.290 401.600 71.505 401.725 ;
      LAYER Pwell ;
        RECT 6.290 398.080 1155.710 401.600 ;
      LAYER Nwell ;
        RECT 6.290 397.955 26.145 398.080 ;
        RECT 6.290 393.885 1155.710 397.955 ;
        RECT 6.290 393.760 308.945 393.885 ;
      LAYER Pwell ;
        RECT 6.290 390.240 1155.710 393.760 ;
      LAYER Nwell ;
        RECT 6.290 390.115 371.665 390.240 ;
        RECT 6.290 386.045 1155.710 390.115 ;
        RECT 6.290 385.920 45.185 386.045 ;
      LAYER Pwell ;
        RECT 6.290 382.400 1155.710 385.920 ;
      LAYER Nwell ;
        RECT 6.290 382.275 23.905 382.400 ;
        RECT 6.290 378.205 1155.710 382.275 ;
        RECT 6.290 378.080 201.640 378.205 ;
      LAYER Pwell ;
        RECT 6.290 374.560 1155.710 378.080 ;
      LAYER Nwell ;
        RECT 6.290 374.435 33.425 374.560 ;
        RECT 6.290 370.365 1155.710 374.435 ;
        RECT 6.290 370.240 51.905 370.365 ;
      LAYER Pwell ;
        RECT 6.290 366.720 1155.710 370.240 ;
      LAYER Nwell ;
        RECT 6.290 366.595 69.825 366.720 ;
        RECT 6.290 362.525 1155.710 366.595 ;
        RECT 6.290 362.400 388.465 362.525 ;
      LAYER Pwell ;
        RECT 6.290 358.880 1155.710 362.400 ;
      LAYER Nwell ;
        RECT 6.290 358.755 51.905 358.880 ;
        RECT 6.290 354.685 1155.710 358.755 ;
        RECT 6.290 354.560 127.505 354.685 ;
      LAYER Pwell ;
        RECT 6.290 351.040 1155.710 354.560 ;
      LAYER Nwell ;
        RECT 6.290 350.915 223.825 351.040 ;
        RECT 6.290 346.845 1155.710 350.915 ;
        RECT 6.290 346.720 72.625 346.845 ;
      LAYER Pwell ;
        RECT 6.290 343.200 1155.710 346.720 ;
      LAYER Nwell ;
        RECT 6.290 343.075 502.705 343.200 ;
        RECT 6.290 339.005 1155.710 343.075 ;
        RECT 6.290 338.880 49.665 339.005 ;
      LAYER Pwell ;
        RECT 6.290 335.360 1155.710 338.880 ;
      LAYER Nwell ;
        RECT 6.290 335.235 146.545 335.360 ;
        RECT 6.290 331.165 1155.710 335.235 ;
        RECT 6.290 331.040 77.665 331.165 ;
      LAYER Pwell ;
        RECT 6.290 327.520 1155.710 331.040 ;
      LAYER Nwell ;
        RECT 6.290 327.395 105.105 327.520 ;
        RECT 6.290 323.325 1155.710 327.395 ;
        RECT 6.290 323.200 50.225 323.325 ;
      LAYER Pwell ;
        RECT 6.290 319.680 1155.710 323.200 ;
      LAYER Nwell ;
        RECT 6.290 319.555 173.985 319.680 ;
        RECT 6.290 315.485 1155.710 319.555 ;
        RECT 6.290 315.360 130.305 315.485 ;
      LAYER Pwell ;
        RECT 6.290 311.840 1155.710 315.360 ;
      LAYER Nwell ;
        RECT 6.290 311.715 59.185 311.840 ;
        RECT 6.290 307.645 1155.710 311.715 ;
        RECT 6.290 307.520 437.185 307.645 ;
      LAYER Pwell ;
        RECT 6.290 304.000 1155.710 307.520 ;
      LAYER Nwell ;
        RECT 6.290 303.875 73.745 304.000 ;
        RECT 6.290 299.805 1155.710 303.875 ;
        RECT 6.290 299.680 128.065 299.805 ;
      LAYER Pwell ;
        RECT 6.290 296.160 1155.710 299.680 ;
      LAYER Nwell ;
        RECT 6.290 296.035 208.705 296.160 ;
        RECT 6.290 291.965 1155.710 296.035 ;
        RECT 6.290 291.840 110.705 291.965 ;
      LAYER Pwell ;
        RECT 6.290 288.320 1155.710 291.840 ;
      LAYER Nwell ;
        RECT 6.290 288.195 73.185 288.320 ;
        RECT 6.290 284.125 1155.710 288.195 ;
        RECT 6.290 284.000 162.785 284.125 ;
      LAYER Pwell ;
        RECT 6.290 280.480 1155.710 284.000 ;
      LAYER Nwell ;
        RECT 6.290 280.355 137.025 280.480 ;
        RECT 6.290 276.285 1155.710 280.355 ;
        RECT 6.290 276.160 98.600 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 1155.710 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 73.745 272.640 ;
        RECT 6.290 268.445 1155.710 272.515 ;
        RECT 6.290 268.320 189.105 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 1155.710 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 140.945 264.800 ;
        RECT 6.290 260.605 1155.710 264.675 ;
        RECT 6.290 260.480 121.905 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 1155.710 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 339.185 256.960 ;
        RECT 6.290 252.765 1155.710 256.835 ;
        RECT 6.290 252.640 90.200 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 1155.710 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 103.425 249.120 ;
        RECT 6.290 244.925 1155.710 248.995 ;
        RECT 6.290 244.800 123.585 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 1155.710 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 185.400 241.280 ;
        RECT 6.290 237.085 1155.710 241.155 ;
        RECT 6.290 236.960 95.240 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 1155.710 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 144.305 233.440 ;
        RECT 6.290 229.245 1155.710 233.315 ;
        RECT 6.290 229.120 168.040 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 1155.710 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 253.160 225.600 ;
        RECT 6.290 221.405 1155.710 225.475 ;
        RECT 6.290 221.280 405.965 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 1155.710 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 345.475 217.760 ;
        RECT 6.290 213.565 1155.710 217.635 ;
        RECT 6.290 213.440 165.025 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 1155.710 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 213.185 209.920 ;
        RECT 6.290 205.725 1155.710 209.795 ;
        RECT 6.290 205.600 476.600 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 1155.710 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 326.305 202.080 ;
        RECT 6.290 197.885 1155.710 201.955 ;
        RECT 6.290 197.760 163.905 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 1155.710 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 196.600 194.240 ;
        RECT 6.290 190.045 1155.710 194.115 ;
        RECT 6.290 189.920 361.240 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 1155.710 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 299.985 186.400 ;
        RECT 6.290 182.205 1155.710 186.275 ;
        RECT 6.290 182.080 171.745 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 1155.710 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 191.345 178.560 ;
        RECT 6.290 174.365 1155.710 178.435 ;
        RECT 6.290 174.240 238.385 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 1155.710 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 544.145 170.720 ;
        RECT 6.290 166.525 1155.710 170.595 ;
        RECT 6.290 166.400 390.360 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 1155.710 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 260.225 162.880 ;
        RECT 6.290 158.685 1155.710 162.755 ;
        RECT 6.290 158.560 189.665 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 1155.710 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 227.960 155.040 ;
        RECT 6.290 150.845 1155.710 154.915 ;
        RECT 6.290 150.720 328.545 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 1155.710 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 496.545 147.200 ;
        RECT 6.290 143.005 1155.710 147.075 ;
        RECT 6.290 142.880 204.225 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 1155.710 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 221.585 139.360 ;
        RECT 6.290 135.165 1155.710 139.235 ;
        RECT 6.290 135.040 238.385 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 1155.710 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 334.145 131.520 ;
        RECT 6.290 127.325 1155.710 131.395 ;
        RECT 6.290 127.200 278.285 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 1155.710 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 210.945 123.680 ;
        RECT 6.290 119.485 1155.710 123.555 ;
        RECT 6.290 119.360 238.385 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 1155.710 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 292.705 115.840 ;
        RECT 6.290 111.645 1155.710 115.715 ;
        RECT 6.290 111.520 228.305 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 1155.710 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 260.225 108.000 ;
        RECT 6.290 103.805 1155.710 107.875 ;
        RECT 6.290 103.680 242.865 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 1155.710 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 541.000 100.160 ;
        RECT 6.290 95.965 1155.710 100.035 ;
        RECT 6.290 95.840 326.305 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 1155.710 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 267.505 92.320 ;
        RECT 6.290 88.125 1155.710 92.195 ;
        RECT 6.290 88.000 446.145 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 1155.710 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 685.825 84.480 ;
        RECT 6.290 80.285 1155.710 84.355 ;
        RECT 6.290 80.160 426.545 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 1155.710 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 339.745 76.640 ;
        RECT 6.290 72.445 1155.710 76.515 ;
        RECT 6.290 72.320 357.105 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 1155.710 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 428.925 68.800 ;
        RECT 6.290 64.605 1155.710 68.675 ;
        RECT 6.290 64.480 709.500 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 1155.710 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 379.505 60.960 ;
        RECT 6.290 56.765 1155.710 60.835 ;
        RECT 6.290 56.640 360.465 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 1155.710 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 414.785 53.120 ;
        RECT 6.290 48.925 1155.710 52.995 ;
        RECT 6.290 48.800 489.480 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 1155.710 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 570.465 45.280 ;
        RECT 6.290 41.085 1155.710 45.155 ;
        RECT 6.290 40.960 364.945 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 1155.710 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 457.345 37.440 ;
        RECT 6.290 33.245 1155.710 37.315 ;
        RECT 6.290 33.120 424.305 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 1155.710 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 809.240 29.600 ;
        RECT 6.290 25.405 1155.710 29.475 ;
        RECT 6.290 25.280 435.160 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 1155.710 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 410.305 21.760 ;
        RECT 6.290 17.565 1155.710 21.635 ;
        RECT 6.290 17.440 775.985 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 1155.710 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 1155.280 1167.450 ;
      LAYER Metal2 ;
        RECT 7.980 1175.940 31.060 1176.980 ;
        RECT 32.220 1175.940 64.660 1176.980 ;
        RECT 65.820 1175.940 75.860 1176.980 ;
        RECT 77.020 1175.940 87.060 1176.980 ;
        RECT 88.220 1175.940 98.260 1176.980 ;
        RECT 99.420 1175.940 109.460 1176.980 ;
        RECT 110.620 1175.940 120.660 1176.980 ;
        RECT 121.820 1175.940 131.860 1176.980 ;
        RECT 133.020 1175.940 143.060 1176.980 ;
        RECT 144.220 1175.940 154.260 1176.980 ;
        RECT 155.420 1175.940 165.460 1176.980 ;
        RECT 166.620 1175.940 176.660 1176.980 ;
        RECT 177.820 1175.940 187.860 1176.980 ;
        RECT 189.020 1175.940 199.060 1176.980 ;
        RECT 200.220 1175.940 210.260 1176.980 ;
        RECT 211.420 1175.940 221.460 1176.980 ;
        RECT 222.620 1175.940 232.660 1176.980 ;
        RECT 233.820 1175.940 243.860 1176.980 ;
        RECT 245.020 1175.940 255.060 1176.980 ;
        RECT 256.220 1175.940 266.260 1176.980 ;
        RECT 267.420 1175.940 277.460 1176.980 ;
        RECT 278.620 1175.940 288.660 1176.980 ;
        RECT 289.820 1175.940 299.860 1176.980 ;
        RECT 301.020 1175.940 311.060 1176.980 ;
        RECT 312.220 1175.940 322.260 1176.980 ;
        RECT 323.420 1175.940 333.460 1176.980 ;
        RECT 334.620 1175.940 344.660 1176.980 ;
        RECT 345.820 1175.940 355.860 1176.980 ;
        RECT 357.020 1175.940 367.060 1176.980 ;
        RECT 368.220 1175.940 378.260 1176.980 ;
        RECT 379.420 1175.940 389.460 1176.980 ;
        RECT 390.620 1175.940 400.660 1176.980 ;
        RECT 401.820 1175.940 411.860 1176.980 ;
        RECT 413.020 1175.940 423.060 1176.980 ;
        RECT 424.220 1175.940 434.260 1176.980 ;
        RECT 435.420 1175.940 445.460 1176.980 ;
        RECT 446.620 1175.940 456.660 1176.980 ;
        RECT 457.820 1175.940 467.860 1176.980 ;
        RECT 469.020 1175.940 479.060 1176.980 ;
        RECT 480.220 1175.940 490.260 1176.980 ;
        RECT 491.420 1175.940 501.460 1176.980 ;
        RECT 502.620 1175.940 512.660 1176.980 ;
        RECT 513.820 1175.940 523.860 1176.980 ;
        RECT 525.020 1175.940 535.060 1176.980 ;
        RECT 536.220 1175.940 546.260 1176.980 ;
        RECT 547.420 1175.940 557.460 1176.980 ;
        RECT 558.620 1175.940 568.660 1176.980 ;
        RECT 569.820 1175.940 579.860 1176.980 ;
        RECT 581.020 1175.940 591.060 1176.980 ;
        RECT 592.220 1175.940 602.260 1176.980 ;
        RECT 603.420 1175.940 613.460 1176.980 ;
        RECT 614.620 1175.940 624.660 1176.980 ;
        RECT 625.820 1175.940 635.860 1176.980 ;
        RECT 637.020 1175.940 647.060 1176.980 ;
        RECT 648.220 1175.940 658.260 1176.980 ;
        RECT 659.420 1175.940 669.460 1176.980 ;
        RECT 670.620 1175.940 680.660 1176.980 ;
        RECT 681.820 1175.940 691.860 1176.980 ;
        RECT 693.020 1175.940 703.060 1176.980 ;
        RECT 704.220 1175.940 714.260 1176.980 ;
        RECT 715.420 1175.940 725.460 1176.980 ;
        RECT 726.620 1175.940 736.660 1176.980 ;
        RECT 737.820 1175.940 747.860 1176.980 ;
        RECT 749.020 1175.940 759.060 1176.980 ;
        RECT 760.220 1175.940 770.260 1176.980 ;
        RECT 771.420 1175.940 781.460 1176.980 ;
        RECT 782.620 1175.940 792.660 1176.980 ;
        RECT 793.820 1175.940 803.860 1176.980 ;
        RECT 805.020 1175.940 815.060 1176.980 ;
        RECT 816.220 1175.940 826.260 1176.980 ;
        RECT 827.420 1175.940 837.460 1176.980 ;
        RECT 838.620 1175.940 848.660 1176.980 ;
        RECT 849.820 1175.940 859.860 1176.980 ;
        RECT 861.020 1175.940 871.060 1176.980 ;
        RECT 872.220 1175.940 882.260 1176.980 ;
        RECT 883.420 1175.940 893.460 1176.980 ;
        RECT 894.620 1175.940 904.660 1176.980 ;
        RECT 905.820 1175.940 915.860 1176.980 ;
        RECT 917.020 1175.940 927.060 1176.980 ;
        RECT 928.220 1175.940 938.260 1176.980 ;
        RECT 939.420 1175.940 949.460 1176.980 ;
        RECT 950.620 1175.940 960.660 1176.980 ;
        RECT 961.820 1175.940 971.860 1176.980 ;
        RECT 973.020 1175.940 983.060 1176.980 ;
        RECT 984.220 1175.940 994.260 1176.980 ;
        RECT 995.420 1175.940 1005.460 1176.980 ;
        RECT 1006.620 1175.940 1016.660 1176.980 ;
        RECT 1017.820 1175.940 1027.860 1176.980 ;
        RECT 1029.020 1175.940 1039.060 1176.980 ;
        RECT 1040.220 1175.940 1050.260 1176.980 ;
        RECT 1051.420 1175.940 1061.460 1176.980 ;
        RECT 1062.620 1175.940 1072.660 1176.980 ;
        RECT 1073.820 1175.940 1083.860 1176.980 ;
        RECT 1085.020 1175.940 1095.060 1176.980 ;
        RECT 1096.220 1175.940 1106.260 1176.980 ;
        RECT 1107.420 1175.940 1117.460 1176.980 ;
        RECT 1118.620 1175.940 1128.660 1176.980 ;
        RECT 1129.820 1175.940 1153.460 1176.980 ;
        RECT 7.980 4.010 1153.460 1175.940 ;
      LAYER Metal3 ;
        RECT 7.930 4.060 1153.510 1175.300 ;
      LAYER Metal4 ;
        RECT 121.100 1164.840 1128.820 1173.110 ;
        RECT 121.100 15.080 175.540 1164.840 ;
        RECT 177.740 15.080 252.340 1164.840 ;
        RECT 254.540 15.080 329.140 1164.840 ;
        RECT 331.340 15.080 405.940 1164.840 ;
        RECT 408.140 15.080 482.740 1164.840 ;
        RECT 484.940 15.080 559.540 1164.840 ;
        RECT 561.740 15.080 636.340 1164.840 ;
        RECT 638.540 15.080 713.140 1164.840 ;
        RECT 715.340 15.080 789.940 1164.840 ;
        RECT 792.140 15.080 866.740 1164.840 ;
        RECT 868.940 15.080 943.540 1164.840 ;
        RECT 945.740 15.080 1020.340 1164.840 ;
        RECT 1022.540 15.080 1097.140 1164.840 ;
        RECT 1099.340 15.080 1128.820 1164.840 ;
        RECT 121.100 4.570 1128.820 15.080 ;
  END
END user_proj_cpu
END LIBRARY

