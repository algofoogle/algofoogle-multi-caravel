* NGSPICE file created from top_raybox_zero_fsm.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_2 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

.subckt top_raybox_zero_fsm i_clk i_debug_map_overlay i_debug_trace_overlay i_debug_vec_overlay
+ i_gpout0_sel[0] i_gpout0_sel[1] i_gpout0_sel[2] i_gpout0_sel[3] i_gpout1_sel[0]
+ i_gpout1_sel[1] i_gpout1_sel[2] i_gpout1_sel[3] i_gpout2_sel[0] i_gpout2_sel[1]
+ i_gpout2_sel[2] i_gpout2_sel[3] i_mode[0] i_mode[1] i_mode[2] i_reg_csb i_reg_mosi
+ i_reg_outs_enb i_reg_sclk i_reset i_tex_in[0] i_tex_in[1] i_tex_in[2] i_tex_in[3]
+ i_vec_csb i_vec_mosi i_vec_sclk o_gpout[0] o_gpout[1] o_gpout[2] o_hsync o_rgb[0]
+ o_rgb[1] o_rgb[2] o_rgb[3] o_rgb[4] o_rgb[5] o_tex_csb o_tex_oeb0 o_tex_out0 o_tex_sclk
+ o_vsync vdd vss
XFILLER_0_185_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18869_ _11787_ _11788_ _11789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_222_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20900_ _01914_ _01989_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_21880_ _02905_ _02919_ _02922_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20831_ _12841_ _01920_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_210_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_176_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23550_ _03713_ _04150_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20762_ _01810_ _01812_ _01852_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__20353__A1 _12955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22501_ _03422_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_23481_ _04320_ _04334_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20693_ _01666_ _01771_ _01783_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19346__I0 rbzero.tex_b1\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21978__S _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_213_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25220_ _06003_ _06000_ _06004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_31_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22432_ _01892_ _03363_ _03375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_230_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25151_ _05933_ _05934_ _05935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__20656__A2 _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22363_ _03306_ _03311_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25249__I _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24102_ _04809_ _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_21314_ _02225_ _02239_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25082_ _05825_ _05826_ _05865_ _05866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_143_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14335__A2 _08022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22294_ _11179_ _03254_ _03255_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24033_ net46 _04814_ _04815_ _04816_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_103_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21245_ _02187_ _02202_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_102_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14612__C _07604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_228_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21176_ _02256_ _02259_ _02263_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__13509__B gpout0.vinf vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20127_ _12893_ _12898_ _12899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_244_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25984_ _06686_ _06638_ _06762_ _06703_ _06763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__13228__C _07041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22030__A1 _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20058_ _12758_ _12829_ _12830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24935_ _05308_ _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_70_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22401__I _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_241_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22581__A2 _10072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24866_ _05644_ _05646_ _05649_ _05650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__20592__A1 _12403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24858__A1 _05640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26605_ _00515_ clknet_leaf_170_i_clk rbzero.tex_b0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_197_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23817_ _04646_ _04649_ _04650_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_213_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24797_ _05526_ _05580_ _05581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15015__I _08813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14059__C _07868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14550_ _07665_ _08358_ _08359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26536_ _00446_ clknet_leaf_22_i_clk rbzero.pov.spi_buffer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23748_ rbzero.wall_tracer.trackDistY\[-3\] _03053_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13501_ _07272_ _07276_ _07311_ _07312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_82_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14481_ rbzero.tex_g0\[33\] _08288_ _08289_ _08290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14023__A1 rbzero.tex_r1\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26467_ _00377_ clknet_leaf_44_i_clk rbzero.debug_overlay.playerY\[-7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23679_ _02750_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_165_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16220_ rbzero.spi_registers.buf_texadd1\[21\] _09730_ _09735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_101_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17760__A2 rbzero.pov.ready_buffer\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25418_ _06031_ _06102_ _06202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13432_ _07242_ _07243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_180_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26398_ _00308_ clknet_leaf_3_i_clk rbzero.spi_registers.buf_texadd2\[18\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_182_i_clk clknet_5_2__leaf_i_clk clknet_leaf_182_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_107_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16151_ _08922_ _09676_ _09684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25349_ _05982_ _06032_ _06133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_13363_ gpout0.vpos\[8\] _07175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xrebuffer7 _05577_ net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_248_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15102_ rbzero.spi_registers.spi_counter\[1\] _08891_ _08892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_107_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_248_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_248_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16082_ rbzero.spi_registers.buf_texadd0\[11\] _09622_ _09631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13294_ _07036_ _07108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_106_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19910_ _12677_ _12681_ _12682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_27019_ _00929_ clknet_leaf_169_i_clk rbzero.tex_g0\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_15033_ rbzero.spi_registers.spi_cmd\[1\] _08826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_239_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_197_i_clk clknet_5_12__leaf_i_clk clknet_leaf_197_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19841_ _12546_ _12566_ _12613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_236_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13419__B _07178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18996__I _11871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19772_ _12468_ _12485_ _12544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_219_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16984_ _10373_ _10391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_120_i_clk clknet_5_18__leaf_i_clk clknet_leaf_120_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_108_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22021__A1 rbzero.wall_tracer.stepDistY\[-10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15935_ _09517_ _09519_ _09520_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18723_ _11689_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_218_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_18654_ _11649_ _11650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15866_ _09467_ _09468_ _09448_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_88_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17605_ _10834_ _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14817_ _08622_ _08623_ _07149_ _07194_ _08624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_118_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18585_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _11608_ _11611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_135_i_clk clknet_5_15__leaf_i_clk clknet_leaf_135_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_204_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15797_ rbzero.spi_registers.buf_texadd3\[16\] _09409_ _09416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17536_ rbzero.tex_b0\[28\] rbzero.tex_b0\[27\] _10791_ _10795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14748_ rbzero.tex_b0\[27\] _08554_ _08459_ _08555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_clkbuf_leaf_148_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17467_ _10753_ _10746_ _10754_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14679_ rbzero.color_floor\[3\] _07966_ _07670_ _08486_ _08487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_104_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16418_ rbzero.spi_registers.buf_texadd3\[23\] _09874_ _09883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19206_ _12044_ _12049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17398_ _10702_ _10700_ _10703_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_171_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20638__A2 _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19137_ _11916_ _11980_ _11981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_15_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21835__A1 rbzero.debug_overlay.vplaneX\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16349_ _09806_ _09833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_119_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_200_i_clk_I clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19068_ _11912_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_18019_ rbzero.wall_tracer.trackDistX\[3\] _11163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_23_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21030_ _12705_ _01805_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15817__A2 _09032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14004__I _07501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16490__A2 _08099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22981_ _03683_ _03697_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24720_ _05327_ _05435_ _05436_ _05504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_21932_ _01662_ _02967_ _02970_ _02887_ _02971_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_179_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_20__f_i_clk clknet_3_5_0_i_clk clknet_5_20__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_24651_ _05286_ _05313_ _05332_ _05335_ _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_21863_ _11020_ _11072_ _08122_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_195_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23602_ _04402_ _04452_ _04453_ _04407_ _04400_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_27370_ _01275_ clknet_leaf_97_i_clk rbzero.wall_tracer.trackDistY\[-10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20814_ _01902_ _01903_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24582_ _05238_ _05305_ _05366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13999__B _07808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21794_ _10463_ _10448_ _02842_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26321_ _00231_ clknet_leaf_236_i_clk rbzero.spi_registers.buf_mapdx\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_212_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23533_ _04179_ _02293_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20745_ _12284_ _01729_ _01722_ _12264_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_147_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14005__B2 _07814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22079__A1 _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26252_ _00162_ clknet_leaf_2_i_clk rbzero.spi_registers.texadd2\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14607__C _07868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23464_ _04309_ _04317_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20676_ _01738_ _01767_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14556__A2 _08364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25203_ _05981_ _05984_ _05985_ _05987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22415_ _03351_ _03358_ _03359_ _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26183_ _00093_ clknet_leaf_235_i_clk rbzero.spi_registers.vshift\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_66_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23395_ _04247_ _04248_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25134_ _05331_ _05917_ _05888_ _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_189_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25568__A2 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22346_ _03296_ _03243_ _03297_ _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__22626__I0 rbzero.wall_tracer.texu\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25065_ _05411_ net91 _05849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22277_ _11191_ _03226_ _03240_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24016_ _04798_ _04800_ _08811_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_21228_ _02179_ _02289_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_236_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_243_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21159_ _02110_ _02123_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_208_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_208_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25967_ _06650_ _06640_ _06747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13981_ _07684_ _07219_ _07790_ _07791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14492__A1 rbzero.tex_g0\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_52_i_clk clknet_5_23__leaf_i_clk clknet_leaf_52_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15720_ rbzero.spi_registers.texadd2\[20\] _09350_ _09359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_198_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24918_ _05419_ _05695_ _05698_ _05699_ _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_25898_ _06672_ _06680_ _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_87_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15651_ rbzero.spi_registers.texadd2\[2\] _09303_ _09308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24849_ _05343_ _05490_ _05542_ _05633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_73_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19440__I _12211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22306__A2 _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14602_ _08406_ _08407_ _08409_ _07861_ _07638_ _08410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_18370_ _11488_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_201_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15582_ rbzero.spi_registers.texadd1\[9\] _09255_ _09256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_67_i_clk clknet_5_21__leaf_i_clk clknet_leaf_67_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17321_ _10611_ _10646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__20868__A2 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26519_ _00429_ clknet_leaf_57_i_clk rbzero.debug_overlay.vplaneY\[-3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14533_ _07459_ _08342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_141_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17252_ rbzero.pov.spi_buffer\[17\] _10591_ _10588_ _10595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14547__A2 _08354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14464_ _07574_ _08246_ _08256_ _08263_ _08272_ _08273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__23806__A2 _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16203_ _09711_ _09723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13415_ gpout0.vpos\[6\] _07226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_180_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17183_ _10541_ _10542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19486__A2 _12245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14395_ rbzero.tex_g0\[28\] _07461_ _08204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16134_ _08843_ _09669_ _09670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13346_ _07157_ net12 _07158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__22490__A1 rbzero.wall_tracer.size\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16065_ _08946_ _09612_ _09619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13277_ _06975_ _06944_ _06974_ _07091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_15016_ _08811_ _08814_ _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_224_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_114_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17844__B _10988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_74_i_clk_I clknet_5_29__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19824_ _12595_ _12199_ _12596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_166_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19755_ _12298_ _12527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16967_ _10377_ _10378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_34_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23742__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18706_ rbzero.tex_r1\[23\] rbzero.tex_r1\[22\] _11677_ _11680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_190_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15918_ _09507_ _09508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19686_ _12449_ _12457_ _12458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_79_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16898_ _10314_ _10315_ _10318_ _10319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_204_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20020__A3 _12789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18637_ _11640_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15849_ rbzero.spi_registers.buf_sky\[5\] _09438_ _09455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20308__A1 _12986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18568_ rbzero.tex_r0\[28\] rbzero.tex_r0\[27\] _11597_ _11601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15983__A1 _08973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17519_ _10785_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_138_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18499_ _11561_ _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20530_ _01610_ _01622_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_156_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14538__A2 _07901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20461_ _01455_ _01549_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24470__A2 _05205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22200_ _03108_ _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23180_ _03918_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__21284__A2 _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20392_ _12933_ _01383_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22131_ _03120_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16160__A1 _09542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19229__A2 _12051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_22062_ rbzero.wall_tracer.rcp_fsm.o_data\[3\] rbzero.wall_tracer.stepDistY\[3\]
+ _03033_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_199_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14710__A2 _08233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_225_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19525__I _12296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21013_ _02086_ _02100_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_184_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_225_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23981__A1 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26870_ _00780_ clknet_leaf_165_i_clk rbzero.tex_r0\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_25821_ _05988_ _05993_ _06603_ _06604_ _06605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_149_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25752_ _06528_ _06535_ _06536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22964_ _03691_ _03694_ _03821_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__25262__I _06045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24703_ _05486_ _05452_ _05487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_203_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21915_ _10483_ _10474_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25683_ _06426_ _06466_ _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_179_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22895_ _02573_ _02686_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_27422_ _01327_ clknet_leaf_84_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24634_ _05241_ _05418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14777__A2 _07930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21846_ _02888_ _02890_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_72_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27353_ _01258_ clknet_leaf_81_i_clk rbzero.wall_tracer.trackDistX\[-5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24565_ _05347_ _05348_ _05349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_148_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21777_ _02703_ _02827_ _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26304_ _00214_ clknet_leaf_232_i_clk rbzero.spi_registers.buf_othery\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23516_ _04155_ _04275_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20728_ _01817_ _01818_ _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_27284_ _01189_ clknet_leaf_212_i_clk gpout0.hpos\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24496_ _05058_ _05157_ _05189_ _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16774__I0 rbzero.pov.ready_buffer\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_26235_ _00145_ clknet_leaf_240_i_clk rbzero.spi_registers.texadd2\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23447_ _04280_ _04300_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_123_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20659_ _01749_ _01750_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_162_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13200_ _06997_ _07014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_151_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21275__A2 _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26166_ _00076_ clknet_leaf_223_i_clk rbzero.floor_leak\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__22472__A1 _08750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14180_ _07210_ _07989_ _07976_ _07990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_23378_ _04143_ _04232_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25117_ _05893_ _05900_ _05901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13131_ rbzero.texu_hot\[4\] _06943_ _06945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22329_ _11155_ _03270_ _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16151__A1 _08922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26097_ _00007_ clknet_leaf_229_i_clk rbzero.spi_registers.ss_buffer\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22224__A1 _11391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25048_ _05566_ _05576_ _05832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_13062_ _06877_ _06878_ _06879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__25961__A2 _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14701__A2 _08506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17870_ rbzero.wall_tracer.rayAddendX\[1\] _11014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16821_ _10249_ _10245_ _10251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14465__A1 _08201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26999_ _00909_ clknet_leaf_193_i_clk rbzero.tex_g0\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13268__A2 _07076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19540_ _10289_ _12312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16752_ _10168_ _10190_ _10191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13964_ rbzero.trace_state\[1\] _07774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_233_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15703_ rbzero.spi_registers.texadd2\[16\] _09338_ _09346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_214_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19471_ rbzero.wall_tracer.stepDistX\[-5\] _12243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_16683_ _10093_ _10127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_85_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14217__A1 _07706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13895_ _07705_ _07706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14217__B2 _07685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15634_ rbzero.spi_registers.texadd1\[22\] _09291_ _09295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18422_ rbzero.tex_g1\[29\] rbzero.tex_g1\[28\] _11517_ _11518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15965__A1 _09542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19156__A1 _08149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21205__I _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18353_ _11477_ _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15565_ _09205_ _09243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18903__A1 rbzero.traced_texa\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17304_ _10632_ _10630_ _10633_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14516_ _08295_ _08320_ _08324_ _08325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_18284_ _11419_ _11424_ _11425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15496_ _09150_ _09192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_151_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17235_ rbzero.pov.spi_buffer\[12\] _10582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14447_ _08249_ _08251_ _08254_ _08255_ _08222_ _08256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17166_ _10522_ _10528_ _10529_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_14378_ _07699_ _08023_ _08036_ _08180_ _08187_ _08188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_51_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16117_ _09599_ _09657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13329_ _06884_ _06887_ _06889_ _07143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_229_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17097_ _08126_ _10477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16048_ rbzero.spi_registers.buf_texadd0\[2\] _09597_ _09606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24251__I _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13900__B1 _07706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19807_ rbzero.wall_tracer.size\[7\] rbzero.wall_tracer.size\[6\] _12579_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17999_ _11142_ _11143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__13393__I gpout0.vpos\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19738_ _12449_ _12457_ _12509_ _12510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__13326__C _07139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_239_Right_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15822__B _09430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19669_ _12319_ _12321_ _10217_ _12324_ _12441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_204_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21700_ _02760_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_22680_ rbzero.wall_tracer.trackDistX\[-8\] _03539_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19147__A1 _08155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24140__A1 _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21631_ _09899_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_192_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13431__A2 _07241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24350_ _05044_ _05061_ _05072_ _05133_ _05134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_21562_ _12238_ _02336_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_16_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23301_ _04040_ _04152_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20513_ _01521_ _01522_ _01605_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_144_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24281_ _04988_ _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_21493_ _02525_ _02535_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26020_ _06739_ _06644_ _06655_ _06737_ _06796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_16_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21257__A2 _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20444_ _01518_ _01537_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_23232_ _04084_ _04087_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22454__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24362__S _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23163_ _04018_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_20375_ _01468_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_207_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19870__A2 _12639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22390__B _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22114_ _11081_ _03092_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23094_ _03945_ _03950_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_101_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22045_ rbzero.wall_tracer.stepDistY\[-3\] _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26922_ _00832_ clknet_leaf_130_i_clk rbzero.tex_r1\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_101_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_205_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_205_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26853_ _00763_ clknet_leaf_191_i_clk rbzero.tex_r0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_25804_ _06578_ _06587_ _06588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26784_ _00694_ clknet_leaf_126_i_clk rbzero.tex_g1\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_242_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23996_ _08810_ _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_203_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25735_ _06478_ _06482_ _06519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_173_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22947_ _03782_ _03799_ _03804_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_67_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_206_Right_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13670__A2 _07338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_238_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25666_ _06154_ _05972_ _06407_ _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_197_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13680_ rbzero.tex_r0\[49\] _07484_ _07491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22878_ _02530_ _03736_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27405_ _01310_ clknet_leaf_113_i_clk rbzero.wall_tracer.stepDistX\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_22_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24617_ _05219_ _05366_ _05401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16119__I _08931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21829_ _02859_ _02864_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25597_ _06350_ _06380_ _06381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_65_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24682__A2 _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27336_ _01241_ clknet_leaf_92_i_clk rbzero.trace_state\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15350_ rbzero.mapdxw\[0\] _09075_ _09085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20864__I _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24548_ _05236_ _05331_ _05332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_183_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22693__A1 _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21496__A2 _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14301_ rbzero.debug_overlay.vplaneY\[-4\] _08111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_202_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27267_ _01172_ clknet_leaf_116_i_clk rbzero.wall_tracer.visualWallDist\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15281_ _07165_ _09034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24479_ _05261_ _05215_ _05263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17020_ _08157_ _10410_ _10419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26218_ _00128_ clknet_leaf_16_i_clk rbzero.spi_registers.texadd1\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14232_ rbzero.debug_overlay.playerY\[-7\] _08042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27198_ _01103_ clknet_leaf_77_i_clk rbzero.wall_tracer.size_full\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14163_ _07775_ net2 _07243_ _07972_ _07973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_26149_ _00059_ clknet_leaf_216_i_clk rbzero.map_overlay.i_mapdx\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_247_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13114_ _06927_ rbzero.wall_hot\[1\] _06928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_104_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14094_ _07896_ _07903_ _07904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15907__B _09491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18971_ rbzero.tex_g0\[22\] rbzero.tex_g0\[21\] _11856_ _11858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_221_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17922_ _10999_ _11063_ _11065_ _11066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13045_ _06861_ _06862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_218_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17624__A1 _10845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17853_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] _10997_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_234_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16804_ _09139_ _10236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14996_ _07175_ _08779_ _08775_ _08798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17784_ _10951_ _10695_ _10947_ _10953_ _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_221_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24370__A1 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16738__B _08882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19523_ rbzero.wall_tracer.stepDistY\[-4\] _12256_ _12294_ _12295_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_220_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13947_ _07244_ rbzero.map_overlay.i_mapdy\[0\] _07758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16735_ _10165_ _10173_ _10175_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__21184__A1 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16666_ _10092_ _08116_ _10110_ _10111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__15938__A1 _09522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19454_ _10331_ _12006_ _12226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_158_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13878_ _07684_ _07685_ _07676_ _07686_ _07688_ _07689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__24122__A1 _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15617_ _09280_ _09282_ _09278_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18405_ _11508_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16597_ _10044_ _10045_ _10046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19385_ _07233_ _11380_ _12157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_57_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14610__A1 rbzero.tex_g1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22684__A1 _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18336_ _07214_ _11466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15548_ _09205_ _09230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_84_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18267_ _11409_ _11410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15479_ _09064_ _09180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16363__A1 _08948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17218_ _10567_ _10559_ _10569_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_181_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18198_ _11335_ _11339_ _11341_ _11342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_142_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17149_ _10513_ _10515_ _10516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__26561__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20160_ _12928_ _12931_ _12932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_122_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20091_ _12858_ _12828_ _12863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_181_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19604__A2 _11988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13337__B _07150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23850_ rbzero.wall_tracer.stepDistY\[10\] _04678_ _04679_ _04680_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_240_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22801_ _02098_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15552__B _09229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_23781_ _04586_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21175__A1 _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20993_ _02076_ _02081_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_196_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25520_ _06302_ _06303_ _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_200_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22732_ _03591_ _03593_ _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__15929__A1 _09515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25451_ _06228_ _06232_ _06234_ _06235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_0_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22663_ rbzero.wall_tracer.trackDistX\[-10\] _12214_ _03526_ _03534_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_165_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_196_i_clk_I clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19678__C _12334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24402_ _05011_ _05186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_168_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_21614_ rbzero.wall_tracer.rayAddendX\[-9\] _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25382_ _05982_ _06040_ _06166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22675__A1 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22594_ _12231_ _03089_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_233_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27121_ _01031_ clknet_leaf_117_i_clk rbzero.traced_texVinit\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_233_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24333_ _04940_ _05023_ _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_192_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21545_ _02509_ _02512_ _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_145_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13800__B _07580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13168__A1 rbzero.spi_registers.texadd2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27052_ _00962_ clknet_leaf_144_i_clk rbzero.tex_b1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__22427__A1 rbzero.wall_tracer.texu\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24264_ _05040_ _05041_ _05042_ _05043_ _05045_ _05047_ _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_65_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14904__A2 _07597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21476_ _02560_ _02561_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26003_ _06629_ _06711_ _06781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_121_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23215_ _04047_ _04049_ _04070_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20427_ _12282_ _13023_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24195_ _04852_ _04978_ _04979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_95_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17854__A1 _08071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__27119__D _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23146_ _03899_ _04002_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20358_ _01365_ _01452_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_113_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21650__A2 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14668__B2 _07955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23077_ _03822_ _03827_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20289_ _12235_ _01383_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22028_ rbzero.wall_tracer.stepDistY\[-8\] _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13247__B _07060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26905_ _00815_ clknet_leaf_125_i_clk rbzero.tex_r1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_227_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold41 i_gpout1_sel[3] net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__13891__A2 _07044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_199_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14850_ rbzero.tex_b1\[15\] _08496_ _08339_ _08656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26836_ _00746_ clknet_leaf_196_i_clk rbzero.tex_r0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_188_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23155__A2 _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13801_ rbzero.tex_r0\[9\] _07584_ _07612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_203_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14781_ rbzero.tex_b0\[9\] _08300_ _08588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26767_ _00677_ clknet_leaf_125_i_clk rbzero.tex_g1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23979_ _04739_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_203_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__21166__A1 _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13643__A2 _07448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16520_ _09973_ _09974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25718_ _06385_ _06501_ _06502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_13732_ _07531_ _07543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19869__B _12171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26698_ _00608_ clknet_leaf_62_i_clk rbzero.pov.ready_buffer\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20913__A1 _12661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16451_ _09908_ _09909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_25649_ _06396_ _06414_ _06433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13663_ _07458_ _07473_ _07441_ _07474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__22115__B1 _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15402_ _09064_ _09124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19170_ _12013_ _12014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__22666__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16382_ rbzero.spi_registers.buf_texadd3\[13\] _09851_ _09857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13594_ _07079_ _07393_ _07394_ _06872_ _07404_ _07405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_53_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18121_ _07694_ _11263_ rbzero.map_rom.b6 _10352_ _11264_ _11265_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_27319_ _01224_ clknet_leaf_116_i_clk rbzero.traced_texa\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15333_ _09054_ _09073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13710__B _07520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18052_ rbzero.wall_tracer.trackDistY\[-6\] _11196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_13_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15264_ _07722_ _09019_ _09020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17003_ _10405_ _10406_ _10386_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14215_ _08024_ _08014_ _08025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23091__A1 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15195_ rbzero.spi_registers.spi_buffer\[12\] _08960_ _08967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24015__B _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14146_ _07951_ _07952_ _07954_ _07955_ _07913_ _07956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_6_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16312__I _09746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18954_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _11845_ _11848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14077_ _07854_ _07886_ _07478_ _07887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24591__A1 _05304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23394__A2 _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17905_ _08082_ rbzero.wall_tracer.rayAddendX\[-1\] _11049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_219_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18885_ _11799_ _11800_ _11802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_218_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21944__A3 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21374__B _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17836_ _10857_ rbzero.pov.ready_buffer\[71\] _10986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24343__A1 _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer17 _05525_ net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_222_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18239__I _11382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xrebuffer28 _05382_ net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17767_ _10937_ rbzero.pov.ready_buffer\[46\] _10942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xrebuffer39 _05335_ net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_14979_ _08778_ _08780_ _08781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__13671__I _07481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13634__A2 _07444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14831__A1 rbzero.tex_b1\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19506_ rbzero.wall_tracer.visualWallDist\[-9\] _12277_ _12278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__18022__A1 _11163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16718_ _10159_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_141_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20904__A1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22984__I _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17698_ _10872_ _10896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19437_ _12208_ _12209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_186_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16649_ _10074_ _10091_ _10094_ _10095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24646__A2 _05429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16915__C _10221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19368_ rbzero.tex_b1\[59\] rbzero.tex_b1\[58\] _12146_ _12149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_44_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15598__I _09254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_215_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18319_ _11431_ _11453_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_174_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19299_ rbzero.tex_b1\[29\] rbzero.tex_b1\[28\] _12109_ _12110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_21330_ _02276_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__22409__A1 _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14898__A1 rbzero.tex_b1\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21261_ _02338_ _02347_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__23082__A1 _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23000_ _03729_ _03740_ _03857_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20212_ _12900_ _12922_ _12983_ _12984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_163_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16639__A2 _09971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17836__A1 _10857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21192_ _12299_ _01466_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15547__B _09229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20143_ rbzero.wall_tracer.stepDistY\[1\] _12906_ _12910_ _12914_ _12915_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_110_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_229_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13322__A1 _07045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20074_ _12819_ _12820_ _12846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24951_ _05710_ _05712_ _05735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_23902_ _03019_ _04711_ _04713_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24882_ _05663_ _05664_ _05665_ _05666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_99_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26621_ _00531_ clknet_leaf_162_i_clk rbzero.tex_b0\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_225_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_213_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23833_ _04661_ _04664_ _02730_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_224_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26552_ _00462_ clknet_leaf_66_i_clk rbzero.pov.spi_buffer\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23764_ _04598_ _04589_ _04604_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20976_ _01938_ _01939_ _02064_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_235_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25503_ _06165_ _06168_ _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_211_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17988__I _11131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22715_ _02746_ _02033_ _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__16575__A1 _10024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26483_ _00393_ clknet_leaf_57_i_clk rbzero.debug_overlay.facingX\[-6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_193_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23695_ _11207_ _03037_ _04543_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_25434_ _06214_ _06215_ _06217_ _06218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_22646_ _12775_ _12864_ _02750_ _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_192_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22648__A1 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14050__A2 _07810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19364__I1 rbzero.tex_b1\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25365_ _06111_ _06112_ _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_97_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22577_ _03468_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_134_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27104_ _01014_ clknet_leaf_139_i_clk rbzero.tex_b1\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24316_ _05099_ net93 _05100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_21528_ _02472_ _02475_ _02612_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_133_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25296_ _05945_ _06080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_181_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14889__B2 _08558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27035_ _00945_ clknet_leaf_137_i_clk rbzero.tex_g0\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24247_ _05003_ _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_161_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21459_ _02261_ _12958_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19816__A2 _12587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14000_ _07628_ _07810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_24178_ _04806_ _04948_ _04915_ _04916_ _04962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_31_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput31 net31 o_gpout[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_75_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput42 net42 o_tex_out0 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_102_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17228__I _10564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23129_ _02404_ _03736_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_246_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15951_ _09515_ _09528_ _09533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13864__A2 rbzero.debug_overlay.playerY\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18252__A1 _11391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14902_ _08704_ _08705_ _08707_ _08564_ _07839_ _08708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_15882_ _09457_ _09443_ _09480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18670_ _11659_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17621_ rbzero.pov.spi_done _10843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13705__B _07492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26819_ _00729_ clknet_leaf_180_i_clk rbzero.tex_g1\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14833_ rbzero.tex_b1\[27\] _08568_ _08638_ _08639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_144_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14764_ rbzero.tex_b0\[20\] _08518_ _08570_ _08571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17552_ _10804_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_106_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19752__A1 _12522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16503_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.wall_tracer.rayAddendY\[-3\] _09958_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13715_ _07331_ _07526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17483_ _10759_ _10765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14695_ _07808_ _08502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_128_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19222_ _12059_ _12063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_156_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16434_ _09893_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13646_ _07432_ _07456_ _07457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19153_ _11986_ _11988_ _11989_ _11996_ _11997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_156_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16365_ _09841_ _09843_ _09844_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_156_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13577_ _07356_ _07387_ _07388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15211__I rbzero.spi_registers.spi_buffer\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18104_ _11139_ _11140_ _11237_ _11247_ _11248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_15316_ _08884_ _09060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19084_ rbzero.debug_overlay.facingY\[-8\] _09991_ _11928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_16296_ rbzero.spi_registers.buf_texadd2\[16\] _09791_ _09792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_227_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23064__A1 _12676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18035_ rbzero.wall_tracer.trackDistY\[-2\] _11179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15247_ _09008_ _09001_ _09009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15178_ _08933_ _08954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13666__I _07326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_144_i_clk_I clknet_5_14__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__17138__I _10491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14129_ rbzero.tex_r1\[55\] _07938_ _07917_ _07939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19986_ _12752_ _12753_ _12757_ _12758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_120_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13304__A1 _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18937_ _11838_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18868_ rbzero.traced_texa\[0\] rbzero.texV\[0\] _11785_ _11788_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_193_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24316__A1 _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17819_ _10973_ rbzero.pov.ready_buffer\[64\] _10976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_206_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18799_ _11732_ _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14804__A1 _07803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20830_ _01919_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25090__I _05856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14280__A2 _08064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19743__A1 _12514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_217_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20761_ _01829_ _01851_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__21550__A1 _12777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22500_ rbzero.wall_tracer.size\[7\] _03417_ _03418_ rbzero.row_render.size\[7\]
+ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_69_i_clk_I clknet_5_29__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23480_ _04323_ _04333_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20692_ _01782_ _01770_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19346__I1 rbzero.tex_b1\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22431_ _02033_ _03373_ _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_230_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_230_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25150_ _05887_ _05901_ _05934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_21_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22362_ _03307_ _03309_ _03310_ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_143_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24101_ _04884_ _04885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_28_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19528__I _12299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21313_ _02398_ _02284_ _02399_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_170_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25081_ _05863_ _05864_ _05865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25974__B _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22293_ _11173_ _03239_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24032_ _04772_ _04768_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_13_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22802__A1 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21605__A2 _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21244_ _02330_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_57_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21175_ _02260_ _02262_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_228_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20126_ _12894_ _12897_ _12898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25983_ _06686_ _06732_ _06762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16887__I _10271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20057_ _12742_ _12749_ _12829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24934_ _05687_ _05718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__18234__A1 _11248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_241_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24865_ _05647_ _05648_ _05649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20592__A2 _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23816_ _04646_ _04649_ _04594_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26604_ _00514_ clknet_leaf_36_i_clk rbzero.pov.spi_buffer\[73\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__22869__A1 _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24796_ _05365_ _05470_ _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13244__C _07057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26535_ _00445_ clknet_leaf_22_i_clk rbzero.pov.spi_buffer\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23747_ _04586_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20344__A2 _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21541__A1 _12300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20959_ _01998_ _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_138_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13500_ _07277_ _07310_ _07311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14480_ _07549_ _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26466_ _00376_ clknet_leaf_44_i_clk rbzero.debug_overlay.playerY\[-8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__22129__I _09982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23678_ _04528_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14023__A2 _07832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25417_ _06200_ _06201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13431_ net2 _07241_ _07242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_101_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22629_ _03506_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26397_ _00307_ clknet_leaf_3_i_clk rbzero.spi_registers.buf_texadd2\[17\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_46_Left_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16150_ rbzero.spi_registers.buf_texadd1\[3\] _09672_ _09683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25348_ _06072_ _06093_ _06131_ _06132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13362_ net19 _07154_ _07161_ net27 _07173_ _07174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xrebuffer8 _05435_ net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15101_ _08888_ _08890_ _08891_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_1_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_248_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16081_ _09629_ _09630_ _09626_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_248_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25279_ _06029_ _06062_ _06063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_51_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13293_ _07065_ _06968_ _07104_ _07106_ _07107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__16720__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_248_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27018_ _00928_ clknet_leaf_169_i_clk rbzero.tex_g0\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_15032_ _08823_ _08824_ _08825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19840_ _12601_ _12612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15287__A1 rbzero.spi_registers.buf_othery\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23349__A2 _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20280__A1 _12962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19771_ _12539_ _12540_ _12541_ _12542_ _12543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_16983_ _10389_ _10390_ _10386_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13298__B1 _07035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24012__C _11473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18722_ rbzero.tex_r1\[30\] rbzero.tex_r1\[29\] _11687_ _11689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_108_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15934_ _09504_ _09520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20112__I _12409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18653_ _11478_ _11649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15865_ _08924_ _09459_ _09468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16787__A1 _07700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17604_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _10833_ _10834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14816_ _07789_ _07798_ _08623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18584_ _11610_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_121_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15796_ rbzero.spi_registers.texadd3\[16\] _09407_ _09415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17535_ _10794_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_158_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14747_ _07811_ _08554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_70_i_clk_I clknet_5_29__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14678_ _08485_ _07668_ _08486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17466_ rbzero.pov.spi_buffer\[72\] _10544_ _10751_ _10754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14014__A2 _07821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19205_ rbzero.wall_tracer.mapY\[7\] _12048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_104_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16417_ _09881_ _09882_ _09878_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13629_ _07435_ _07440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17397_ rbzero.pov.spi_buffer\[54\] _10697_ _10693_ _10703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_171_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19136_ _11955_ _11979_ _11945_ _11980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24254__I _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16348_ _08926_ _09831_ _09832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19067_ net25 rbzero.tex_g0\[63\] _11908_ _11912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16279_ _09778_ _09779_ _09773_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18018_ _11161_ _11162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_160_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19969_ _12682_ _12720_ _12740_ _12741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15825__B _09430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22502__I _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22980_ _03721_ _03836_ _03837_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_52_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19964__A1 _12728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21931_ _02963_ _10087_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_241_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_242_i_clk clknet_5_0__leaf_i_clk clknet_leaf_242_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_24650_ _05340_ _05339_ _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21862_ _02891_ _02900_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__19716__A1 _12261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23601_ _03713_ _04308_ _04406_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20813_ _01857_ _01884_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24581_ _05364_ _05365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21793_ _08131_ rbzero.debug_overlay.vplaneX\[-9\] _02841_ _02842_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_26320_ _00230_ clknet_leaf_236_i_clk rbzero.spi_registers.buf_mapdx\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__21989__S _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23532_ _03861_ _04180_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20744_ _12696_ _12593_ _01620_ _01834_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_9_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__25265__A2 _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26251_ _00161_ clknet_leaf_2_i_clk rbzero.spi_registers.texadd2\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23463_ _04311_ _04316_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20675_ _01741_ _01766_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16950__A1 _10358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25202_ _05981_ _05984_ _05985_ _05986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_162_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22414_ _03346_ _03358_ _03323_ _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26182_ _00092_ clknet_leaf_188_i_clk rbzero.spi_registers.vshift\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_23394_ _04124_ _04125_ _04128_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14904__B _08603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25133_ _05915_ _05916_ _05917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22345_ _11147_ _03245_ _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14690__I _07546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18162__I _11256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23028__A1 _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25064_ _05413_ _05332_ _05848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22276_ _11190_ _03239_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24015_ rbzero.wall_tracer.rcp_fsm.i_start _06895_ _04799_ _04800_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_72_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21227_ _02293_ _02299_ _02313_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_243_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20262__A1 _12955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21158_ _02244_ _02245_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_208_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20109_ _12627_ _12630_ _12881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_205_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16410__I _09855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13980_ _07196_ _07790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25966_ _06627_ _06733_ _06624_ _06622_ _06697_ _06699_ _06746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_21089_ _02054_ _02164_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_245_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14492__A2 _08300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23751__A2 _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24917_ _05661_ _05662_ _05664_ _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_25897_ _06666_ _06675_ _06679_ _06680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_232_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21762__A1 _09945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15650_ _09304_ _09307_ _09301_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24848_ _05599_ _05631_ _05632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_38_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19707__A1 _12439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24700__A1 _05460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14601_ rbzero.tex_g1\[10\] _07635_ _08408_ _08409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_201_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15581_ _09254_ _09255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24779_ _05283_ net65 _05563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17320_ rbzero.pov.spi_buffer\[34\] _10645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14532_ rbzero.tex_g0\[61\] _08340_ _08341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26518_ _00428_ clknet_leaf_57_i_clk rbzero.debug_overlay.vplaneY\[-4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_83_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_54_Left_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14463_ _08264_ _08271_ _08272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17251_ _10571_ _10594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26449_ _00359_ clknet_leaf_88_i_clk rbzero.wall_tracer.rayAddendY\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15744__A2 _09373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16941__A1 rbzero.pov.ready_buffer\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16202_ _08990_ _09721_ _09722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13414_ _07224_ _07225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_153_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17182_ rbzero.pov.ss_buffer\[1\] _10514_ _10541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_221_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14394_ rbzero.tex_g0\[29\] _08202_ _08203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16133_ rbzero.spi_registers.spi_done _08833_ _09669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_13345_ net13 _07157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16064_ rbzero.spi_registers.buf_texadd0\[6\] _09610_ _09618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13276_ _06945_ _06973_ _07090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15015_ _08813_ _08814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_114_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_17_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Left_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_131_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19823_ rbzero.wall_tracer.visualWallDist\[-10\] _12595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_235_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25192__A1 _05333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19754_ _12382_ _12525_ _12526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16966_ _08876_ _10163_ _10377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_223_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14483__A2 _08291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19946__A1 _12714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18705_ _11679_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15917_ _09497_ _09507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19685_ _12450_ _12451_ _12457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_223_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18213__A4 _11308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16897_ _10295_ _10317_ _10318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21753__A1 _10466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19631__I _12402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18636_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _11639_ _11640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_189_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15848_ _09140_ _09453_ _09454_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_8_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__18247__I _11390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18567_ _11600_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15779_ rbzero.spi_registers.buf_texadd3\[11\] _09398_ _09403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_72_Left_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17518_ rbzero.tex_b0\[20\] rbzero.tex_b0\[19\] _10781_ _10785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18498_ rbzero.tex_g1\[62\] rbzero.tex_g1\[61\] _11559_ _11561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17449_ _10739_ _10735_ _10741_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16932__A1 _10346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20460_ _09939_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19119_ _08160_ rbzero.wall_tracer.rayAddendY\[-1\] _11963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20391_ _01483_ _01484_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22130_ _03089_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20017__I _12706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_81_Left_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22061_ _03063_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14015__I _07492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_225_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21012_ _02086_ _02100_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_184_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_225_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23981__A2 _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22232__I _11248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15555__B _09229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16999__A1 rbzero.pov.ready_buffer\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13854__I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25820_ _06582_ _06598_ _06596_ _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_149_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16230__I _09741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23772__B _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17660__A2 rbzero.pov.ready_buffer\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_181_i_clk clknet_5_8__leaf_i_clk clknet_leaf_181_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25751_ _06531_ _06534_ _06535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_208_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input29_I i_vec_sclk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22963_ _02501_ _02115_ _03692_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_65_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18204__A4 _11107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24702_ _05454_ _05485_ _05486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_21914_ _10483_ _10474_ _10471_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_25682_ _06427_ _06465_ _06466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__20687__I _09939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_203_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22894_ _03750_ _03752_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_27421_ _01326_ clknet_leaf_84_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24633_ _05409_ _05415_ _05416_ _05417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23497__A1 _11410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13803__B _07613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21845_ _02888_ _02890_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18157__I _11269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15974__A2 _08831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_196_i_clk clknet_5_12__leaf_i_clk clknet_leaf_196_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_172_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27352_ _01257_ clknet_leaf_80_i_clk rbzero.wall_tracer.trackDistX\[-6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24564_ _05313_ _05328_ _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_66_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21776_ _10022_ _02821_ _02826_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_23515_ _04155_ _04031_ _04162_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_26303_ _00213_ clknet_leaf_236_i_clk rbzero.spi_registers.buf_otherx\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_65_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20727_ _12885_ _12645_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27283_ _01188_ clknet_leaf_212_i_clk gpout0.hpos\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24495_ _05256_ _05277_ _05278_ _05279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_175_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16774__I1 _10208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26234_ _00144_ clknet_leaf_247_i_clk rbzero.spi_registers.texadd2\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23446_ _04283_ _04299_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_163_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20658_ _12208_ _01641_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_135_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26165_ _00075_ clknet_leaf_184_i_clk rbzero.floor_leak\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23377_ _04190_ _04231_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20589_ _01606_ _01623_ _01680_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25116_ _05894_ _05899_ _05900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13130_ rbzero.texu_hot\[4\] _06943_ _06944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22328_ rbzero.wall_tracer.trackDistY\[5\] _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26096_ _00006_ clknet_leaf_230_i_clk rbzero.spi_registers.mosi vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_134_i_clk clknet_5_15__leaf_i_clk clknet_leaf_134_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25047_ _05767_ _05799_ _05831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13061_ gpout0.hpos\[4\] _06878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__22224__A2 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22259_ _03203_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13764__I _07482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17236__I _10571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16820_ _10249_ _10245_ _10250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__16140__I _09675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_149_i_clk clknet_5_11__leaf_i_clk clknet_leaf_149_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_26998_ _00908_ clknet_leaf_172_i_clk rbzero.tex_g0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14465__A2 _08273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15662__A1 rbzero.spi_registers.texadd2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__23724__A2 _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16751_ _08172_ _10189_ _10190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25949_ _06677_ _06673_ _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13963_ _07186_ _07772_ _07773_ net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__19451__I _12222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15702_ _09344_ _09345_ _09337_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19470_ _12241_ _12242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_232_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_214_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16682_ _10126_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_85_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13894_ rbzero.debug_overlay.playerY\[-3\] _07705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14217__A2 _08023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_243_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18421_ _11501_ _11517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15633_ _09292_ _09294_ _09290_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18352_ _11474_ rbzero.spi_registers.sclk_buffer\[1\] _11477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_57_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15564_ _09238_ _09239_ _09242_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22160__A1 _11287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22160__B2 _11070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17303_ rbzero.pov.spi_buffer\[30\] _10627_ _10624_ _10633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_230_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14515_ _08321_ _08322_ _08323_ _08324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_185_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15495_ _09188_ _09189_ _09191_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18283_ _11399_ _11424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_232_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16914__A1 rbzero.pov.ready_buffer\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17234_ _10579_ _10572_ _10581_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22317__I _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14446_ _07601_ _08255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_181_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21221__I _09900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16315__I _09806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17165_ rbzero.pov.spi_counter\[3\] _10527_ _10529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_80_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14377_ _08183_ _08185_ _08186_ _08187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_12_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16116_ rbzero.spi_registers.buf_texadd0\[20\] _09655_ _09656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13328_ _06871_ _06861_ _06879_ _07142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_17096_ _10475_ _10476_ _10462_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19626__I _12397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16047_ _09604_ _09605_ _09603_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13259_ _06990_ _06995_ _07073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20226__A1 _12486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13900__A1 gpout0.vpos\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13900__B2 _07707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19806_ _12577_ _11068_ _12180_ _12578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__17642__A2 rbzero.pov.ready_buffer\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22987__I _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17998_ rbzero.wall_tracer.trackDistY\[9\] _11142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14456__A2 _07816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19737_ _12450_ _12451_ _12509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16949_ rbzero.pov.ready_buffer\[56\] _10260_ _10360_ _10362_ _10293_ _10363_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__21726__A1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_220_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_220_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19668_ rbzero.wall_tracer.visualWallDist\[-3\] _11381_ _11382_ _12440_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_126_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15405__A1 _08485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18619_ _11630_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_189_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19599_ _12353_ _12370_ _12371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_56_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24140__A2 _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21630_ _02308_ _02706_ _02707_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22151__A1 _11989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21561_ _02496_ _02516_ _02645_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_16_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23300_ _03918_ _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13719__A1 _07480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20512_ _12685_ _01523_ _01604_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_24280_ _05013_ _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_28_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21492_ _02521_ _02557_ _02576_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23231_ _04085_ _04086_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20443_ _01520_ _01523_ _01536_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__21257__A3 _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_51_i_clk clknet_5_23__leaf_i_clk clknet_leaf_51_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23162_ _03908_ _03995_ _04017_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_20374_ rbzero.wall_tracer.visualWallDist\[4\] _12199_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22113_ _03104_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_219_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23093_ _03946_ _03949_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__15892__A1 _08928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_192_i_clk_I clknet_5_9__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22044_ _03052_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26921_ _00831_ clknet_leaf_130_i_clk rbzero.tex_r1\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
Xclkbuf_leaf_66_i_clk clknet_5_21__leaf_i_clk clknet_leaf_66_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_205_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_26852_ _00762_ clknet_leaf_191_i_clk rbzero.tex_r0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__17633__A2 _10538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_205_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25803_ _06579_ _06586_ _06587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_23995_ rbzero.wall_tracer.rcp_fsm.i_data\[6\] _04770_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26783_ _00693_ clknet_leaf_126_i_clk rbzero.tex_g1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_203_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19271__I _12093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_170_Right_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25734_ _06506_ _06516_ _06517_ _06518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22946_ _03800_ _03803_ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22390__A1 _12577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_23__f_i_clk_I clknet_3_5_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14629__B _07819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_238_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25665_ _06154_ _05972_ _06407_ _06449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_197_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22877_ _01380_ _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_238_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_197_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27404_ _01309_ clknet_leaf_111_i_clk rbzero.wall_tracer.stepDistX\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24616_ _05295_ _05399_ _05400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_21828_ _10481_ _11075_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25596_ _06277_ _06378_ _06379_ _06380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_155_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24547_ _05230_ _05331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_27335_ _01240_ clknet_leaf_93_i_clk rbzero.trace_state\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21759_ _09923_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18897__A1 rbzero.traced_texa\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22693__A2 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14300_ _08109_ _08110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15280_ rbzero.spi_registers.buf_otherx\[4\] _09032_ _09033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24478_ _05261_ _05216_ _05262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_191_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22137__I _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27266_ _01171_ clknet_leaf_96_i_clk rbzero.wall_tracer.visualWallDist\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13759__I _07348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14231_ rbzero.debug_overlay.playerY\[-6\] _08041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_26217_ _00127_ clknet_leaf_16_i_clk rbzero.spi_registers.texadd1\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_19_i_clk clknet_5_5__leaf_i_clk clknet_leaf_19_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_23429_ _04176_ _04281_ _04282_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_27197_ _01102_ clknet_leaf_74_i_clk rbzero.wall_tracer.size_full\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22581__B _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14162_ _07717_ _07800_ _07970_ _07971_ _07972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_26148_ _00058_ clknet_leaf_216_i_clk rbzero.map_overlay.i_mapdx\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14135__A1 rbzero.tex_r1\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13113_ rbzero.wall_hot\[0\] _06927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26079_ _06802_ _03019_ _06844_ _06845_ _06810_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_21_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14093_ _07897_ _07899_ _07900_ _07902_ _07638_ _07903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_18970_ _11857_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_111_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17921_ _08071_ _11064_ _11065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_hold37_I i_gpout0_sel[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13044_ gpout0.hpos\[6\] _06861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19074__A1 _08151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17852_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] _10996_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_227_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_245_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16803_ _09462_ _10227_ _10235_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_206_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17783_ _10952_ rbzero.pov.ready_buffer\[51\] _10953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14995_ _08775_ _08794_ _08795_ _08796_ _08797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_19522_ _11383_ _12294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_205_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24370__A2 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16734_ _08182_ _10165_ _10174_ _10175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13946_ _07756_ _07757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_159_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19453_ _12194_ _12225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16665_ _10092_ _08103_ _10110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13877_ _07687_ _06864_ _07688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_18404_ rbzero.tex_g1\[21\] rbzero.tex_g1\[20\] _11507_ _11508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15616_ rbzero.spi_registers.buf_texadd1\[17\] _09281_ _09282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_243_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19384_ rbzero.hsync _11826_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22133__A1 _11992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16596_ _10005_ _10026_ _10023_ _10045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14610__A2 _07563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18335_ _11462_ _11463_ _11465_ _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_15547_ _09227_ _09228_ _09229_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__18888__A1 rbzero.traced_texa\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23881__A1 rbzero.wall_tracer.stepDistX\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22684__A2 _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18266_ _11397_ _11409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_170_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15478_ _09177_ _09179_ _09175_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13669__I _07479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17217_ rbzero.pov.spi_buffer\[8\] _10568_ _10565_ _10569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14429_ _07574_ _08231_ _08237_ _08238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_114_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18197_ _11111_ _11340_ _11341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23633__A1 _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17148_ _10514_ _10515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24262__I _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14126__B2 _07912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17079_ _10463_ _10443_ _10464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20090_ _12768_ _12772_ _12862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_181_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13885__B1 _07677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22800_ _03650_ _03653_ _03658_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23780_ _11167_ _04589_ _04618_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_211_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20992_ _02077_ _02080_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_200_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22731_ _03591_ _03593_ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_200_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15124__I _08805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25450_ _06233_ _06199_ _06234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_177_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22662_ rbzero.wall_tracer.stepDistX\[-9\] _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_133_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_139_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24401_ _05118_ _05183_ _05184_ _05185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__13404__A3 _07214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14601__A2 _07635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21613_ _02692_ _02693_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25381_ _05948_ _06046_ _06165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23872__A1 rbzero.wall_tracer.rcp_fsm.o_data\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22593_ _03321_ _03475_ _03479_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_233_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24332_ _05100_ _05102_ _05115_ _05082_ _05004_ _05116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_146_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27120_ _01030_ clknet_leaf_118_i_clk rbzero.traced_texVinit\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_233_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21544_ _02510_ _02511_ _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_192_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27051_ _00961_ clknet_leaf_121_i_clk rbzero.wall_tracer.mapY\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24263_ _05046_ _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__23624__A1 _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21475_ _02459_ _02559_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26002_ _06629_ _06778_ _06779_ _06780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23214_ _04057_ _04061_ _04069_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20426_ _01415_ _01418_ _01519_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24194_ _04858_ _04859_ _04978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_114_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14117__A1 _07889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25377__A1 _06148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23145_ _03997_ _04001_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20357_ _01369_ _01451_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23927__A2 _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23076_ _03915_ _03932_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20288_ _12448_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21938__A1 _10478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_22027_ _02990_ _03031_ _03040_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26904_ _00814_ clknet_leaf_125_i_clk rbzero.tex_r1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__20610__A1 _12731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold42 net11 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_243_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_199_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15743__B _09372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26835_ _00745_ clknet_leaf_196_i_clk rbzero.tex_r0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__16290__A1 rbzero.spi_registers.spi_buffer\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13800_ rbzero.tex_r0\[10\] _07460_ _07580_ _07611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_230_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14780_ rbzero.tex_b0\[8\] _07629_ _08587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26766_ _00676_ clknet_leaf_230_i_clk rbzero.spi_registers.sclk_buffer\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_203_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23978_ rbzero.wall_tracer.rcp_fsm.operand\[2\] _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13643__A3 _07449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14840__A2 _07595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25717_ _06496_ _06500_ _06501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13731_ _07533_ _07536_ _07538_ _07540_ _07541_ _07542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_22929_ _01948_ _01952_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26697_ _00607_ clknet_leaf_63_i_clk rbzero.pov.ready_buffer\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16042__A1 _09591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16450_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] _09907_
+ _09908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25648_ _06396_ _06414_ _06432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__24347__I _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13662_ _07422_ _07472_ rbzero.row_render.texu\[0\] _07473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_85_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22115__A1 _11994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22115__B2 rbzero.wall_tracer.visualWallDist\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15401_ _09114_ _09122_ _09123_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_16381_ _09852_ _09854_ _09856_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13593_ _07402_ _07403_ _07404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25579_ _05234_ _06041_ _06363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23863__A1 _12214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18120_ rbzero.debug_overlay.playerX\[4\] _11259_ _11264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27318_ _01223_ clknet_leaf_117_i_clk rbzero.traced_texa\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14806__C _08357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15332_ rbzero.spi_registers.buf_mapdy\[1\] _09060_ _09072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18051_ rbzero.wall_tracer.trackDistX\[-6\] _11195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_163_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27249_ _01154_ clknet_leaf_99_i_clk rbzero.wall_tracer.visualWallDist\[-11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15263_ _08878_ _09019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17002_ rbzero.pov.ready_buffer\[40\] _10383_ _10406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14214_ _07999_ _08000_ _08024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_112_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21626__B1 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15194_ _08964_ _08966_ _08954_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_50_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__23091__A2 _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25368__A1 _06034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14145_ _07539_ _07955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14659__A2 _07641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18953_ _11847_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14076_ _07803_ _07862_ _07869_ _07875_ _07885_ _07886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_238_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19904__I _12430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17904_ rbzero.debug_overlay.facingX\[-8\] _11047_ _11048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_219_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14113__I _07546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18884_ _11799_ _11800_ _11801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_128_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17835_ _10979_ _10750_ _10982_ _10985_ _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_222_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24343__A2 _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer18 _05024_ net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17766_ _10935_ _10679_ _10939_ _10941_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xrebuffer29 _05811_ net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_14978_ net8 _08780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_222_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19505_ _12256_ _12277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14831__A2 _08518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16717_ _10150_ _10158_ _10125_ _10159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_18_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13929_ rbzero.map_overlay.i_mapdx\[5\] _07740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_17697_ _10889_ _10610_ _10892_ _10895_ _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__20904__A2 _11390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16033__A1 _09515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19436_ _12203_ _12207_ _12208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_186_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16648_ _10093_ _10073_ _10094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_140_i_clk_I clknet_5_14__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22106__A1 _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15879__I _08908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19367_ _12148_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23854__A1 _09896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16579_ _10023_ _10026_ _10028_ _10029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_44_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18255__I _11397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18318_ _07712_ _11449_ _11445_ _11452_ _11453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19298_ _12093_ _12109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_84_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_199_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18249_ rbzero.wall_tracer.rcp_done _11392_ _11393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14898__A2 _08631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21260_ _02339_ _02346_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_163_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20211_ _12883_ _12899_ _12983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21093__A1 _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21191_ _12713_ _01469_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_14__f_i_clk clknet_3_3_0_i_clk clknet_5_14__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_229_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20840__A1 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20142_ _12911_ _12913_ _12277_ _12914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_65_i_clk_I clknet_5_21__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20073_ _12832_ _12840_ _12844_ _12845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24950_ _05727_ _05732_ _05733_ _05734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_244_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22593__A1 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23901_ _04009_ _04704_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22240__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24881_ _05661_ _05662_ _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_225_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16272__A1 _08955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24876__B _05640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26620_ _00530_ clknet_leaf_162_i_clk rbzero.tex_b0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23832_ _04662_ _04663_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_213_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24368__S _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23763_ _04533_ _04603_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26551_ _00461_ clknet_leaf_65_i_clk rbzero.pov.spi_buffer\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_200_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20975_ _12429_ _01712_ _01940_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_164_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_194_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_235_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25502_ _06166_ _06167_ _06286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_194_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22714_ rbzero.wall_tracer.trackDistX\[-3\] _12374_ _03578_ _03579_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_178_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23694_ _11209_ rbzero.wall_tracer.stepDistY\[-10\] _04538_ _04543_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_26482_ _00392_ clknet_leaf_62_i_clk rbzero.debug_overlay.facingX\[-7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16575__A2 _08105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25433_ _06029_ _06062_ _06216_ _06217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_22645_ rbzero.wall_tracer.trackDistX\[-11\] _12395_ _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25364_ _06142_ _06144_ _06147_ _06148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_36_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22576_ _11296_ _09974_ _01553_ rbzero.traced_texa\[10\] _03468_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_146_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27103_ _01013_ clknet_leaf_138_i_clk rbzero.tex_b1\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_21527_ _02473_ _02474_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_24315_ _05056_ _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_134_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25295_ _05910_ _06079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_35_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24246_ _04940_ _04992_ _04995_ _05030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_27034_ _00944_ clknet_leaf_137_i_clk rbzero.tex_g0\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_21458_ _02379_ _02380_ _02543_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15738__B _09372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20409_ _01501_ _01412_ _01502_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_24177_ _04881_ _04850_ _04887_ _04960_ _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_0_31_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21389_ _02473_ _02474_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_75_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput32 net32 o_gpout[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23128_ _02250_ _03734_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20831__A1 _12841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net45 o_tex_sclk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_246_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_246_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23059_ _03793_ _03796_ _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15950_ rbzero.spi_registers.buf_vshift\[1\] _09531_ _09532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__21387__A2 _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14901_ rbzero.tex_b1\[50\] _07829_ _08706_ _08707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__18252__A2 _11394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15881_ _08912_ _09477_ _09479_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_204_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16263__A1 _08944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17620_ _10842_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26818_ _00728_ clknet_leaf_181_i_clk rbzero.tex_g1\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14832_ rbzero.tex_b1\[26\] _08291_ _08638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_216_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13077__A1 _06892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14089__B _07819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13616__A3 _07425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17551_ rbzero.tex_b0\[34\] rbzero.tex_b0\[33\] _10802_ _10804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__19201__A1 _12036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19052__I1 rbzero.tex_g0\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14763_ rbzero.tex_b0\[21\] _08448_ _08570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_86_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_106_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26749_ _00659_ clknet_leaf_119_i_clk rbzero.wall_tracer.mapX\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_230_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16502_ rbzero.debug_overlay.vplaneY\[-3\] _09948_ _09957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20898__A1 _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13714_ rbzero.tex_r0\[60\] _07523_ _07524_ _07525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__24089__A1 _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17482_ _10764_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14694_ rbzero.tex_b0\[52\] _08499_ _08500_ _08501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14817__B _07149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19221_ _12056_ _12062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16433_ _09892_ net27 _09893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13645_ _07447_ _07455_ _07456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_184_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19152_ _11990_ _11991_ _11992_ _11995_ _11996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_186_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16364_ _09806_ _09844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13576_ _07362_ _07386_ _07387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_156_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18103_ _11246_ _11247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15315_ _07736_ _09058_ _09059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19083_ rbzero.debug_overlay.facingY\[-7\] _10007_ _11927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16295_ _09741_ _09791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18034_ rbzero.wall_tracer.trackDistY\[-1\] _11178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_151_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15246_ rbzero.spi_registers.spi_buffer\[21\] _09008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15177_ _08950_ _08952_ _08953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20822__A1 _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14128_ _07513_ _07938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19985_ _12754_ _12755_ _12756_ _12757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__24013__A1 rbzero.wall_tracer.rcp_done vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24564__A2 _05328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18936_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _11835_ _11838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14059_ _07863_ _07864_ _07866_ _07867_ _07868_ _07869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_182_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input3_I i_debug_vec_overlay vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18867_ rbzero.traced_texa\[1\] rbzero.texV\[1\] _11787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_118_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13682__I _07492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17818_ _09035_ _10975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_234_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22327__A1 _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18798_ rbzero.tex_r1\[63\] rbzero.tex_r1\[62\] _11729_ _11732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20338__B1 _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17749_ _10915_ _10930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_178_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19743__A2 _12171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_217_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20760_ _01831_ _01850_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_176_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19419_ rbzero.wall_tracer.stepDistX\[-11\] _12161_ _12190_ _12191_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_159_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20691_ _01668_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15402__I _09064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22430_ _03321_ _07700_ _03372_ _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_230_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_230_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22361_ rbzero.mapdxw\[0\] _03307_ _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13791__A2 _07600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24100_ _04843_ _04883_ _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_32_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21312_ _02266_ _02285_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25080_ _05827_ _05802_ _05862_ _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_22292_ _03220_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15558__B _09229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13857__I _07425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24031_ rbzero.wall_tracer.rcp_fsm.operand\[0\] rbzero.wall_tracer.rcp_fsm.operand\[-1\]
+ rbzero.wall_tracer.rcp_fsm.operand\[-2\] rbzero.wall_tracer.rcp_fsm.operand\[-3\]
+ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_142_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21243_ _02328_ _02329_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14740__A1 rbzero.tex_b0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21174_ _02261_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_228_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20125_ _12895_ _12896_ _12897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_229_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25982_ _06727_ _06728_ _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22566__A1 _11283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22566__B2 rbzero.traced_texa\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20056_ _12825_ _12827_ _12828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_24933_ _05692_ _05715_ _05716_ _05717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__18234__A2 _11377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19431__A1 _12194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_70_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_241_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24864_ _05644_ _05646_ _05648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_240_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__27413__D _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26603_ _00513_ clknet_leaf_38_i_clk rbzero.pov.spi_buffer\[72\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23815_ _04647_ _04648_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24795_ _04919_ _05530_ _05579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_213_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26534_ _00444_ clknet_leaf_22_i_clk rbzero.pov.spi_buffer\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_240_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23746_ _11179_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_184_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20958_ _01991_ _02025_ _02046_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16408__I _09818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26465_ _00375_ clknet_leaf_44_i_clk rbzero.debug_overlay.playerY\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20889_ rbzero.wall_tracer.stepDistY\[8\] _01838_ _01839_ _01978_ _01979_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_23677_ _04527_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25416_ _06037_ _06103_ _06199_ _06200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_166_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13430_ _07240_ _07241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19498__A1 rbzero.wall_tracer.size\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22628_ rbzero.wall_tracer.texu\[4\] rbzero.texu_hot\[4\] _03503_ _03506_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_26396_ _00306_ clknet_leaf_3_i_clk rbzero.spi_registers.buf_texadd2\[16\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13361_ net14 _07172_ _07173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25347_ _06071_ _06060_ _06131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_180_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22559_ _03458_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13782__A2 _07592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_101_Left_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15100_ rbzero.spi_registers.spi_counter\[0\] _08889_ _08891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xrebuffer9 net52 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_248_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16080_ _08965_ _09624_ _09630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13292_ _07049_ _07105_ _07045_ _07106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_248_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25278_ _06060_ _06061_ _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_210_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16720__A2 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_248_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27017_ _00927_ clknet_leaf_169_i_clk rbzero.tex_g0\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_15031_ rbzero.spi_registers.spi_cmd\[2\] _08824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24229_ _04986_ _05013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14731__B2 _07463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19670__A1 rbzero.debug_overlay.playerX\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19770_ _12461_ _12505_ _12542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_219_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16982_ rbzero.pov.ready_buffer\[36\] _10383_ _10390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18721_ _11688_ _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15933_ _09518_ _09508_ _09519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18652_ _11648_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15864_ rbzero.spi_registers.buf_floor\[2\] _09464_ _09467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22309__A1 rbzero.wall_tracer.trackDistY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17603_ _10822_ _10833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14815_ _07764_ _07776_ _08622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_204_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18583_ rbzero.tex_r0\[34\] rbzero.tex_r0\[33\] _11608_ _11610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15795_ _09413_ _09414_ _09406_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_121_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17702__I _10884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17534_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _10791_ _10794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14746_ rbzero.tex_b0\[26\] _08528_ _08553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14547__B _08355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17465_ rbzero.pov.spi_buffer\[71\] _10753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14677_ rbzero.color_sky\[3\] _08485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_86_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19204_ _12033_ _12034_ _12045_ _12046_ _12047_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_16416_ rbzero.spi_registers.spi_buffer\[22\] _09876_ _09882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13628_ _07438_ _07439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_41_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17396_ rbzero.pov.spi_buffer\[53\] _10702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_19135_ _11956_ _11977_ _11978_ _11979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_171_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14970__A1 _08747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16347_ _09819_ _09831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13559_ rbzero.row_render.size\[0\] _07370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18161__A1 _11300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19066_ _11911_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__23037__A2 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16278_ rbzero.spi_registers.spi_buffer\[11\] _09771_ _09779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13677__I _07335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18017_ rbzero.wall_tracer.trackDistY\[4\] _11161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15229_ _08994_ _08984_ _08995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_238_i_clk_I clknet_5_4__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16988__I _10377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16475__A1 _09928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19968_ _12725_ _12739_ _12740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22548__A1 _11287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_226_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18919_ _11456_ _11827_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_226_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19899_ _12611_ _12655_ _12670_ _12671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_52_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19964__A2 _12733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21930_ _02951_ _10478_ _02959_ _02969_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_179_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21861_ _10482_ _02904_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23600_ _03713_ _04308_ _04406_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__15450__A2 _09159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20812_ _01858_ _01883_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_222_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24580_ _05238_ _05363_ _05282_ _05364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_21792_ _02836_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_148_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22720__A1 _11175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_159_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20743_ rbzero.wall_tracer.stepDistX\[6\] _01715_ _01833_ _01834_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_147_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23531_ _04293_ _04296_ _04383_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23462_ _04312_ _04315_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_161_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26250_ _00160_ clknet_leaf_2_i_clk rbzero.spi_registers.texadd2\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24445__I _05228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20674_ _01742_ _01765_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16950__A2 _10283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25201_ _05978_ _05985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_190_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19539__I _12310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22413_ _03354_ _03357_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_23393_ _04124_ _04125_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14961__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26181_ _00091_ clknet_leaf_188_i_clk rbzero.spi_registers.vshift\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_45_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25132_ _05783_ _05321_ _05916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22344_ rbzero.wall_tracer.trackDistY\[8\] _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__24225__A1 _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25063_ _05778_ _05779_ _05847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22275_ _03205_ _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24014_ _06901_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_72_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21226_ _02296_ _02297_ _02295_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_72_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_243_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21157_ _02142_ _02158_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20108_ _12627_ _12630_ _12880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_208_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_233_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25965_ _05058_ _06745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21088_ _02054_ _02164_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_232_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20039_ _12810_ _12808_ _12811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24916_ _05698_ _05699_ _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25896_ _06666_ _06678_ _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_217_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_24847_ _05603_ _05628_ _05630_ _05631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_198_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22011__I0 rbzero.wall_tracer.rcp_fsm.o_data\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14600_ rbzero.tex_g1\[11\] _07591_ _08408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_103_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15580_ _09204_ _09254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_205_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24778_ _05505_ _05506_ _05562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26517_ _00427_ clknet_leaf_58_i_clk rbzero.debug_overlay.vplaneY\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14531_ _07831_ _08340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_23729_ _04542_ _04573_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_187_i_clk_I clknet_5_9__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14086__C _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17250_ rbzero.pov.spi_buffer\[16\] _10593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_26448_ _00358_ clknet_leaf_88_i_clk rbzero.wall_tracer.rayAddendY\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14462_ _08262_ _08267_ _08270_ _08271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_138_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16201_ _09674_ _09721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15977__I _09504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13413_ _06866_ gpout0.hpos\[8\] _06882_ _07224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_183_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17181_ _10538_ _10539_ _10540_ _10357_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_221_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26379_ _00289_ clknet_leaf_250_i_clk rbzero.spi_registers.buf_texadd1\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14393_ _07916_ _08202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16132_ _09666_ _09668_ _09661_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13344_ _07153_ _07154_ _07155_ _07156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14704__A1 _08264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16063_ _09616_ _09617_ _09615_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13275_ _07084_ _07085_ _07087_ _07088_ _07074_ _07053_ _07089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_15014_ _08812_ _08813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_184_Right_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_131_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19822_ _12520_ _12594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_224_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_208_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19753_ _12262_ _12525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16965_ _08082_ _10375_ _10376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16209__A1 _08997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_223_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15916_ rbzero.spi_registers.buf_otherx\[3\] _09495_ _09506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18704_ rbzero.tex_r1\[22\] rbzero.tex_r1\[21\] _11677_ _11679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_19684_ _12394_ _12454_ _12455_ _12456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_204_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16896_ rbzero.debug_overlay.playerY\[-4\] _10316_ _10317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_204_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18635_ _11628_ _11639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15847_ _08937_ _09446_ _09454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15432__A2 _08885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18566_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _11597_ _11600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_188_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15778_ rbzero.spi_registers.texadd3\[11\] _09396_ _09402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17517_ _10784_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14729_ rbzero.tex_b0\[45\] _08529_ _08536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_86_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18497_ _11560_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17448_ rbzero.pov.spi_buffer\[67\] _10732_ _10740_ _10741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14943__A1 rbzero.hsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17379_ _10687_ _10688_ _10689_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_132_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19118_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] _11962_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20390_ _12690_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16696__A1 _09998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19049_ rbzero.tex_g0\[56\] rbzero.tex_g0\[55\] _11898_ _11902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25096__I _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22060_ rbzero.wall_tracer.rcp_fsm.o_data\[2\] rbzero.wall_tracer.stepDistY\[2\]
+ _03051_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__19634__A1 rbzero.wall_tracer.visualWallDist\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22513__I _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14740__B _07861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21011_ _02089_ _02099_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_151_Right_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16448__A1 rbzero.debug_overlay.vplaneY\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20244__A2 _11039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_206_Left_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_184_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_225_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25750_ _06495_ _06532_ _06533_ _06534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14031__I _07468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22962_ _03813_ _03819_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_5_13__f_i_clk_I clknet_3_3_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24701_ _05457_ _05484_ _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_241_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21913_ _02951_ _02952_ _02953_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_25681_ _06431_ _06464_ _06465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_223_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22893_ _02575_ _02684_ _03751_ _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_210_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_203_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27420_ _01325_ clknet_leaf_84_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__16620__A1 _10067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24632_ _05412_ _05414_ _05416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21844_ _02864_ _02875_ _02889_ _02859_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_33_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27351_ _01256_ clknet_leaf_98_i_clk rbzero.wall_tracer.trackDistX\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_215_Left_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24563_ _05264_ _05347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_148_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21775_ _10121_ _02825_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26302_ _00212_ clknet_leaf_215_i_clk rbzero.spi_registers.buf_otherx\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20726_ _12989_ _12585_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23514_ _04365_ _04300_ _04366_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_37_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15187__A1 _08959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27282_ _01187_ clknet_leaf_213_i_clk gpout0.hpos\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24494_ _05259_ _05276_ _05267_ _05274_ _05278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_163_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14915__B _08214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26233_ _00143_ clknet_leaf_1_i_clk rbzero.spi_registers.texadd2\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13737__A2 _07532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20657_ _01747_ _01748_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_23445_ _04284_ _04298_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_190_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23376_ _04193_ _04230_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_26164_ _00074_ clknet_leaf_184_i_clk rbzero.floor_leak\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24903__I _05298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20588_ _01610_ _01622_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_33_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25115_ _05895_ _05898_ _05899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22327_ _03281_ _03282_ _03252_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26095_ _00005_ clknet_leaf_225_i_clk rbzero.spi_registers.mosi_buffer\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24124__B _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13060_ gpout0.hpos\[3\] _06877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__19625__A1 _12206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22258_ _03201_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25046_ _05829_ _05830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_224_Left_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15746__B _09372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21209_ _01905_ _13012_ _02141_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_217_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22189_ _03162_ _03164_ _03168_ _03109_ rbzero.wall_tracer.rcp_fsm.i_data\[3\] _03169_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_100_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26997_ _00907_ clknet_leaf_172_i_clk rbzero.tex_g0\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__23185__A1 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23185__B2 _12428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16750_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] _10189_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25948_ _06727_ _06728_ _06700_ _06729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13962_ reg_rgb\[0\] _07186_ _07773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22932__A1 _12733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15701_ rbzero.spi_registers.buf_texadd2\[15\] _09340_ _09345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16681_ _10107_ _10124_ _10125_ _10126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_25879_ _05020_ _06662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_85_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13893_ rbzero.debug_overlay.playerY\[-2\] _07704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_214_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18420_ _11516_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_154_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15632_ rbzero.spi_registers.buf_texadd1\[21\] _09293_ _09294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_233_Left_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__24685__A1 _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18351_ _11476_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15563_ _09241_ _09242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17302_ rbzero.pov.spi_buffer\[29\] _10632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14514_ rbzero.tex_g0\[55\] _08317_ _08323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18282_ _11419_ _11406_ _11422_ _11423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_15494_ _09190_ _09191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_194_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17233_ rbzero.pov.spi_buffer\[12\] _10580_ _10577_ _10581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14925__A1 _08364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14445_ rbzero.tex_g0\[3\] _08252_ _08253_ _08254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17164_ rbzero.pov.spi_counter\[3\] _10527_ _10528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14376_ _07694_ _08058_ _08055_ _07687_ _08186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_133_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16678__A1 _10121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16115_ _09595_ _09655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_241_i_clk clknet_5_0__leaf_i_clk clknet_leaf_241_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13327_ _06879_ _07080_ _07141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__21671__A1 _11360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_242_Left_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_150_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17095_ rbzero.pov.ready_buffer\[19\] _10460_ _10476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16046_ _09515_ _09601_ _09605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15350__A1 rbzero.mapdxw\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13258_ _07070_ _07071_ _07072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21423__A1 _12777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16331__I _09818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13900__A2 _07704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13189_ _06991_ _07003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_237_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_166_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19805_ _12345_ _12577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17997_ rbzero.wall_tracer.trackDistX\[9\] _11141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_236_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19736_ _12506_ _12507_ _12508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24912__A2 _05296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16948_ _10295_ _10361_ _10362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_223_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_220_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16487__B _09942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19667_ _07705_ _12013_ _12254_ _12438_ _12439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_16879_ rbzero.pov.ready_buffer\[47\] _10252_ _10302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13690__I _07488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_144_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18618_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _11629_ _11630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19598_ _12356_ _12358_ _12361_ _12369_ _12370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_176_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18549_ _11590_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_220_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24209__B _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21560_ _02499_ _02515_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_47_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14735__B _08316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20511_ _01535_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13719__A2 _07506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_220_Right_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_173_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21491_ _02523_ _02556_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13275__S0 _07074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23230_ _03844_ _02075_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20442_ _12523_ _01535_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__21257__A4 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_209_i_clk clknet_5_7__leaf_i_clk clknet_leaf_209_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_23161_ _03909_ _03994_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_20373_ _12403_ _01466_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22112_ _03082_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23092_ _03947_ _03948_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14144__A2 _07919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_135_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17337__I _06897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22043_ rbzero.wall_tracer.rcp_fsm.o_data\[-4\] _03050_ _03051_ _03052_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__21414__A1 _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26920_ _00830_ clknet_leaf_130_i_clk rbzero.tex_r1\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_100_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17094__A1 _10474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26851_ _00761_ clknet_leaf_191_i_clk rbzero.tex_r0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_215_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_205_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_205_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25802_ _06581_ _06585_ _06586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_227_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26782_ _00692_ clknet_leaf_127_i_clk rbzero.tex_g1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23994_ rbzero.wall_tracer.rcp_fsm.operand\[6\] _04776_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21717__A2 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18043__B1 _11163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25733_ _06476_ _06504_ _06517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_22945_ _02621_ _03802_ _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_242_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22390__A2 _08182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25664_ _06403_ _06410_ _06447_ _06448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_195_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_238_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22876_ _02262_ _03734_ _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_238_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27403_ _01308_ clknet_leaf_111_i_clk rbzero.wall_tracer.stepDistX\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24615_ _05397_ _05398_ _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_168_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24131__A3 _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21827_ _02869_ _02871_ _02873_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_25595_ _06355_ _06353_ _06379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__18346__A1 _07179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24119__B _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27334_ _01239_ clknet_leaf_91_i_clk rbzero.trace_state\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_80_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24546_ _05329_ _05330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_183_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21758_ _09998_ _02809_ _02810_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20709_ _01711_ _01733_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27265_ _01170_ clknet_leaf_116_i_clk rbzero.wall_tracer.visualWallDist\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24477_ _05083_ _05261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14907__B2 _08558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21689_ _11260_ _12051_ _12024_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_0_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26216_ _00126_ clknet_leaf_10_i_clk rbzero.spi_registers.texadd1\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14230_ _08039_ _08040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_123_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23428_ _04178_ _04185_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_27196_ _01101_ clknet_leaf_75_i_clk rbzero.wall_tracer.size_full\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19846__B2 _12475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23642__A2 _12229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19727__I rbzero.wall_tracer.stepDistX\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14161_ _07257_ _07971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26147_ _00057_ clknet_leaf_214_i_clk rbzero.map_overlay.i_mapdx\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23359_ _04050_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13112_ rbzero.spi_registers.texadd3\[15\] _06922_ _06925_ rbzero.spi_registers.texadd2\[15\]
+ _06913_ _06926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_104_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26078_ _06662_ _06682_ _06692_ _06842_ _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_14092_ rbzero.tex_r1\[37\] _07901_ _07630_ _07902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_111_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17247__I _10555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25029_ _05545_ _05597_ _05813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_17920_ rbzero.wall_tracer.rayAddendX\[7\] _11064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13043_ _06858_ _06859_ _06860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_17851_ _10995_ _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__26500__D _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15990__I _09550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16802_ rbzero.pov.ready_buffer\[67\] _10228_ _10229_ _10234_ _10235_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_17782_ _10936_ _10952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_179_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14994_ net27 _08779_ _08781_ net19 _08796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_31_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19521_ rbzero.wall_tracer.size\[4\] _12181_ _12292_ _12252_ _12293_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_161_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16733_ _08908_ _10174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13945_ rbzero.map_overlay.i_mapdy\[3\] _07756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_233_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19452_ _12223_ _12224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_198_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16664_ _10108_ _10103_ _10109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13876_ rbzero.debug_overlay.playerX\[3\] _07687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_202_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15615_ _09258_ _09281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18403_ _11501_ _11507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_243_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19383_ net88 _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16595_ _10027_ _10005_ _10026_ _10044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18806__I _08752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18334_ _11464_ _11465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20144__A1 rbzero.wall_tracer.stepDistX\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15546_ _09190_ _09229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16899__A1 _08061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18265_ _11403_ _11406_ _11407_ _11408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_15477_ rbzero.spi_registers.buf_texadd0\[5\] _09178_ _09179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17216_ _10555_ _10568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14428_ _08232_ _08234_ _08236_ _08215_ _08222_ _08237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_71_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_180_i_clk clknet_5_8__leaf_i_clk clknet_leaf_180_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_18196_ rbzero.map_rom.b6 _11340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17147_ rbzero.pov.sclk_buffer\[2\] _09015_ _10514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__21644__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14359_ _07979_ _07202_ _08093_ _08168_ _08169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17078_ _08132_ _10463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_122_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16029_ rbzero.spi_registers.spi_buffer\[0\] _09591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_195_i_clk clknet_5_12__leaf_i_clk clknet_leaf_195_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_181_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_139_Left_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13885__B2 _07102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25138__A2 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_225_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19719_ _12490_ _12491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20991_ _01956_ _01604_ _02079_ _12790_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22730_ _11172_ _12511_ _03592_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_200_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20383__A1 _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25310__A2 _06093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22661_ _03532_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_133_i_clk clknet_5_15__leaf_i_clk clknet_leaf_133_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__18328__A1 _07205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24400_ _04719_ _05114_ _05023_ _05184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_148_Left_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21612_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_34_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25380_ _06162_ _06129_ _06163_ _06164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_clkbuf_leaf_61_i_clk_I clknet_5_21__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22592_ rbzero.side_hot _03475_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_192_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17000__A1 _10345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24331_ _05103_ _05113_ _05114_ _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_233_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21543_ _02624_ _02627_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__16236__I _09747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_233_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_148_i_clk clknet_5_11__leaf_i_clk clknet_leaf_148_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27050_ _00960_ clknet_leaf_121_i_clk rbzero.wall_tracer.mapY\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24262_ _05012_ _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_160_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21474_ _02459_ _02559_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_132_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26001_ _06645_ _06648_ _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20425_ _01416_ _01417_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21635__A1 _08128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23213_ _04068_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24193_ _04976_ _04977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_95_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23144_ _03768_ _03999_ _04000_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_20356_ _01447_ _01450_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13809__B _07587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__23388__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23075_ _03928_ _03931_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20287_ _01379_ _01381_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_140_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22026_ _03037_ _03039_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26903_ _00813_ clknet_leaf_125_i_clk rbzero.tex_r1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_41_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20610__A2 _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26834_ _00744_ clknet_leaf_199_i_clk rbzero.tex_r0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
Xhold43 net100 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_199_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21317__I _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26765_ _00675_ clknet_leaf_229_i_clk rbzero.spi_registers.sclk_buffer\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_242_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23977_ _04769_ _04771_ _04767_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_203_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22363__A2 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25716_ _06498_ _06499_ _06500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13730_ _07444_ _07541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_230_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22928_ _12791_ _01956_ _03669_ _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26696_ _00606_ clknet_leaf_67_i_clk rbzero.pov.ready_buffer\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16855__B _09028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25647_ _06383_ _06418_ _06430_ _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13661_ _07470_ _07471_ _07472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_168_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22859_ _03716_ _03717_ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_79_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15400_ rbzero.spi_registers.buf_sky\[2\] _09119_ _09123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17790__A2 rbzero.pov.ready_buffer\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16380_ _09855_ _09856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25578_ _06359_ _06360_ _06361_ _06362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13592_ _07077_ _07398_ _07393_ _06886_ _07403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_94_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27317_ _01222_ clknet_leaf_118_i_clk rbzero.traced_texa\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15331_ rbzero.map_overlay.i_mapdy\[1\] _09058_ _09071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24529_ _05244_ _05313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21874__A1 _10072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21874__B2 _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18050_ _11190_ _11191_ _11192_ _11193_ _11194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_108_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27248_ _01153_ clknet_leaf_77_i_clk rbzero.wall_tracer.rcp_fsm.i_start vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15262_ _09016_ _09017_ _09018_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19819__A1 _12160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17001_ _08079_ _10381_ _10405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14213_ _08022_ _08023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__21626__A1 _09900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15193_ _08965_ _08952_ _08966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27179_ _01084_ clknet_leaf_47_i_clk rbzero.wall_tracer.rayAddendX\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__18098__A3 _11227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14108__A2 _07916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14144_ rbzero.tex_r1\[58\] _07919_ _07953_ _07954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_238_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18952_ rbzero.tex_g0\[14\] rbzero.tex_g0\[13\] _11845_ _11847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14075_ _07841_ _07884_ _07885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23707__I _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17903_ rbzero.wall_tracer.rayAddendX\[0\] _11047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_18883_ rbzero.traced_texa\[3\] rbzero.texV\[3\] _11798_ _11800_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_238_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19192__I _12035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17834_ _10980_ rbzero.pov.ready_buffer\[70\] _10985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_128_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13619__A1 rbzero.floor_leak\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14977_ _08778_ net8 _08779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_88_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17765_ _10937_ rbzero.pov.ready_buffer\[45\] _10941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xrebuffer19 _05206_ net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_233_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23551__A1 _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19504_ _12275_ _12276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_50_i_clk clknet_5_17__leaf_i_clk clknet_leaf_50_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_107_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16716_ _10151_ _10156_ _10157_ _10158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13928_ _07736_ _06890_ _07738_ _07739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_159_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17696_ _10890_ rbzero.pov.ready_buffer\[22\] _10895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_141_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16647_ _10092_ _10093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19435_ _12204_ _11098_ _12205_ _12206_ _12207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_201_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13859_ _07430_ _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14044__A1 _07803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16578_ _10027_ _10005_ _10028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19366_ rbzero.tex_b1\[58\] rbzero.tex_b1\[57\] _12146_ _12148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_65_i_clk clknet_5_21__leaf_i_clk clknet_leaf_65_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_44_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18317_ _11450_ _11451_ _11452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15529_ _09190_ _09217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19297_ _12108_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_215_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__18581__I1 rbzero.tex_r0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18248_ rbzero.wall_tracer.rcp_fsm.i_start _11392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24273__I _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18179_ _11317_ _11319_ _11322_ _11323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_114_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20210_ _12902_ _12980_ _12981_ _12982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_52_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21190_ _02277_ _01474_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22290__A1 _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21093__A2 _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20141_ rbzero.wall_tracer.size\[9\] _12640_ _12912_ _12913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_204_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20072_ _12843_ _12844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_237_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23900_ _03017_ _04711_ _04712_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24880_ _05653_ _05654_ _05655_ _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__21137__I _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23831_ _03292_ _03072_ _04656_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_212_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_i_clk clknet_5_5__leaf_i_clk clknet_leaf_18_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__22345__A2 _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15135__I _08916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26550_ _00460_ clknet_leaf_66_i_clk rbzero.pov.spi_buffer\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23762_ _04568_ _04602_ _03590_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19210__A2 _12051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20974_ _02061_ _02062_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_156_Left_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25501_ _06282_ _06284_ _06285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_194_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_235_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22713_ _11190_ _12287_ _03577_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_221_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_194_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26481_ _00391_ clknet_leaf_57_i_clk rbzero.debug_overlay.facingX\[-8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23693_ _04535_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25432_ _06203_ _06209_ _06216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14907__C _08595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22644_ rbzero.wall_tracer.w\[2\] _03515_ _03517_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14586__A2 _07563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25363_ _06003_ _05973_ _06126_ _06145_ _06146_ _06147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_36_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22575_ _03467_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_97_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27102_ _01012_ clknet_leaf_138_i_clk rbzero.tex_b1\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24314_ _05033_ _05050_ _05055_ _05097_ _05098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_21526_ _02214_ _02489_ _02610_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_69_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25294_ _06027_ _06076_ _06077_ _06078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27033_ _00943_ clknet_leaf_137_i_clk rbzero.tex_g0\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24245_ _04844_ _04972_ _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_21457_ _02146_ _02377_ _02381_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_165_Left_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20408_ _12412_ _12562_ _12548_ _12298_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_21388_ _01947_ _01982_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24176_ _04860_ _04959_ _04960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_160_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23127_ _12961_ _03852_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput33 net33 o_hsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_20339_ rbzero.wall_tracer.stepDistX\[3\] _12280_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput44 net44 o_vsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_246_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_246_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23058_ _03913_ _03914_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15754__B _09384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14510__A2 _07617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14900_ rbzero.tex_b1\[51\] _07561_ _08706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22009_ rbzero.wall_tracer.size_full\[9\] _03020_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15880_ rbzero.spi_registers.buf_leak\[0\] _09476_ _09478_ _09479_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_216_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14831_ rbzero.tex_b1\[24\] _08518_ _08289_ _08637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26817_ _00727_ clknet_leaf_181_i_clk rbzero.tex_g1\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_208_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_174_Left_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_4_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17550_ _10803_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14762_ rbzero.tex_b0\[23\] _08568_ _08280_ _08569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26748_ _00658_ clknet_leaf_120_i_clk rbzero.wall_tracer.mapX\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_203_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19201__A2 _12044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16501_ rbzero.wall_tracer.rayAddendY\[-2\] _09956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_123_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13713_ _07442_ _07524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20898__A2 _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17481_ rbzero.tex_b0\[4\] rbzero.tex_b0\[3\] _10760_ _10764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14693_ rbzero.tex_b0\[53\] _07930_ _08500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__18356__I _11479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26679_ _00589_ clknet_leaf_23_i_clk rbzero.pov.ready_buffer\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__17763__A2 rbzero.pov.ready_buffer\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16432_ _08806_ _09892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19220_ rbzero.wall_tracer.mapY\[9\] _12061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_116_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13644_ rbzero.row_render.wall\[0\] _07454_ _07455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14577__A2 _07810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19151_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendY\[-2\] _11993_
+ _11994_ _11995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_109_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16363_ _08948_ _09842_ _09843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13575_ rbzero.row_render.size\[4\] _07372_ _07385_ _07386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_240_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18102_ _11144_ _11239_ _11244_ _11245_ _11246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_26_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15314_ _08878_ _09058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19082_ rbzero.debug_overlay.facingY\[-6\] _10030_ _11926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_136_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16294_ _09789_ _09790_ _09784_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_183_Left_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18033_ rbzero.wall_tracer.trackDistX\[-1\] _11177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_15245_ rbzero.spi_registers.spi_buffer\[22\] _08917_ _09007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25917__I _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15176_ _08951_ _08952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_151_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14127_ rbzero.tex_r1\[54\] _07641_ _07937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20822__A2 _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19984_ _12736_ _12738_ _12756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25210__A1 _05880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18935_ _11837_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14501__A2 _07600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14058_ _07526_ _07868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_123_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__23772__A1 _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18866_ _08753_ _11786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_192_Left_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_175_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17817_ _10972_ _10731_ _10968_ _10974_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_18797_ _11731_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_221_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20338__A1 rbzero.wall_tracer.stepDistY\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17748_ _10927_ _10661_ _10923_ _10929_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_221_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_234_i_clk_I clknet_5_3__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18266__I _11397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17679_ _08809_ _10884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__17754__A2 rbzero.pov.ready_buffer\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19418_ _12162_ _12189_ _12190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20690_ _01665_ _01779_ _01780_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_119_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19349_ _12138_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_230_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_230_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22360_ rbzero.mapdyw\[0\] _12038_ _03308_ _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_198_Right_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21311_ _02269_ _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22291_ _03201_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_245_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24252__A2 _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24030_ rbzero.wall_tracer.rcp_fsm.operand\[-4\] rbzero.wall_tracer.rcp_fsm.operand\[-5\]
+ rbzero.wall_tracer.rcp_fsm.operand\[-6\] rbzero.wall_tracer.rcp_fsm.operand\[-7\]
+ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_21242_ _02222_ _02241_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22263__A1 rbzero.wall_tracer.visualWallDist\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21173_ _12587_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_57_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_228_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20124_ _12495_ _12297_ _12896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25981_ _06757_ _06760_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23763__A1 _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20055_ _12826_ _12805_ _12827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24932_ _05713_ _05714_ _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__19431__A2 _12196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_241_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24863_ _05371_ _05493_ _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_225_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26602_ _00512_ clknet_leaf_38_i_clk rbzero.pov.spi_buffer\[71\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_213_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23814_ rbzero.wall_tracer.trackDistY\[5\] _03067_ _04642_ _04648_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24794_ _05531_ _05532_ _05578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26533_ _00443_ clknet_leaf_22_i_clk rbzero.pov.spi_buffer\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23745_ _04587_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__25268__A1 _06051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18176__I _11249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20957_ _01992_ _02024_ _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26464_ _00374_ clknet_leaf_206_i_clk rbzero.debug_overlay.playerX\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23676_ _04526_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20888_ _01976_ _01977_ _01525_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_193_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25415_ _06183_ _06192_ _06198_ _06199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_192_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22627_ _03505_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_101_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26395_ _00305_ clknet_leaf_19_i_clk rbzero.spi_registers.buf_texadd2\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25346_ _06115_ _06116_ _06129_ _06130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_180_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13360_ _07171_ _07158_ _07172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_192_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20501__A1 _12422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22558_ _11291_ _03455_ _03456_ rbzero.traced_texa\[2\] _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_134_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15749__B _09372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_165_Right_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21509_ _02340_ _02343_ _01944_ _01966_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_133_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25277_ _06043_ _06058_ _06061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16181__A1 _08968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13291_ rbzero.texu_hot\[0\] _06965_ _07105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_248_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22489_ _03415_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_248_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_248_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15030_ rbzero.spi_registers.spi_cmd\[3\] _08823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_27016_ _00926_ clknet_leaf_169_i_clk rbzero.tex_g0\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24228_ _04988_ _04989_ _04990_ _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_47_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_2__f_i_clk_I clknet_3_0_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24159_ _04920_ _04885_ _04901_ _04943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_20_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_183_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16981_ _08085_ _10381_ _10389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13298__A2 _07111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18720_ rbzero.tex_r1\[29\] rbzero.tex_r1\[28\] _11687_ _11688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15932_ rbzero.spi_registers.spi_buffer\[2\] _09518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13716__C _07526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15863_ _09462_ _09465_ _09466_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_18651_ _07171_ rbzero.tex_r0\[63\] _11644_ _11648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_203_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17602_ _10832_ _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14814_ _08371_ _08620_ _08621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18582_ _11609_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15794_ rbzero.spi_registers.buf_texadd3\[15\] _09409_ _09414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_231_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17533_ _10793_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14745_ _07888_ _08511_ _08524_ _08539_ _08551_ _08552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_169_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25259__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17464_ _10750_ _10746_ _10752_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14676_ _07801_ _08480_ _08483_ _08484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16415_ rbzero.spi_registers.buf_texadd3\[22\] _09874_ _09881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19203_ rbzero.wall_tracer.mapY\[6\] _12047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13627_ _07433_ _07436_ _07437_ _07438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17395_ _10699_ _10700_ _10701_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_229_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24037__B _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_212_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19134_ _11943_ _11978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_171_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16346_ rbzero.spi_registers.buf_texadd3\[4\] _09829_ _09830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13558_ _07039_ _07368_ _07369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18161__A2 _11260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19065_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _11908_ _11911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_136_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16334__I _09806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16277_ rbzero.spi_registers.buf_texadd2\[11\] _09769_ _09778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13489_ rbzero.texV\[3\] _07291_ _07300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_180_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18016_ rbzero.wall_tracer.trackDistX\[4\] _11160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__22245__A1 _12595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21048__A2 _12383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15228_ rbzero.spi_registers.spi_buffer\[17\] _08994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_140_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22796__A2 _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15159_ _08937_ _08929_ _08938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19967_ _12727_ _12736_ _12738_ _12739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_201_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24942__B1 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18918_ gpout2.clk_div\[0\] gpout2.clk_div\[1\] _11827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_19898_ _12665_ _12669_ _12670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_207_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18849_ _11767_ _11770_ _11771_ _11772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_207_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21860_ _11025_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14789__A2 _07930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15986__A1 _08977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19177__A1 _11269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21415__I _12684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20811_ _01793_ _01887_ _01900_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_132_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21791_ _08133_ _08139_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13461__A2 rbzero.spi_registers.vshift\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23530_ _04179_ _04382_ _04294_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_20742_ _12444_ _01720_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_159_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23461_ _04313_ _04314_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14029__I _07541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20673_ _01755_ _01764_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_161_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25200_ _05983_ _05984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_175_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22412_ _03355_ _03356_ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26180_ _00090_ clknet_leaf_188_i_clk rbzero.spi_registers.vshift\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__22484__A1 rbzero.wall_tracer.size\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23392_ rbzero.wall_tracer.stepDistX\[8\] _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25131_ _05236_ _05889_ _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22343_ _03274_ _03294_ _03295_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16163__A1 _08939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13089__B _06900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25062_ _05775_ _05780_ _05846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22274_ _03225_ _03236_ _03238_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14713__A2 _08291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19101__A1 rbzero.debug_overlay.facingY\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23984__A1 _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24013_ rbzero.wall_tracer.rcp_done _04722_ _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21225_ _02175_ _02310_ _02311_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_130_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_243_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_243_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21156_ _02145_ _02157_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14699__I _07566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23736__A1 _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14477__B2 _08284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20107_ _12632_ _12650_ _12878_ _12879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_208_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25964_ _06694_ _02994_ _06736_ _06744_ _06719_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_176_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21087_ _02047_ _02050_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20038_ _12666_ _12697_ _12810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24915_ _05329_ _05607_ _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25895_ _06676_ _06677_ _06678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_213_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24846_ _05626_ _05629_ _05630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14648__B _07946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_234_Right_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24777_ _05503_ _05507_ _05561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_69_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21989_ rbzero.wall_tracer.rcp_fsm.o_data\[2\] rbzero.wall_tracer.size\[10\] _03002_
+ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13452__A2 rbzero.spi_registers.vshift\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15323__I _09064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26516_ _00426_ clknet_leaf_60_i_clk rbzero.debug_overlay.vplaneY\[-6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14530_ _07489_ _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14367__C _07218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23728_ _04568_ _04572_ _03567_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_25_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26447_ _00357_ clknet_leaf_86_i_clk rbzero.wall_tracer.rayAddendY\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14461_ _07838_ _08268_ _08269_ _08270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_166_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23659_ _04469_ _04510_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_166_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16200_ rbzero.spi_registers.buf_texadd1\[16\] _09719_ _09720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13412_ _07195_ _07206_ _07222_ _07223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_181_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17180_ rbzero.pov.mosi _10539_ _10540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_165_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26378_ _00288_ clknet_leaf_250_i_clk rbzero.spi_registers.buf_texadd1\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14392_ _07928_ _08201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_153_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14952__A2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13778__I _07449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16131_ _09667_ _09657_ _09668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25329_ _06111_ _06112_ _06113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13343_ net14 _07155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25413__A1 _05605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19891__A2 _12192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__26072__B _09113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22227__A1 _11392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16062_ _09542_ _09612_ _09617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14704__A2 _08503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13274_ _06979_ _06982_ _07088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__25964__A2 _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15013_ rbzero.wall_tracer.rcp_fsm.i_start rbzero.wall_tracer.rcp_fsm.state\[0\]
+ _08812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19465__I _12236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15993__I _09564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19821_ _12592_ _12593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_120_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19752_ _12522_ _12523_ _12524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14402__I _07946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16964_ _10374_ _10375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13446__C _07256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18703_ _11678_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_34_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15915_ _09502_ _09503_ _09505_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19683_ _12436_ _12453_ _12455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_16895_ rbzero.debug_overlay.playerY\[-5\] _10303_ _10316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_232_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_189_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18634_ _11638_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15846_ rbzero.spi_registers.buf_sky\[4\] _09439_ _09453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_189_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14558__B _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24152__A1 _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_201_Right_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18565_ _11599_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15777_ _09400_ _09401_ _09395_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__18906__A1 rbzero.traced_texa\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17516_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _10781_ _10784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14728_ rbzero.tex_b0\[47\] _08241_ _07867_ _08535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18496_ rbzero.tex_g1\[61\] rbzero.tex_g1\[60\] _11559_ _11560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14659_ rbzero.tex_g1\[54\] _07641_ _08467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17447_ _10705_ _10740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17378_ rbzero.pov.spi_buffer\[49\] _10685_ _10682_ _10689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13688__I _07498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19117_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] _11961_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_144_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16145__A1 _08913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16329_ rbzero.spi_registers.buf_texadd3\[0\] _09816_ _09817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__26564__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19048_ _11901_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22769__A2 rbzero.wall_tracer.stepDistX\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19634__A2 _11381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_120_Left_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_54_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21010_ _12836_ _02098_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__18693__I0 rbzero.tex_r1\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22961_ _03816_ _03818_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24700_ _05460_ _05463_ _05483_ _05484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__17623__I _10844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21912_ _02941_ _02947_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25680_ _06434_ _06463_ _06464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22892_ _02574_ _02685_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_179_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_203_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21145__I _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24631_ _05412_ _05414_ _05415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21843_ _08121_ _11075_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_222_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27350_ _01255_ clknet_leaf_90_i_clk rbzero.wall_tracer.trackDistX\[-8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_195_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24562_ _05325_ _05341_ _05346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_38_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_131_i_clk_I clknet_5_14__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21774_ _10471_ _12216_ _02824_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_33_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26301_ _00211_ clknet_leaf_215_i_clk rbzero.spi_registers.buf_otherx\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23513_ _04271_ _04279_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20725_ _01693_ _01694_ _01815_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27281_ _01186_ clknet_leaf_213_i_clk gpout0.hpos\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24493_ _05259_ _05267_ _05274_ _05276_ _05277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_65_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26232_ _00142_ clknet_leaf_1_i_clk rbzero.spi_registers.texadd1\[23\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23444_ _04289_ _04291_ _04297_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_147_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20656_ _12658_ _01478_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26163_ _00073_ clknet_leaf_184_i_clk rbzero.floor_leak\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23375_ _04197_ _04229_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_162_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20587_ _01584_ _01677_ _01678_ _01625_ _01582_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_162_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25114_ _05896_ _05897_ _05898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_61_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17884__A1 rbzero.debug_overlay.facingX\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22326_ _11284_ _03250_ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26094_ _06855_ _06856_ _08811_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14931__B _08198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25045_ _05770_ _05798_ _05829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22257_ _03202_ _03223_ _03224_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13370__A1 _07179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21208_ _02135_ _02140_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13370__B2 _07180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22188_ _03165_ _03167_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_56_i_clk_I clknet_5_23__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21139_ _12779_ _01484_ _01924_ _01925_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_26996_ _00906_ clknet_leaf_172_i_clk rbzero.tex_g0\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__24382__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13961_ _07232_ _07771_ _07772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__15762__B _09384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25947_ _06676_ _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_233_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14870__A1 _08295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15700_ rbzero.spi_registers.texadd2\[15\] _09338_ _09344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_216_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16680_ _10086_ _10125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_25878_ _06903_ _02980_ _06658_ _06661_ _10992_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_13892_ _07191_ _07698_ _07700_ _07041_ _07702_ _07703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_214_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21991__I0 rbzero.wall_tracer.rcp_fsm.o_data\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24829_ _05418_ _05310_ _05613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_15631_ _09258_ _09293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_198_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18350_ _11474_ rbzero.spi_registers.sclk_buffer\[0\] _11476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15562_ _09240_ _09241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17301_ _10629_ _10630_ _10631_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15988__I _09547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14513_ rbzero.tex_g0\[54\] _07872_ _08322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15493_ _08986_ _09190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18281_ rbzero.wall_tracer.mapX\[8\] _11420_ _11421_ _11422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14444_ rbzero.tex_g0\[2\] _08206_ _08253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17232_ _10555_ _10580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17163_ _10512_ _10526_ _10527_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_36_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14375_ _07677_ _08053_ _08026_ _08184_ _08185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__21120__A1 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16114_ _09653_ _09654_ _09648_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13326_ _07107_ _07118_ _07138_ _07063_ _07139_ _07140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_134_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17094_ _10474_ _10458_ _10475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16045_ rbzero.spi_registers.buf_texadd0\[1\] _09597_ _09604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13257_ _06906_ _07002_ _07071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13361__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13188_ _06996_ _07001_ _07002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19804_ _12248_ _11985_ _12576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_224_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17996_ rbzero.wall_tracer.trackDistX\[10\] _11140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__24373__A1 _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19735_ _12384_ _12388_ _12507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16947_ _10359_ _10353_ _10361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_220_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19666_ _11952_ _11998_ _10323_ _12003_ _12438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_16878_ _10282_ _10301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_205_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18617_ _11628_ _11629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15829_ rbzero.spi_registers.buf_sky\[0\] _09439_ _09440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16059__I _09614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19597_ _12368_ _12369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_231_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22687__A1 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18548_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _11587_ _11590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24276__I _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20162__A2 _12667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18479_ _11550_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20510_ _01587_ _01602_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14916__A2 _08226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21490_ _02457_ _02562_ _02560_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_16_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13275__S1 _07053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20441_ _01534_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19855__A2 _12382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16950__C _09441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23160_ _03904_ _03907_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_125_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20372_ _01376_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22524__I _09938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22111_ _03079_ _03103_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23091_ _02271_ _02115_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22042_ _03038_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20044__I _12788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26850_ _00760_ clknet_leaf_192_i_clk rbzero.tex_r0\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_205_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25801_ _06582_ _06584_ _06585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_177_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16841__A2 _07687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26781_ _00691_ clknet_leaf_127_i_clk rbzero.tex_g1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23993_ _04782_ _04783_ _04767_ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_242_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25732_ _06476_ _06504_ _06516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_173_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22944_ _03661_ _03662_ _03801_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_98_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19791__A1 _12476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25663_ _06406_ _06409_ _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22875_ _02546_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14604__A1 rbzero.tex_g1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_238_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_238_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27402_ _01307_ clknet_leaf_109_i_clk rbzero.wall_tracer.stepDistX\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24614_ _05363_ _05356_ _05386_ _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_168_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_5__f_i_clk clknet_3_1_0_i_clk clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21826_ _02872_ _02857_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25594_ _06355_ _06353_ _06378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27333_ _01238_ clknet_leaf_35_i_clk rbzero.side_hot vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24545_ _05328_ _05329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21757_ rbzero.wall_tracer.rayAddendX\[-4\] _02722_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24419__A2 _05202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20708_ _01714_ _01732_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27264_ _01169_ clknet_leaf_116_i_clk rbzero.wall_tracer.visualWallDist\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24476_ _05213_ _05260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_21688_ _02750_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_163_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26215_ _00125_ clknet_leaf_16_i_clk rbzero.spi_registers.texadd1\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23427_ _04178_ _04185_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_27195_ _01100_ clknet_leaf_74_i_clk rbzero.wall_tracer.size\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_20639_ _01727_ _01730_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_191_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23642__A3 _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14160_ _07431_ _07965_ _07969_ _07970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26146_ _00056_ clknet_leaf_216_i_clk rbzero.map_overlay.i_mapdx\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13591__A1 _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23358_ _04053_ _04055_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__21653__A2 _08194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13111_ _06924_ _06925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_22309_ rbzero.wall_tracer.trackDistY\[1\] _03243_ _03244_ _03267_ _03268_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_132_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26077_ _06660_ _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14091_ _07459_ _07901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23289_ _04033_ _04046_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25028_ _05809_ _05810_ _05811_ _05812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_30_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13042_ gpout0.hpos\[9\] _06859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XTAP_TAPCELL_ROW_111_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17850_ _09892_ rbzero.pov.mosi_buffer\[0\] _10995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24355__A1 _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16801_ _10171_ _10232_ _10233_ _10234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17781_ _10934_ _10951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14993_ _07171_ _08782_ _08795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26979_ _00889_ clknet_leaf_123_i_clk rbzero.texV\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__17263__I _10602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19520_ _12289_ _11989_ _12290_ _12291_ _12292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_31_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16732_ rbzero.pov.ready_buffer\[59\] _10169_ _10172_ _10173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_161_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13944_ _07214_ _07753_ _07754_ _07755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__24297__S _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19782__A1 _12553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19782__B2 _12401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19451_ _12222_ _12223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16663_ _10099_ _10100_ _10108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13875_ _07197_ _07686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__20392__A2 _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18402_ _11506_ _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15614_ rbzero.spi_registers.texadd1\[17\] _09279_ _09280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19382_ _11474_ net87 _12156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_202_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16594_ _10041_ _10042_ _10043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_243_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14836__B _07826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18333_ _07220_ _11460_ _11464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15545_ rbzero.spi_registers.buf_texadd1\[0\] _09220_ _09228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16348__A1 _08926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14359__B1 _08093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15476_ _09153_ _09178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18264_ rbzero.wall_tracer.mapX\[6\] _11404_ _11128_ _11407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_13_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__19918__I _12501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14427_ rbzero.tex_g0\[19\] _08210_ _08235_ _08236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17215_ rbzero.pov.spi_buffer\[7\] _10567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__23094__A1 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18195_ _11304_ _11336_ _11338_ _11339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17146_ rbzero.pov.spi_counter\[0\] _10513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14358_ _08089_ _08147_ _08167_ _08168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_52_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13309_ rbzero.spi_registers.texadd0\[2\] _07123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17077_ _10459_ _10461_ _10462_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14289_ _08098_ _08099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_21_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13334__A1 _07060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16028_ rbzero.spi_registers.buf_mapdyw\[0\] _09583_ _09590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13885__A2 _07693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17979_ _11108_ _11122_ _11123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14834__B2 _08294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19718_ _12337_ _12339_ _12342_ _12490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_79_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20990_ _02078_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__20907__A1 _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19773__A1 _12468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19649_ _12420_ _12421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_200_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16587__B2 _10036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22660_ _03531_ rbzero.wall_tracer.trackDistX\[-10\] _11400_ _03532_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21611_ _08933_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_22591_ _07028_ _03475_ _03478_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_62_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24330_ _05010_ _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_192_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21542_ _02625_ _02626_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_8_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_233_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_99_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24261_ _05044_ _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_145_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21473_ _02519_ _02558_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_26000_ _06747_ _06708_ _06778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23212_ _04063_ _04067_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20424_ _01516_ _01438_ _01517_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24192_ _04933_ _04973_ _04974_ _04975_ _04976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA__22832__A1 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14481__B _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23143_ _03998_ _03881_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20355_ _12952_ _01448_ _01449_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_229_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23074_ _03667_ _03930_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_20286_ _12816_ _12960_ _01380_ _12750_ _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22025_ _03038_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26902_ _00812_ clknet_leaf_132_i_clk rbzero.tex_r1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_228_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_216_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20071__A1 _12841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26833_ _00743_ clknet_leaf_199_i_clk rbzero.tex_r0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
Xhold44 _12156_ net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_243_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23976_ rbzero.wall_tracer.rcp_fsm.i_data\[1\] _04770_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26764_ _00674_ clknet_leaf_230_i_clk rbzero.spi_registers.sclk_buffer\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_231_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25715_ _06451_ _06457_ _06499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_22927_ _03650_ _03783_ _03784_ _03659_ _03664_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_26695_ _00605_ clknet_leaf_67_i_clk rbzero.pov.ready_buffer\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20374__A2 _12199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_240_i_clk clknet_5_1__leaf_i_clk clknet_leaf_240_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13660_ rbzero.row_render.texu\[4\] _07452_ _07417_ _07451_ _07471_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_25646_ _06428_ _06416_ _06365_ _06429_ _06430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_196_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22858_ _01996_ _01953_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21809_ _02852_ _02855_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_25577_ _05977_ _06013_ _06361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13591_ _07062_ _07397_ _07398_ _06885_ _07401_ _07402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_22789_ _02599_ _02604_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__21323__A1 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13800__A2 _07460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15330_ _09069_ _09070_ _09055_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24528_ _05310_ _05311_ _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27316_ _01221_ clknet_leaf_94_i_clk rbzero.traced_texa\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15261_ _08987_ _09018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24459_ _05242_ _05003_ _05025_ _05054_ _05243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_27247_ _01152_ clknet_leaf_81_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15553__A2 _09230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17000_ _10345_ _10402_ _10404_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14212_ _07998_ _08021_ _08022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_27178_ _01083_ clknet_leaf_48_i_clk rbzero.wall_tracer.rayAddendX\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15192_ rbzero.spi_registers.spi_buffer\[10\] _08965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14391__B _08198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13786__I _07576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17258__I _10564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14143_ rbzero.tex_r1\[59\] _07583_ _07953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_26129_ _00039_ clknet_leaf_250_i_clk rbzero.spi_registers.spi_buffer\[21\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18951_ _11846_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14074_ _07868_ _07880_ _07883_ _07884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_120_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17902_ rbzero.debug_overlay.facingX\[-7\] _11014_ _11046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_120_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_163_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18882_ rbzero.traced_texa\[4\] rbzero.texV\[4\] _11799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__24328__A1 _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24328__B2 _05111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17833_ _10979_ _10748_ _10982_ _10984_ _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_128_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13619__A2 _07326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17764_ _10935_ _10676_ _10939_ _10940_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_16_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14976_ net9 _08778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19503_ _12274_ _12275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23723__I _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16715_ _10145_ _10136_ _09934_ _10067_ _10157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_13927_ _07737_ _07373_ _06890_ _07736_ _07738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_208_i_clk clknet_5_7__leaf_i_clk clknet_leaf_208_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__21562__A1 _12238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17695_ _10889_ _10608_ _10892_ _10894_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_18_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19434_ _11387_ _12206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_186_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_179_Right_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16646_ _08095_ _10092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13858_ _07668_ _07669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__19507__A1 _08048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19365_ _12147_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16577_ _08112_ _08098_ _10002_ _10027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_clkbuf_leaf_178_i_clk_I clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13789_ _07599_ _07600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__23854__A3 _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18316_ _11433_ _07181_ _07712_ _11451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15528_ rbzero.spi_registers.buf_texadd0\[19\] _09209_ _09216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_44_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19296_ rbzero.tex_b1\[28\] rbzero.tex_b1\[27\] _12104_ _12108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_215_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18247_ _11390_ _11391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15459_ _09164_ _09166_ _09162_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_199_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18178_ rbzero.map_overlay.i_otherx\[3\] _11320_ _11106_ _09027_ _11321_ _11322_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_41_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13696__I _07479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17129_ rbzero.pov.ready_buffer\[5\] _10379_ _10502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_230_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20140_ _12247_ _12912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20071_ _12841_ _12817_ _12842_ _12843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14807__A1 _07802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23830_ _03292_ _03072_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23761_ _04598_ _03058_ _04601_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20973_ _01943_ _01960_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25819__A1 _05951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17631__I _10844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_23__f_i_clk clknet_3_5_0_i_clk clknet_5_23__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25500_ _06110_ _06117_ _06283_ _06284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_22712_ _11225_ rbzero.wall_tracer.stepDistX\[-4\] _03572_ _03577_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_194_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26480_ _00390_ clknet_leaf_58_i_clk rbzero.debug_overlay.facingX\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_235_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23692_ _11210_ _04529_ _04541_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_146_Right_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25431_ _06201_ _06210_ _06213_ _06215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_138_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22643_ rbzero.wall_tracer.w\[1\] _03508_ _03512_ rbzero.wall_tracer.w\[2\] _03517_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_137_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25362_ _06085_ _06086_ _06125_ _06009_ _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_22574_ _11278_ _09974_ _01553_ rbzero.traced_texa\[9\] _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__18182__B1 _11106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24313_ _05074_ _05084_ _05087_ _05096_ _05097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_152_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27101_ _01011_ clknet_leaf_138_i_clk rbzero.tex_b1\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_21525_ _12837_ _02489_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25293_ _06020_ _05974_ _06022_ _06077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_90_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16732__A1 rbzero.pov.ready_buffer\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27032_ _00942_ clknet_leaf_134_i_clk rbzero.tex_g0\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24244_ _05027_ _05028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21456_ _02425_ _02426_ _02541_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20407_ _12562_ _12548_ _12297_ _12412_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_121_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24175_ _04761_ _04856_ _04959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_21387_ _01951_ _01845_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23126_ _03816_ _03818_ _03982_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_31_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20338_ rbzero.wall_tracer.stepDistY\[3\] _12906_ _01429_ _01432_ _01433_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xoutput34 net34 o_rgb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_246_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23057_ _03799_ _03804_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23230__A1 _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20269_ _13037_ _13039_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_101_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22008_ rbzero.wall_tracer.rcp_fsm.o_data\[9\] _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_216_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15326__I _09067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26816_ _00726_ clknet_leaf_180_i_clk rbzero.tex_g1\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14830_ rbzero.tex_b1\[25\] _08252_ _08636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_231_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14761_ _07835_ _08568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26747_ _00657_ clknet_leaf_119_i_clk rbzero.wall_tracer.mapX\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_230_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23959_ rbzero.wall_tracer.rcp_fsm.operand\[-2\] _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16500_ _09924_ _09954_ _09955_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_123_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13712_ _07340_ _07523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22159__I _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17480_ _10763_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14692_ _07535_ _08499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26678_ _00588_ clknet_leaf_23_i_clk rbzero.pov.ready_buffer\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_224_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14026__A2 _07835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_224_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16431_ _08841_ _09886_ _09891_ _08888_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_25629_ _06025_ _05970_ _06412_ _06413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__16157__I _09660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13643_ _07417_ _07448_ _07449_ _07451_ _07453_ _07454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xclkbuf_leaf_194_i_clk clknet_5_12__leaf_i_clk clknet_leaf_194_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19150_ _08160_ _09965_ _11994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_16362_ _09819_ _09842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13574_ rbzero.row_render.size\[2\] rbzero.row_render.size\[1\] rbzero.row_render.size\[0\]
+ _07385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_54_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18173__B1 _11251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18101_ _11159_ _11231_ _11245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15313_ _09056_ _09031_ _09057_ _09036_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_19081_ _11923_ _11924_ _11925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16293_ rbzero.spi_registers.spi_buffer\[15\] _09782_ _09790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18032_ _11173_ rbzero.wall_tracer.trackDistY\[-2\] _11174_ _11175_ _11176_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15244_ _09004_ _09006_ _09003_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15175_ _08905_ _08951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__17523__I0 rbzero.tex_b0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14405__I _07448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14126_ _07929_ _07931_ _07934_ _07912_ _07935_ _07936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_104_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19983_ _12736_ _12738_ _12755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18321__B _10256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_132_i_clk clknet_5_15__leaf_i_clk clknet_leaf_132_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__18228__A1 rbzero.map_overlay.i_mapdx\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18934_ rbzero.tex_g0\[6\] rbzero.tex_g0\[5\] _11835_ _11837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14057_ _07501_ _07867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_238_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_248_Right_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_207_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_207_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18865_ _11779_ _11784_ _11785_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_207_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19028__I0 rbzero.tex_g0\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17816_ _10973_ rbzero.pov.ready_buffer\[63\] _10974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_238_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18796_ rbzero.tex_r1\[62\] rbzero.tex_r1\[61\] _11729_ _11731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_147_i_clk clknet_5_11__leaf_i_clk clknet_leaf_147_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__19728__A1 _12499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24721__A1 _05257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17747_ _10928_ rbzero.pov.ready_buffer\[39\] _10929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20338__A2 _12906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14959_ _07074_ _08749_ _08756_ _07153_ _08762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__17451__I _10543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17678_ _10881_ _10590_ _10877_ _10883_ _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_217_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19417_ rbzero.wall_tracer.stepDistY\[-11\] _12169_ _12188_ _12189_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_9_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16629_ _10038_ _10063_ _08095_ _10076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16962__A1 _08881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19348_ rbzero.tex_b1\[50\] rbzero.tex_b1\[49\] _12136_ _12138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24284__I _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_230_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_230_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19279_ _12098_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_245_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13528__A1 _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21310_ _02331_ _02396_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__24788__A1 _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22290_ _03247_ _03251_ _03252_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21241_ _02183_ _02184_ _02221_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_170_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_92_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21172_ _01483_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_57_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17626__I rbzero.pov.spi_done vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20123_ _12568_ _12380_ _12895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_228_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25980_ _06758_ rbzero.wall_tracer.rcp_fsm.o_data\[-7\] _06759_ _06760_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_217_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_215_Right_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20054_ _12799_ _12804_ _12826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24931_ _05713_ _05714_ _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_237_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__21774__A1 _10471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24862_ _05315_ _05645_ _05312_ _05646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_241_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26601_ _00511_ clknet_leaf_38_i_clk rbzero.pov.spi_buffer\[70\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23813_ _03283_ _03067_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24793_ _05560_ _05566_ _05576_ _05577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_139_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23744_ _11174_ _04585_ _04586_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14918__C _08334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26532_ _00442_ clknet_leaf_28_i_clk rbzero.pov.spi_buffer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20956_ _01909_ _02043_ _02044_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_49_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23675_ _12042_ _12043_ _04525_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_26463_ _00373_ clknet_leaf_208_i_clk rbzero.debug_overlay.playerX\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_20887_ rbzero.wall_tracer.size_full\[8\] _01975_ _01528_ _01977_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16953__A1 _07685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25414_ _06193_ _06196_ _06197_ _06198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_76_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22626_ rbzero.wall_tracer.texu\[3\] rbzero.texu_hot\[3\] _03503_ _03505_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_26394_ _00304_ clknet_leaf_18_i_clk rbzero.spi_registers.buf_texadd2\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_192_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21611__I _08933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25345_ _06119_ _06122_ _06128_ _06129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_9_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22557_ _03457_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21508_ _02071_ _02481_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25276_ _06059_ _06060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_20_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13290_ _06966_ _06967_ _07104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_248_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22488_ rbzero.wall_tracer.size\[2\] _03410_ _03412_ _07365_ _03415_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_248_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_248_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24227_ _05010_ _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_161_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27015_ _00925_ clknet_leaf_149_i_clk rbzero.tex_g0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14192__A1 _07212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21439_ _12238_ _02524_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18920__I _10757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24158_ _04941_ _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17130__A1 _06900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15765__B _09384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_219_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_126_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23109_ _03848_ _03854_ _03850_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_9_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24089_ _04852_ _04872_ _04873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_16980_ _10387_ _10388_ _10386_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_9_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15931_ rbzero.spi_registers.buf_othery\[2\] _09510_ _09517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_64_i_clk clknet_5_21__leaf_i_clk clknet_leaf_64_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_18650_ _11647_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_216_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15862_ _08920_ _09460_ _09466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17601_ rbzero.tex_b0\[56\] rbzero.tex_b0\[55\] _10828_ _10832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14813_ _07431_ _08493_ _08619_ _08620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_192_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18581_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _11608_ _11609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_188_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15793_ rbzero.spi_registers.texadd3\[15\] _09407_ _09413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_24_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_192_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_79_i_clk clknet_5_30__leaf_i_clk clknet_leaf_79_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17532_ rbzero.tex_b0\[26\] rbzero.tex_b0\[25\] _10791_ _10793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14744_ _08264_ _08545_ _08550_ _08355_ _08551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_197_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17463_ rbzero.pov.spi_buffer\[71\] _10743_ _10751_ _10752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_196_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15747__A2 _09373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14675_ _07475_ _08481_ _08482_ _07437_ _08483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_50_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19202_ _12044_ _12046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16414_ _09879_ _09880_ _09878_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13626_ net18 _07437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17394_ rbzero.pov.spi_buffer\[53\] _10697_ _10693_ _10701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19133_ _11957_ _11975_ _11976_ _11977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18316__B _07712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_212_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16345_ _09815_ _09829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_171_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23690__A1 _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13557_ _07367_ _07056_ _07368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18161__A3 _11251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19064_ _11910_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16276_ _09776_ _09777_ _09773_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13488_ _07296_ _07297_ _07298_ _07299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_164_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18015_ _11154_ _11158_ _11159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15227_ rbzero.spi_registers.spi_buffer\[18\] _08992_ _08993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_17_i_clk clknet_5_5__leaf_i_clk clknet_leaf_17_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_160_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15158_ rbzero.spi_registers.spi_buffer\[4\] _08937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_239_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25195__A1 _05977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14109_ _07523_ _07919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_19966_ _12737_ _12738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15089_ _07790_ _08872_ _08873_ _08874_ _08881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_239_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19949__A1 _12426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18917_ gpout2.clk_div\[0\] _11826_ _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19897_ _12667_ _12668_ _12669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_38_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21756__A1 _09927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19661__I _12432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18848_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] _11771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__21508__A1 _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18779_ _11721_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14738__C _08245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20810_ _01796_ _01886_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_21790_ _02833_ _02835_ _02839_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22181__A1 _12005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20741_ _01702_ _01706_ _01703_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_187_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16935__A1 rbzero.pov.ready_buffer\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23460_ _04199_ _04080_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20672_ _01637_ _01763_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14754__B _07955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22411_ _03326_ _03339_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23391_ rbzero.wall_tracer.trackDistX\[8\] _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23681__A1 _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25130_ _05893_ _05900_ _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22342_ _11281_ _03290_ _03278_ _03295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25422__A2 _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25061_ _05839_ _05844_ _05845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22273_ rbzero.wall_tracer.visualWallDist\[-5\] _03237_ _03229_ _03238_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14045__I _07599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20247__A1 rbzero.wall_tracer.size\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24012_ _04796_ _08814_ _04797_ _11473_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_41_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21224_ _02178_ _02301_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22262__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_243_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21155_ _02182_ _02242_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_243_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20106_ _12617_ _12631_ _12878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25963_ _06738_ _06741_ _06743_ _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_208_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21086_ _02041_ _02172_ _02173_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19571__I _12342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24410__C _05163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20037_ _12780_ _12686_ _12809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24914_ _05419_ _05695_ _05697_ _05698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_25894_ _06649_ _06646_ _06677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_225_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_213_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24845_ _05627_ _05629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__18187__I rbzero.map_rom.f4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24161__A2 _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17179__A1 rbzero.pov.ss_buffer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21988_ _03013_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_24776_ _05508_ _05517_ _05559_ _05560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26515_ _00425_ clknet_leaf_31_i_clk rbzero.debug_overlay.vplaneY\[-7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_23727_ _11221_ _03048_ _04571_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20939_ _01899_ _01901_ _02028_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_25_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18915__I _07167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_26446_ _00356_ clknet_leaf_86_i_clk rbzero.wall_tracer.rayAddendY\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_52_i_clk_I clknet_5_23__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14460_ rbzero.tex_g0\[10\] _07816_ _08269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23042__B _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23658_ _04500_ _04503_ _04509_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_36_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13411_ net3 _07212_ _07215_ _07221_ _07222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_22609_ _03490_ _03492_ _03494_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14391_ _08197_ _07669_ _08198_ _08199_ _08200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_23589_ _04255_ _04341_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_153_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26377_ _00287_ clknet_leaf_248_i_clk rbzero.spi_registers.buf_texadd1\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16130_ rbzero.spi_registers.spi_buffer\[23\] _09667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13342_ net13 net12 _07154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_25328_ _06050_ _06046_ _06112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16061_ rbzero.spi_registers.buf_texadd0\[5\] _09610_ _09616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13273_ _06989_ _07086_ _07087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25259_ _06031_ _06033_ _06042_ _06043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13912__A1 _07720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15012_ _08810_ _08811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__22172__I _10151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13912__B2 _07678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21986__A1 _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19820_ _08181_ _12160_ _12591_ _12592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_209_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16170__I _09675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18851__A1 _11769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_236_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19751_ _12302_ _12523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23727__A2 _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16963_ _10373_ _10374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21738__A1 _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18702_ rbzero.tex_r1\[21\] rbzero.tex_r1\[20\] _11677_ _11678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15914_ _09504_ _09505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_235_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19682_ _12436_ _12453_ _12454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_194_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16894_ rbzero.pov.ready_buffer\[49\] _10252_ _10315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_204_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18633_ rbzero.tex_r0\[56\] rbzero.tex_r0\[55\] _11634_ _11638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_204_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15845_ _09451_ _09452_ _09448_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_204_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18564_ rbzero.tex_r0\[26\] rbzero.tex_r0\[25\] _11597_ _11599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15776_ rbzero.spi_registers.buf_texadd3\[10\] _09398_ _09401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17515_ _10783_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14727_ rbzero.tex_b0\[46\] _08248_ _08534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18825__I _11737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18495_ _11543_ _11559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16917__A1 _07704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24048__B _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17446_ rbzero.pov.spi_buffer\[66\] _10739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_129_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22347__I _09926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14658_ _07841_ _08460_ _08465_ _08466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_145_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13609_ _07419_ _07420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16345__I _09815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17377_ _10665_ _10688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_171_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14589_ rbzero.tex_g1\[29\] _07845_ _08397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19116_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] _11960_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16328_ _09815_ _09816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19656__I _12414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19047_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _11898_ _11901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_180_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16259_ rbzero.spi_registers.buf_texadd2\[6\] _09757_ _09765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13903__A1 _07712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19095__A1 rbzero.debug_overlay.facingY\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25168__A1 _05951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17645__A2 rbzero.pov.ready_buffer\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18693__I1 rbzero.tex_r1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14459__A2 _07626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19949_ _12426_ _12414_ _12721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_149_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21729__A1 _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24391__A2 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22960_ _02540_ _03817_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21911_ rbzero.wall_tracer.rayAddendX\[8\] _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_241_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22891_ _03632_ _03633_ _03749_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__15424__I _09139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24143__A2 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_203_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24630_ _05351_ _05413_ _05354_ _05414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_21842_ _08121_ _11020_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_139_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14631__A2 _07901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25891__A2 _06652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24561_ _05342_ _05344_ _05345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_33_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16908__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21773_ _02817_ _02822_ _02823_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_194_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26300_ _00210_ clknet_leaf_217_i_clk rbzero.spi_registers.buf_otherx\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20724_ _12424_ _12646_ _01695_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_23512_ _04280_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_93_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6_0_i_clk clknet_0_i_clk clknet_3_6_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_24492_ _05275_ _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_147_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27280_ _01185_ clknet_leaf_214_i_clk gpout0.hpos\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21161__I _12237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25643__A2 _06382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26231_ _00141_ clknet_leaf_1_i_clk rbzero.spi_registers.texadd1\[22\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23443_ _04293_ _04296_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20655_ _12929_ _12489_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23374_ _04208_ _04228_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_144_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26162_ _00072_ clknet_leaf_184_i_clk rbzero.floor_leak\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20586_ _01603_ _01624_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19566__I _12337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25113_ _05492_ _05333_ _05336_ _05385_ _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_22325_ _11162_ _03206_ _03244_ _03280_ _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_150_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14147__A1 _07555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26093_ _06823_ _06660_ _06827_ _06856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__22209__A2 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24405__C _05163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14698__A2 _08496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25044_ _05763_ _05766_ _05828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22256_ rbzero.wall_tracer.visualWallDist\[-8\] _03218_ _03211_ _03224_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19086__A1 _08157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21207_ _02131_ _02160_ _02294_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_113_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22187_ _11290_ _03166_ _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_245_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__23709__A2 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21138_ _12684_ _01578_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26995_ _00905_ clknet_leaf_172_i_clk rbzero.tex_g0\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_219_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25946_ _06688_ _06640_ _06727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_21069_ _02145_ _02157_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13960_ _07236_ _07243_ _07769_ _07770_ _07771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__22393__A1 _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20240__I _12644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17939__A3 _11079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25877_ _06660_ _06661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13891_ _07701_ _07044_ _07702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_213_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15630_ rbzero.spi_registers.texadd1\[21\] _09291_ _09292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24828_ _05422_ _05423_ _05612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_154_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15561_ _08931_ _09240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24759_ _05490_ _05542_ _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17300_ rbzero.pov.spi_buffer\[29\] _10627_ _10624_ _10631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14512_ _07493_ _08321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_166_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18280_ _11413_ _11415_ _11412_ _11421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15492_ rbzero.spi_registers.buf_texadd0\[10\] _09178_ _09189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13789__I _07599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17231_ rbzero.pov.spi_buffer\[11\] _10579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_127_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26429_ _00339_ clknet_leaf_231_i_clk rbzero.spi_registers.spi_cmd\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14443_ _07543_ _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__26083__B _06842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20459__A1 _09901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17162_ rbzero.pov.spi_counter\[2\] _10524_ _10527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_182_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14374_ rbzero.debug_overlay.playerX\[4\] _08184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_153_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16113_ _09000_ _09646_ _09654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13325_ _07077_ _07139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17093_ _08138_ _10474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__19077__A1 _08153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16044_ _09598_ _09602_ _09603_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13256_ _06996_ _07001_ _07070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_150_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15509__I _09190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13187_ _06991_ _06999_ _07000_ _07001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14413__I _07935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_237_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19803_ rbzero.wall_tracer.stepDistY\[-1\] _12271_ _12575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_202_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17995_ rbzero.wall_tracer.trackDistY\[10\] _11139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_19_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19734_ _12385_ _12387_ _12506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_193_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16946_ _10359_ _10353_ _10360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_208_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22384__A1 _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14861__A2 _08529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19665_ _12405_ _12406_ _12408_ _12222_ _12437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_205_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_220_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16877_ _10272_ _10300_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18616_ _11564_ _11628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15828_ _09438_ _09439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19596_ rbzero.wall_tracer.stepDistX\[-9\] _12202_ _12367_ _12368_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_144_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_248_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_231_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18547_ _11589_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15759_ _09386_ _09388_ _09384_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_220_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20698__A1 _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18478_ rbzero.tex_g1\[53\] rbzero.tex_g1\[52\] _11549_ _11550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17429_ rbzero.pov.spi_buffer\[62\] _10721_ _10718_ _10727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23636__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20440_ _01524_ _01532_ _01533_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_145_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24292__I _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20371_ _01382_ _01394_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__26050__A2 rbzero.wall_tracer.rcp_fsm.o_data\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22110_ rbzero.wall_tracer.rcp_fsm.i_data\[-10\] _03088_ _03102_ _03103_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23090_ _02504_ _02292_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_141_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22041_ rbzero.wall_tracer.stepDistY\[-4\] _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_205_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25800_ _06583_ _06584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_167_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24364__A2 _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26780_ _00690_ clknet_leaf_122_i_clk rbzero.tex_g1\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23992_ rbzero.wall_tracer.rcp_fsm.i_data\[5\] _04770_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22375__A1 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input27_I i_vec_csb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13655__A3 _07463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14852__A2 _08631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25731_ _06470_ _06471_ _06507_ _06515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_22943_ _03670_ _03663_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_223_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15154__I _08933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25662_ _06384_ _06391_ _06446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_67_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22127__A1 _11993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22874_ _02251_ _12961_ _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22127__B2 _11079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14604__A2 _07807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_238_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27401_ _01306_ clknet_leaf_108_i_clk rbzero.wall_tracer.stepDistX\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_238_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24613_ _05098_ _05377_ _05397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_225_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21825_ _08134_ _08140_ _02854_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_25593_ _06297_ _06305_ _06366_ _06330_ _06367_ _06377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__23875__A1 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27332_ _01237_ clknet_leaf_37_i_clk rbzero.wall_hot\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24544_ _05245_ _05328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_164_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21756_ _09927_ _02806_ _02808_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_182_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20707_ _01686_ _01736_ _01797_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27263_ _01168_ clknet_leaf_96_i_clk rbzero.wall_tracer.visualWallDist\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24475_ _05258_ _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_164_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21687_ _11132_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_184_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24416__B _05163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26214_ _00124_ clknet_leaf_13_i_clk rbzero.spi_registers.texadd1\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20638_ _12386_ _01534_ _01729_ _12264_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_23426_ _04271_ _04279_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_150_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27194_ _01099_ clknet_leaf_74_i_clk rbzero.wall_tracer.size\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_34_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23357_ _04098_ _04101_ _04211_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26145_ _00055_ clknet_leaf_215_i_clk rbzero.map_overlay.i_mapdx\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20569_ _09973_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15868__A1 _08928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22308_ _03266_ _03203_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13110_ _06923_ _06924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14090_ rbzero.tex_r1\[36\] _07857_ _07900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26076_ _06802_ _03017_ _06661_ _06843_ _06810_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_23288_ _04073_ _04108_ _04142_ _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13041_ _06857_ _06858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_22239_ _03209_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25027_ _05632_ _05633_ _05811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__14540__A1 _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16293__A1 rbzero.spi_registers.spi_buffer\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16800_ _07708_ _10230_ _10233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_234_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__24355__A2 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17780_ _10943_ _10692_ _10947_ _10950_ _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_206_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14992_ _06894_ _08776_ _08794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26978_ _00888_ clknet_leaf_121_i_clk rbzero.texV\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14843__A2 _07633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16731_ _08182_ _10171_ _10172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25929_ _06710_ _06652_ _06711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13943_ rbzero.map_overlay.i_mapdy\[4\] _07754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_161_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19450_ _12214_ _12162_ _12221_ _12222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_16662_ rbzero.wall_tracer.rayAddendY\[7\] _10107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13874_ rbzero.debug_overlay.playerY\[4\] _07685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_202_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18401_ rbzero.tex_g1\[20\] rbzero.tex_g1\[19\] _11502_ _11506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15613_ _09254_ _09279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19381_ _11456_ net83 _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_232_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23866__A1 _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16593_ rbzero.debug_overlay.vplaneY\[-1\] _08109_ _10042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__18375__I _11480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18332_ _07220_ _11460_ _11463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15544_ rbzero.spi_registers.texadd1\[0\] _09218_ _09227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14359__A1 _07979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18263_ _11405_ _11406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_194_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15475_ rbzero.spi_registers.texadd0\[5\] _09176_ _09177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17214_ _10563_ _10559_ _10566_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_181_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14426_ rbzero.tex_g0\[18\] _07872_ _08235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18194_ _11337_ _11338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_182_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17145_ _09035_ rbzero.pov.ss_buffer\[1\] _10512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_181_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__17848__A2 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14357_ _07203_ _07217_ _08166_ _08167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_52_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13308_ _07119_ _07035_ _07120_ _07121_ _07041_ _07122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_17076_ _10385_ _10462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14288_ rbzero.debug_overlay.vplaneY\[-8\] _08098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15239__I _08987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16027_ _09588_ _09589_ _09587_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13334__A2 _07057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13239_ _07052_ _07053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16779__B _10214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_181_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_174_i_clk_I clknet_5_9__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_146_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17978_ _11110_ _11119_ _11121_ _11122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_224_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19717_ _12275_ _12489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16929_ _09139_ _10345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_224_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20907__A2 _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19773__A2 _12485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19648_ _12417_ _12418_ _12419_ _12267_ _12420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_200_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22109__A1 _12216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16587__A2 _09977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19579_ _12161_ _12350_ _12351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_179_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21610_ gpout1.clk_div\[0\] _11826_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_192_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22590_ rbzero.wall_tracer.wall\[1\] _03476_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_192_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21541_ _12300_ _01803_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17000__A3 _10404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_233_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_99_i_clk_I clknet_5_27__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24260_ _05036_ _05044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21472_ _02521_ _02557_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22535__I _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14762__B _08280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23211_ _04065_ _04066_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_132_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20423_ _01426_ _01427_ _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__17629__I _08809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24191_ _04958_ _04961_ _04962_ _04964_ _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_31_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25846__I _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23142_ _03998_ _03881_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20354_ _12955_ _13033_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24034__A1 _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14522__A1 _08321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23073_ _03668_ _03929_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_178_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20285_ _01378_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_77_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22596__A1 _07241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22024_ _03029_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26901_ _00811_ clknet_leaf_132_i_clk rbzero.tex_r1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_11_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19461__A1 _07701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15078__A2 _07191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16275__A1 _08959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26832_ _00742_ clknet_leaf_199_i_clk rbzero.tex_r0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__22348__A1 _11279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold45 i_gpout0_sel[2] net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_242_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26763_ _00673_ clknet_leaf_221_i_clk gpout0.vpos\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23975_ _04739_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_242_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25714_ _06494_ _06456_ _06497_ _06498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_97_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22926_ _03653_ _03658_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_196_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26694_ _00604_ clknet_leaf_67_i_clk rbzero.pov.ready_buffer\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25645_ _06392_ _06415_ _06429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13841__B _07343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22857_ _02257_ _02403_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_168_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21808_ _02852_ _02855_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25576_ _05949_ _05999_ _06360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_183_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13261__A1 _07053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13590_ _07399_ _07385_ _07400_ _07401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_22788_ _02592_ _02598_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22520__A1 rbzero.wall_tracer.texu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27315_ _01220_ clknet_leaf_94_i_clk rbzero.traced_texa\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__22520__B2 rbzero.row_render.texu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24527_ _05255_ _05311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_148_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21739_ _11103_ _11420_ _11124_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_53_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27246_ _01151_ clknet_leaf_78_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15260_ rbzero.spi_registers.buf_otherx\[0\] _08885_ _09017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24458_ _05002_ _05242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_137_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14211_ _08001_ _08020_ _08021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_23409_ _04189_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27177_ _01082_ clknet_leaf_49_i_clk rbzero.wall_tracer.rayAddendX\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15191_ rbzero.spi_registers.spi_buffer\[11\] _08960_ _08964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16443__I _09900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_229_Right_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24389_ _05144_ _05172_ _05044_ _05173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14142_ rbzero.tex_r1\[57\] _07916_ _07636_ _07952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26128_ _00038_ clknet_leaf_250_i_clk rbzero.spi_registers.spi_buffer\[20\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16502__A2 _09948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26059_ _06828_ _06829_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18950_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _11845_ _11846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14073_ _07848_ _07881_ _07882_ _07883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17901_ rbzero.debug_overlay.facingX\[-6\] _11017_ _11045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18881_ _11786_ _11797_ _11798_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_163_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17274__I _06897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24328__A2 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17832_ _10980_ rbzero.pov.ready_buffer\[69\] _10984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_128_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17763_ _10937_ rbzero.pov.ready_buffer\[44\] _10940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_195_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14975_ _07050_ _08776_ _08777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_221_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19502_ _12273_ _12274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16714_ _10066_ _10150_ _10155_ _10156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_92_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13926_ rbzero.map_overlay.i_mapdx\[0\] _07737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17694_ _10890_ rbzero.pov.ready_buffer\[21\] _10894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16569__A2 _10020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25828__A2 _06605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21562__A2 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19433_ _07708_ _11098_ _12205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16645_ _10077_ _10091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_202_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13857_ _07425_ _07668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_159_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_202_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19364_ rbzero.tex_b1\[57\] rbzero.tex_b1\[56\] _12146_ _12147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16576_ _10025_ _10026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13252__A1 _07065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13788_ _07419_ _07599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18315_ _08870_ _11450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15527_ rbzero.spi_registers.texadd0\[19\] _09206_ _09215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_44_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19295_ _12107_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_215_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18246_ _11389_ _11390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_215_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15458_ rbzero.spi_registers.buf_vshift\[5\] _09165_ _09166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23067__A2 _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14409_ _08215_ _08216_ _08217_ _08218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_41_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18177_ rbzero.map_overlay.i_othery\[0\] _11269_ _11321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15389_ _09113_ _09114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14752__B2 _08558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_22__f_i_clk_I clknet_3_5_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20825__A1 _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17128_ _09928_ _10375_ _10501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14504__A1 _08304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17059_ _08144_ _10448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20070_ _12832_ _12840_ _12842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_204_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16257__A1 _08935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17184__I _10542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25516__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_240_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22050__I0 rbzero.wall_tracer.rcp_fsm.o_data\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23760_ _04599_ _04600_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20972_ _01937_ _01942_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22711_ _03576_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_189_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_194_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23691_ _04536_ _04540_ _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_235_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25430_ _06201_ _06210_ _06213_ _06214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_138_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22642_ _03515_ _03516_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25361_ _06085_ _06086_ _06125_ _05718_ _06145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_22573_ _03466_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18182__B2 _09027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27100_ _01010_ clknet_leaf_139_i_clk rbzero.tex_b1\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_118_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24312_ _05089_ _05093_ _05095_ _05096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_21524_ _02608_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_25292_ _06075_ _05975_ _06022_ _06076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27031_ _00941_ clknet_leaf_134_i_clk rbzero.tex_g0\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24243_ _05026_ _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21455_ _02540_ _12960_ _02427_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_133_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14743__B2 _08522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20406_ _01414_ _01419_ _01499_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24174_ _04826_ _04881_ _04850_ _04879_ _04958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_21386_ _12732_ _02098_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_160_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16496__A1 _08118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20337_ _01430_ _01431_ _12311_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23125_ _03811_ _03812_ _03819_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput35 net35 o_rgb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_246_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_79_Left_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23056_ _03785_ _03798_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20268_ _13037_ _13039_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_179_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13836__B _07646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23230__A2 _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22007_ _03024_ _02986_ _03025_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20199_ _12930_ _12971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14259__B1 _08060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26815_ _00725_ clknet_leaf_180_i_clk rbzero.tex_g1\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_204_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26746_ _00656_ clknet_leaf_229_i_clk rbzero.pov.mosi vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14760_ rbzero.tex_b0\[22\] _08277_ _08567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23958_ _04754_ _04756_ _04752_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_4_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13482__A1 rbzero.texV\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18796__I0 rbzero.tex_r1\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13711_ rbzero.tex_r0\[61\] _07509_ _07522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17043__B _10436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22909_ _03750_ _03752_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_123_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16438__I _09895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14691_ rbzero.tex_b0\[55\] _08496_ _08497_ _08498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26677_ _00587_ clknet_leaf_23_i_clk rbzero.pov.ready_buffer\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23889_ _03010_ _04699_ _04706_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15342__I _09029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16430_ _08839_ _09887_ _09891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_88_Left_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25628_ _05880_ _06328_ _06412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13642_ _07452_ _07453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_122_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13785__A2 _07595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16361_ rbzero.spi_registers.buf_texadd3\[8\] _09840_ _09841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25559_ _06110_ _06118_ _06283_ _06343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_39_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18653__I _11478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13573_ _06882_ _07358_ _07361_ _06858_ _07383_ _07384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_109_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18100_ _11194_ _11208_ _11242_ _11243_ _11244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__18173__B2 rbzero.map_overlay.i_othery\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15312_ rbzero.spi_registers.buf_mapdx\[2\] _09038_ _09057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19080_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] _11924_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_164_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16292_ rbzero.spi_registers.buf_texadd2\[15\] _09780_ _09789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13797__I _07468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18031_ rbzero.wall_tracer.trackDistX\[-3\] _11175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_35_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27229_ _01134_ clknet_leaf_88_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15243_ _09005_ _09001_ _09006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13537__A2 _07347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24797__A2 _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15174_ rbzero.spi_registers.spi_buffer\[7\] _08950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17523__I1 rbzero.tex_b0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19484__I _12255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16487__A1 _09933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14125_ _07495_ _07935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_97_Left_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19982_ _12727_ _12754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14622__S _07928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13746__B _07546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18933_ _11836_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14056_ rbzero.tex_r1\[12\] _07821_ _07865_ _07866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_197_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__23221__A2 _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15517__I _08883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_47_i_clk_I clknet_5_17__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18864_ _11780_ _11783_ _11785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17815_ _10856_ _10973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18795_ _11730_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__19028__I1 rbzero.tex_g0\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20991__B1 _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22032__I0 rbzero.wall_tracer.rcp_fsm.o_data\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19728__A2 _12245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17746_ _10905_ _10928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_221_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14958_ _07050_ _08760_ _08755_ _06892_ _08761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13909_ _07719_ _07720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17677_ _10882_ rbzero.pov.ready_buffer\[15\] _10883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14889_ _08691_ _08692_ _08694_ _08558_ _08595_ _08695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_217_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15214__A2 _08975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19416_ _12168_ _12174_ _12187_ _12188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_16628_ _10053_ _10064_ _10075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_134_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21299__A1 _12222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19659__I _12402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16559_ rbzero.debug_overlay.vplaneY\[0\] _09992_ _10011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19347_ _12137_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_230_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_230_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22085__I _10048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19278_ rbzero.tex_b1\[20\] rbzero.tex_b1\[19\] _12094_ _12098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13528__A2 _07338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18229_ rbzero.map_overlay.i_mapdx\[1\] _11337_ _11373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_143_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21240_ _02243_ _02288_ _02326_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19664__A1 _12425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19394__I _12165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16478__A1 _09933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21171_ _02257_ _02258_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_57_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20122_ _12626_ _12521_ _12894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_74_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15150__A1 _08928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18219__A2 _11360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20053_ _12823_ _12824_ _12825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24930_ _05675_ _05693_ _05652_ _05714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__21774__A2 _12216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24861_ _05330_ _05288_ _05645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24399__S1 _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18738__I _11692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_241_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_26600_ _00510_ clknet_leaf_39_i_clk rbzero.pov.spi_buffer\[69\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23812_ _03287_ _03069_ _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_197_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24712__A2 _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24792_ _05567_ _05575_ _05576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__13464__A1 rbzero.traced_texVinit\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26531_ _00441_ clknet_leaf_39_i_clk rbzero.pov.spi_buffer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23743_ _04535_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_20955_ _02042_ _02027_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15162__I _08917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26462_ _00372_ clknet_leaf_208_i_clk rbzero.debug_overlay.playerX\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_95_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23674_ _12225_ _03472_ _03498_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20886_ rbzero.wall_tracer.size_full\[8\] _01975_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_178_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16953__A2 _10359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25413_ _05605_ _06000_ _06197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14964__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13767__A2 _07577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22625_ _03504_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26393_ _00303_ clknet_leaf_18_i_clk rbzero.spi_registers.buf_texadd2\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25344_ _06124_ _06127_ _06128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22556_ _11292_ _03455_ _03456_ rbzero.traced_texa\[1\] _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_180_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16705__A2 _10145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21507_ _02466_ _02469_ _02467_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_63_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25275_ _06043_ _06058_ _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14506__I _07329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14716__B2 _08522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22487_ _03414_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_248_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_248_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27014_ _00924_ clknet_leaf_187_i_clk rbzero.tex_g0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24226_ _04996_ _05009_ _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21438_ _01953_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_133_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_207_i_clk clknet_5_18__leaf_i_clk clknet_leaf_207_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21462__A1 _12522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24157_ _04818_ _04820_ _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_21369_ _02405_ _02415_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23108_ _02482_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24400__A1 _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24088_ _04865_ _04868_ _04871_ _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_9_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_247_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_229_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15930_ _09514_ _09516_ _09505_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_229_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23039_ _03894_ _03765_ _03895_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__17969__A1 _11112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15861_ rbzero.spi_registers.buf_floor\[1\] _09464_ _09465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17600_ _10831_ _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_0_i_clk i_clk clknet_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_243_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14812_ _07801_ _08614_ _08618_ _07438_ _08198_ _08619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__15444__A2 _09155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18580_ _11607_ _11608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_192_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15792_ _09411_ _09412_ _09406_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__21517__A2 _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17531_ _10792_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14743_ _08546_ _08547_ _08549_ _08522_ _08532_ _08550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_26729_ _00639_ clknet_leaf_32_i_clk rbzero.pov.ready_buffer\[59\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_235_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16168__I _09671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17462_ _06898_ _10751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_158_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13207__A1 rbzero.spi_registers.texadd3\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14674_ _07458_ _07441_ _07473_ _08482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_80_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16413_ rbzero.spi_registers.spi_buffer\[21\] _09876_ _09880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19201_ _12036_ _12044_ _12045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_184_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14955__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13625_ _07434_ _07435_ _07436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22478__B1 _10040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17393_ _10665_ _10700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15800__I _09037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_19132_ _08152_ _11919_ _11976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_41_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16344_ _09827_ _09828_ _09822_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13556_ _07366_ _07367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_212_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19063_ rbzero.tex_g0\[62\] rbzero.tex_g0\[61\] _11908_ _11910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16275_ _08959_ _09771_ _09777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13487_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] _07298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_180_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18014_ rbzero.wall_tracer.trackDistY\[5\] _11155_ _11157_ _11158_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15226_ _08916_ _08992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_124_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19646__A1 rbzero.wall_tracer.visualWallDist\[-5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14860__B _07861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17727__I _10915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15157_ _08935_ _08918_ _08936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14108_ rbzero.tex_r1\[47\] _07916_ _07917_ _07918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_39_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19965_ _12305_ _12306_ _12737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_15088_ _07164_ _08879_ _08880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19949__A2 _12414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18916_ _11825_ _11826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14039_ rbzero.tex_r1\[21\] _07845_ _07849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19896_ _12237_ _12668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input1_I i_debug_map_overlay vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18847_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] _11770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_52_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17462__I _06898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_223_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18778_ rbzero.tex_r1\[54\] rbzero.tex_r1\[53\] _11719_ _11721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_195_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24170__A3 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17729_ _10912_ _10640_ _10916_ _10917_ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_78_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20740_ _01727_ _01830_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__20192__A1 _12236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19389__I _12160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20671_ _01760_ _01762_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14946__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15710__I _09257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22410_ _01661_ _03325_ _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23390_ _11410_ _04243_ _04244_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19885__A1 _10336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22341_ _03292_ _03275_ _03293_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25060_ _05331_ _05641_ _05841_ _05843_ _05844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_22272_ _03209_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14174__A2 _07189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19637__A1 _12405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24630__A1 _05351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24011_ rbzero.wall_tracer.rcp_fsm.i_data\[10\] _08813_ _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21223_ _02178_ _02301_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21154_ _02222_ _02241_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_243_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_243_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20105_ _12633_ _12875_ _12876_ _12877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_10_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2_0_i_clk clknet_0_i_clk clknet_3_2_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_6_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_193_i_clk clknet_5_12__leaf_i_clk clknet_leaf_193_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25962_ _06742_ _06743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21085_ _02045_ _02165_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_208_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20036_ _12433_ _12694_ _12808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24913_ _05310_ _05696_ _05464_ _05418_ _05697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25893_ _06649_ _06642_ _06676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_232_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16623__A1 _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15426__A2 _08885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24844_ _05627_ _05626_ _05628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_213_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_87_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24775_ _05327_ net52 _05436_ _05507_ _05559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_103_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21987_ rbzero.wall_tracer.rcp_fsm.o_data\[1\] rbzero.wall_tracer.size\[9\] _03002_
+ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14010__B _07819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26514_ _00424_ clknet_leaf_32_i_clk rbzero.debug_overlay.vplaneY\[-8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23726_ _04569_ _04570_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_194_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20938_ _01909_ _01911_ _02027_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_56_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26445_ _00355_ clknet_leaf_85_i_clk rbzero.wall_tracer.rayAddendY\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_131_i_clk clknet_5_14__leaf_i_clk clknet_leaf_131_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_23657_ _04505_ _04507_ _04508_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20869_ _01955_ _01958_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13410_ _07194_ _07218_ _07220_ _07221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_126_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22608_ _03493_ _03486_ _03299_ _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14390_ rbzero.color_sky\[2\] _07966_ _08199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26376_ _00286_ clknet_leaf_251_i_clk rbzero.spi_registers.buf_texadd1\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23588_ _04359_ _04361_ _04440_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_148_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25327_ _06110_ _05998_ _06111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13341_ _06883_ _07153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__21683__A1 _08057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22539_ _03446_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_221_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_146_i_clk clknet_5_14__leaf_i_clk clknet_leaf_146_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_118_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16060_ _09611_ _09613_ _09615_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25258_ _06037_ _06041_ _06042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__15362__A1 rbzero.mapdyw\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13272_ _06907_ _07026_ _06919_ _06926_ _07086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_121_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17547__I _10758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15011_ _08809_ _08810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_24209_ _04988_ _04989_ _04990_ _04838_ _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_32_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13912__A2 _07721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25189_ _05972_ _05973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18300__B2 rbzero.vga_sync.vsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16862__A1 _10283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19750_ _12521_ _12522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16962_ _08881_ _10177_ _10373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_18701_ _11671_ _11677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15913_ _09428_ _09504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_120_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19681_ _12425_ _12447_ _12452_ _12453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_200_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16893_ _10281_ _10314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_246_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15844_ _08928_ _09446_ _09452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18632_ _11637_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_235_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_231_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18563_ _11598_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13979__A2 _06884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15775_ rbzero.spi_registers.texadd3\[10\] _09396_ _09400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_232_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23360__A1 _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17514_ rbzero.tex_b0\[18\] rbzero.tex_b0\[17\] _10781_ _10783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14726_ _08525_ _08527_ _08531_ _08522_ _08532_ _08533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_18494_ _11558_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14855__B _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17445_ _10737_ _10735_ _10738_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14657_ _08461_ _08462_ _08464_ _07955_ _07464_ _08465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_138_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23112__A1 _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13608_ _07418_ _07419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17376_ rbzero.pov.spi_buffer\[48\] _10687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_156_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14588_ _08392_ _08393_ _08395_ _08211_ _07589_ _08396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_83_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24860__A1 _05298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23663__A2 _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19115_ rbzero.debug_overlay.facingY\[-4\] _10062_ _11959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16327_ _09814_ _09815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13539_ rbzero.floor_leak\[4\] _07349_ _07329_ rbzero.floor_leak\[3\] _07350_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_131_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19046_ _11900_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_153_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15353__A1 rbzero.mapdxw\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16258_ _09763_ _09764_ _09762_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15209_ _08976_ _08978_ _08971_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13903__A2 _07713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16189_ _09708_ _09710_ _09712_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_239_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21908__S _10125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_225_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19948_ _12703_ _12712_ _12719_ _12720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__21707__I _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19879_ _12632_ _12650_ _12651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__24391__A3 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15705__I _09336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21910_ _02921_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_235_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13419__A1 _07175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22890_ _03638_ _03748_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__24679__A1 _05408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_203_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_203_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21841_ _09989_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_69_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24560_ _05291_ _05294_ _05344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21772_ rbzero.debug_overlay.vplaneX\[-3\] _12184_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23511_ _04302_ _04338_ _04363_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20723_ _01698_ _01707_ _01813_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14919__A1 _07624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24491_ net47 _05275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16536__I _09988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_169_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26230_ _00140_ clknet_leaf_1_i_clk rbzero.spi_registers.texadd1\[21\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23442_ _04294_ _04295_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_190_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20654_ _01649_ _01650_ _01745_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_147_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_i_clk clknet_5_21__leaf_i_clk clknet_leaf_63_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_190_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26161_ _00071_ clknet_leaf_185_i_clk rbzero.floor_leak\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20585_ _01603_ _01624_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_23373_ _04210_ _04212_ _04227_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_33_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25112_ _05393_ _05408_ _05233_ _05301_ _05896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_190_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22324_ _11160_ _03203_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15344__A1 _07757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26092_ rbzero.wall_tracer.rcp_fsm.o_data\[10\] _06846_ _06855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13895__I _07705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25043_ _05760_ _05800_ _05827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_143_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22255_ _11202_ _03204_ _03222_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_78_i_clk clknet_5_28__leaf_i_clk clknet_leaf_78_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13828__C _07638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_221_i_clk_I clknet_5_3__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22090__A1 _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21206_ _02132_ _02159_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22186_ _03104_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_113_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24906__A2 _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21137_ _02224_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13658__A1 rbzero.row_render.texu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26994_ _00904_ clknet_leaf_194_i_clk rbzero.tex_g0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_25945_ _06720_ _06695_ _06725_ _06726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_21068_ _02148_ _02156_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15615__I _09258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20019_ _12790_ _12791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_25876_ _06659_ _06660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_232_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13890_ rbzero.debug_overlay.playerX\[-2\] _07701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output40_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24827_ _05330_ _05492_ _05609_ _05610_ _05611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
Xclkbuf_leaf_16_i_clk clknet_5_4__leaf_i_clk clknet_leaf_16_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_150_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15560_ rbzero.spi_registers.buf_texadd1\[4\] _09232_ _09239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20156__A1 _12660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24758_ _05497_ _05499_ _05541_ _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_69_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14511_ _08316_ _08318_ _08319_ _08320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_23709_ rbzero.wall_tracer.trackDistY\[-8\] _03041_ _04549_ _04556_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15491_ rbzero.spi_registers.texadd0\[10\] _09176_ _09188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24689_ _05472_ _05367_ _05473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_68_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17230_ _10576_ _10572_ _10578_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_194_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26428_ _00338_ clknet_leaf_231_i_clk rbzero.spi_registers.spi_cmd\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14442_ rbzero.tex_g0\[1\] _08250_ _07838_ _08251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19849__A1 _12409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_202_Left_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17161_ rbzero.pov.spi_counter\[2\] _10524_ _10526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20459__A2 _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26359_ _00269_ clknet_leaf_246_i_clk rbzero.spi_registers.buf_texadd1\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14373_ _07708_ _08007_ _08047_ _08182_ _08183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16112_ rbzero.spi_registers.buf_texadd0\[19\] _09644_ _09653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14138__A2 _07920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13324_ _07137_ _07138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_133_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17092_ _10471_ _10397_ _10473_ _09441_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_12_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16043_ _09564_ _09603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22456__I0 _07713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13255_ _07065_ _07013_ _07068_ _07069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_51_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22081__A1 _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13186_ rbzero.spi_registers.texadd0\[17\] _06991_ _07000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19802_ rbzero.wall_tracer.stepDistX\[-1\] _12294_ _12574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_166_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_211_Left_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_166_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17994_ _11137_ _11138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19733_ _12468_ _12485_ _12504_ _12505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__20431__I _12906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16945_ _07681_ _10359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_236_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19664_ _12425_ _12434_ _12435_ _12436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_95_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_220_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16876_ _08042_ _10283_ _10299_ _10300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18615_ _11627_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__26616__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15827_ _09437_ _08852_ _08843_ _09438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_19595_ _12161_ _12366_ _12367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_144_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14074__A1 _07868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18546_ rbzero.tex_r0\[18\] rbzero.tex_r0\[17\] _11587_ _11589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15758_ rbzero.spi_registers.buf_texadd3\[5\] _09387_ _09388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23884__A2 _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14585__B _07580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14709_ _08512_ _08513_ _08515_ _08284_ _08509_ _08516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_18477_ _11543_ _11549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15689_ _09240_ _09336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14077__S _07478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_170_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17428_ rbzero.pov.spi_buffer\[61\] _10726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_16_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17359_ rbzero.pov.spi_buffer\[44\] _10674_ _10671_ _10675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20370_ _01396_ _01444_ _01463_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_160_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14129__A2 _07938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25389__A2 _06093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17187__I _10541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19029_ _11890_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22040_ _03000_ _03045_ _03049_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_207_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22072__A1 _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_17__f_i_clk clknet_3_4_0_i_clk clknet_5_17__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_228_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_215_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_205_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__20341__I _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_95_i_clk_I clknet_5_26__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23991_ _04781_ _04776_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25730_ _06469_ _06512_ _06513_ _06514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_22942_ _02609_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25661_ _06413_ _06443_ _06444_ _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_218_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22873_ _03730_ _03731_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14065__B2 _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27400_ _01305_ clknet_leaf_79_i_clk rbzero.wall_tracer.stepDistX\[-2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__19379__I0 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24612_ _05253_ _05393_ _05394_ _05395_ _05396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_238_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20138__A1 _12907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21824_ _02870_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_25592_ _06327_ _06329_ _06376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13812__A1 _07609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27331_ _01236_ clknet_leaf_37_i_clk rbzero.wall_hot\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24543_ _05275_ _05296_ _05232_ _05300_ _05327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21755_ _10452_ _02697_ _02807_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_149_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20706_ _01687_ _01735_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_164_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27262_ _01167_ clknet_leaf_116_i_clk rbzero.wall_tracer.visualWallDist\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24474_ _05257_ _05258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__24824__A1 _05351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21686_ _11300_ _02729_ _02749_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26213_ _00123_ clknet_leaf_10_i_clk rbzero.spi_registers.texadd1\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23425_ _04272_ _04278_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21638__A1 _09915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27193_ _01098_ clknet_leaf_76_i_clk rbzero.wall_tracer.size\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_20637_ _01715_ _01617_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_150_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26144_ _00054_ clknet_leaf_215_i_clk rbzero.map_overlay.i_othery\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23356_ _04099_ _04100_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_33_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20568_ _01556_ _01660_ _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_150_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22307_ _11168_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26075_ _06842_ _06657_ _06843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23287_ _04029_ _04141_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20499_ _12884_ _12518_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_60_Left_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25026_ _05637_ _05685_ _05748_ _05752_ _05810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_13040_ gpout0.hpos\[8\] _06857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_237_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22238_ _03200_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21810__A1 _10121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22169_ _11983_ _03120_ _03093_ _11067_ _03151_ _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_79_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14991_ _08784_ _08791_ _08792_ _08793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26977_ _00887_ clknet_leaf_122_i_clk rbzero.texV\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13942_ rbzero.map_overlay.i_mapdy\[5\] rbzero.map_overlay.i_mapdy\[3\] _07752_ _07753_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_16730_ _10170_ _10171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25928_ _06649_ _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_191_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_199_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__26078__C _06842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16661_ _09998_ _10105_ _10106_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25859_ _05047_ _06643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13873_ _07213_ _07684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_126_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15612_ _09276_ _09277_ _09278_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18400_ _11505_ _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16592_ _08102_ _08105_ _10041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19380_ _12155_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_158_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15543_ _09225_ _09226_ _09217_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18331_ _10220_ _11462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_167_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_243_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__26094__B _08811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18262_ _11404_ _11405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_166_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15474_ _09150_ _09176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14359__A2 _07202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19487__I _12258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14425_ rbzero.tex_g0\[17\] _08233_ _08220_ _08234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17213_ rbzero.pov.spi_buffer\[7\] _10556_ _10565_ _10566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18193_ _11112_ _11337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_154_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17144_ _10067_ _10393_ _10511_ _10357_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_14356_ _08150_ _08154_ _08158_ _08165_ _08166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_25_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_12__f_i_clk_I clknet_3_3_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13307_ rbzero.spi_registers.texadd3\[3\] _07027_ _07028_ _07121_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14424__I _07484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17075_ rbzero.pov.ready_buffer\[14\] _10460_ _10461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14287_ _08096_ _08078_ _08097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22054__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16026_ _09522_ _09585_ _09589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13238_ _06905_ _07052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_27_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13334__A3 _06905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18340__B _07176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_117_i_clk_I clknet_5_19__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17735__I _10905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_181_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13169_ _06982_ _06983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_225_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_146_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17977_ _11120_ _11101_ _11121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_218_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22357__A2 _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19716_ _12261_ _12487_ _12488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16928_ _07676_ _10328_ _10344_ _10221_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__24568__I _05205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Left_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19647_ _10205_ _10200_ _11096_ _12419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_233_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_205_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16859_ rbzero.pov.ready_buffer\[44\] _10169_ _10284_ _10285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_232_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_200_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19578_ rbzero.wall_tracer.stepDistY\[-8\] _12271_ _12347_ _12349_ _12350_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_179_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14598__A2 _07855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_196_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_196_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18529_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _11576_ _11579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__25059__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21540_ _02016_ _02502_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_233_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21471_ _02523_ _02556_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_160_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Left_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23210_ _03814_ _04058_ _04064_ _01642_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__22293__A1 _11173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20422_ _01426_ _01427_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24190_ _04956_ _04927_ _04974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_44_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23141_ _03769_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_114_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20353_ _12955_ _13033_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24034__A2 _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_211_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23072_ _12733_ _03788_ _03786_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_20284_ _12427_ _12788_ _12958_ _01378_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_12_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22023_ rbzero.wall_tracer.stepDistY\[-9\] _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26900_ _00810_ clknet_leaf_132_i_clk rbzero.tex_r1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_110_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26831_ _00741_ clknet_leaf_199_i_clk rbzero.tex_r0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XPHY_EDGE_ROW_126_Left_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold46 _08765_ net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__23545__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26762_ _00672_ clknet_leaf_221_i_clk gpout0.vpos\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_23974_ _04768_ _04758_ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_230_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25713_ _06453_ _06400_ _06497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_22925_ _03653_ _03658_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_26693_ _00603_ clknet_leaf_65_i_clk rbzero.pov.ready_buffer\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__17775__A2 rbzero.pov.ready_buffer\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25644_ _06392_ _06415_ _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_223_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22856_ _03713_ _03714_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14589__A2 _07845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21807_ _02853_ _02854_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__21859__A1 _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25575_ _06358_ _06359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22787_ _02606_ _03644_ _03645_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_155_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27314_ _01219_ clknet_leaf_110_i_clk rbzero.traced_texa\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24526_ _05259_ _05310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_164_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21738_ _02789_ _02792_ _02793_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__20531__A1 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_135_Left_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_27245_ _01150_ clknet_leaf_78_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24457_ _05240_ _05241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14210__A1 _07101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21669_ _08018_ _02731_ _02728_ _02734_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_191_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14210_ _07101_ _08012_ _08003_ _08020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XPHY_EDGE_ROW_193_Right_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23408_ _04258_ _04261_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_27176_ _01081_ clknet_leaf_49_i_clk rbzero.wall_tracer.rayAddendX\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15190_ _08961_ _08963_ _08954_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24388_ _05135_ _05130_ _05052_ _05172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14141_ rbzero.tex_r1\[56\] _07460_ _07951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26127_ _00037_ clknet_leaf_251_i_clk rbzero.spi_registers.spi_buffer\[19\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23339_ _04171_ _04070_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22036__A1 _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26058_ _04799_ rbzero.wall_tracer.rcp_fsm.o_data\[2\] _08909_ _06829_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14513__A2 _07872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14072_ rbzero.tex_r1\[0\] _07876_ _07882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25009_ _05589_ _05590_ _05587_ _05793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17900_ rbzero.debug_overlay.facingX\[-4\] _11004_ _11044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_238_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18880_ _11795_ _11796_ _11798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_207_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_144_Left_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_219_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17831_ _10979_ _10745_ _10982_ _10983_ _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_128_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17762_ _10915_ _10939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14974_ net9 net8 _08776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_234_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19501_ _12266_ _12267_ _12270_ _12272_ _12273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_156_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16713_ _10152_ _10153_ _10154_ _10155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13925_ rbzero.map_overlay.i_mapdx\[3\] _07736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17693_ _10889_ _10605_ _10892_ _10893_ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_18_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19432_ _10232_ _10233_ _12204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16644_ _10065_ _10089_ _10090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_141_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13856_ _07439_ _07476_ _07666_ _07667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20770__A1 _12660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19363_ _12135_ _12146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16575_ _10024_ _08105_ _10025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13787_ rbzero.tex_r0\[5\] _07597_ _07598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18314_ _11444_ _11449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15526_ _09213_ _09214_ _09202_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_167_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19294_ rbzero.tex_b1\[27\] rbzero.tex_b1\[26\] _12104_ _12107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_43_i_clk_I clknet_5_16__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_215_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18245_ _11388_ _11389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_174_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15457_ _09153_ _09165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_215_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_191_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14408_ rbzero.tex_g0\[26\] _08207_ _08217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_160_Right_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18176_ _11249_ _11320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15388_ _06898_ _09113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_170_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14339_ _08148_ _08149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17127_ _06900_ _10499_ _10500_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_40_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19691__A2 _12419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22027__A1 _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17058_ _06899_ _10447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14504__A2 _08312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13993__I _07329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16009_ _09573_ _09575_ _09576_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19443__A2 _12173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20589__A1 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__25516__A2 _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22050__I1 _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20971_ _01935_ _02058_ _02059_ _01961_ _01986_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_79_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22710_ _03575_ _11225_ _03569_ _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_189_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23690_ _02744_ _04538_ _04539_ _03530_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_164_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_235_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22641_ rbzero.wall_tracer.w\[1\] _03511_ _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25360_ _06143_ _06126_ _06144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_180_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22572_ _11279_ _03461_ _03462_ rbzero.traced_texa\[8\] _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24311_ _05089_ _05094_ _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21523_ _12782_ _02362_ _02607_ _12686_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_75_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25291_ _06020_ _06075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_27030_ _00940_ clknet_leaf_134_i_clk rbzero.tex_g0\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24242_ _05025_ _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_160_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21454_ _02258_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20405_ _01409_ _01413_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_133_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24173_ _04927_ _04956_ _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_21385_ _02465_ _02470_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_32_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16496__A2 _09948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23124_ _03870_ _03871_ _03980_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20336_ rbzero.wall_tracer.size_full\[3\] _13018_ _12912_ _01431_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_222_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput36 net36 o_rgb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_23055_ _03782_ _03910_ _03911_ _03805_ _03831_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_20267_ _12942_ _13038_ _13039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22006_ rbzero.wall_tracer.size_full\[8\] _03020_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_228_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20198_ _12967_ _12969_ _12970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14259__A1 _08057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14259__B2 _08061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26814_ _00724_ clknet_leaf_186_i_clk rbzero.tex_g1\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_99_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19198__A1 _11131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23957_ rbzero.wall_tracer.rcp_fsm.i_data\[-3\] _04755_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26745_ _00655_ clknet_leaf_229_i_clk rbzero.pov.mosi_buffer\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16719__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22741__A2 _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13710_ rbzero.tex_r0\[62\] _07515_ _07520_ _07521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_212_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22908_ _03763_ _03764_ _03765_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_86_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14690_ _07546_ _08497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26676_ _00586_ clknet_leaf_28_i_clk rbzero.pov.ready_buffer\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_123_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23888_ _03599_ _04704_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_196_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13641_ rbzero.row_render.texu\[3\] _07452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25627_ _06403_ _06410_ _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_212_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22839_ _03683_ _03697_ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__14239__I _08048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16360_ _09815_ _09840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25558_ _06339_ _06340_ _06341_ _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_13572_ _07379_ _07381_ _07382_ _07383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_186_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15311_ rbzero.map_overlay.i_mapdx\[2\] _09056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_171_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24509_ _05279_ _05290_ _05293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_87_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16291_ _09787_ _09788_ _09784_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25489_ _05237_ _06020_ _05968_ _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_136_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18030_ rbzero.wall_tracer.trackDistY\[-3\] _11174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15242_ rbzero.spi_registers.spi_buffer\[20\] _09005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_240_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27228_ _01133_ clknet_leaf_81_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26091__C _11825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15173_ _08948_ _08940_ _08949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27159_ _01064_ clknet_leaf_202_i_clk rbzero.wall_tracer.mapY\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14124_ rbzero.tex_r1\[50\] _07932_ _07933_ _07934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16487__A2 _09915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19981_ _12394_ _12454_ _12753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_22_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_152_Left_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14498__A1 _07814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18932_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _11835_ _11836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14055_ rbzero.tex_r1\[13\] _07822_ _07865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_120_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14702__I _07496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18863_ _11780_ _11783_ _11784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__19714__B _12327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17814_ _10848_ _10972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18794_ rbzero.tex_r1\[61\] rbzero.tex_r1\[60\] _11729_ _11730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__20991__A1 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24182__A1 _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__22032__I1 _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17745_ _10903_ _10927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14957_ net5 net4 _08760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14670__A1 _07928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19005__I _11871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15533__I _09208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13908_ gpout0.vpos\[3\] _07719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17676_ _10874_ _10882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_161_Left_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14888_ rbzero.tex_b1\[44\] _07829_ _08693_ _08694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_134_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19415_ _12178_ rbzero.wall_tracer.rayAddendY\[-3\] _12182_ _12186_ _12187_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_176_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16627_ _10065_ _10073_ _10074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13839_ _07639_ _07649_ _07650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__21299__A2 _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19346_ rbzero.tex_b1\[49\] rbzero.tex_b1\[48\] _12136_ _12137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__22496__A1 rbzero.wall_tracer.size\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16558_ rbzero.debug_overlay.vplaneY\[10\] _10008_ _10010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_85_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15509_ _09190_ _09202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_230_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16175__A1 _08955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16364__I _09806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19277_ _12097_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_230_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16489_ _09944_ _09945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__26567__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18228_ rbzero.map_overlay.i_mapdx\[0\] _11347_ _11372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18159_ _11302_ _11303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20274__A3 _13036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21170_ _12522_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15708__I _09349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17195__I _08908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20121_ _12888_ _12892_ _12893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_1_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_228_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_228_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20052_ _12802_ _12803_ _12824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22420__A1 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24860_ _05298_ _05639_ _05643_ _05644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_241_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24173__A1 _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23811_ _04638_ _04619_ _04645_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24791_ _05569_ _05574_ _05575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_240_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13464__A2 rbzero.spi_registers.vshift\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22723__A2 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14487__C _08295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26530_ _00440_ clknet_leaf_38_i_clk rbzero.pov.spi_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23742_ _02761_ _04584_ _03580_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20954_ _02042_ _02027_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26461_ _00371_ clknet_leaf_207_i_clk rbzero.debug_overlay.playerX\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23673_ _11240_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_177_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20885_ _01840_ _01717_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25412_ _06194_ _06195_ _06196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_193_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22624_ rbzero.wall_tracer.texu\[2\] rbzero.texu_hot\[2\] _03503_ _03504_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26392_ _00302_ clknet_leaf_19_i_clk rbzero.spi_registers.buf_texadd2\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13898__I _07708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25343_ _06003_ _05974_ _06126_ _06127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_192_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22555_ _03437_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16166__A1 _08944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21506_ _02589_ _02590_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25274_ _06056_ _06057_ _06058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22486_ rbzero.wall_tracer.size\[1\] _03410_ _03412_ _07367_ _03414_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_20_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_248_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27013_ _00923_ clknet_leaf_191_i_clk rbzero.tex_g0\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24225_ _04862_ _04997_ _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_21437_ _02376_ _02393_ _02522_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14192__A3 _07991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22225__B _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24156_ _04939_ _04893_ _04940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__20265__A3 _13036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21368_ _02408_ _02414_ _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23107_ _03808_ _03830_ _03963_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_82_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20319_ _01409_ _01413_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24087_ _04753_ _04870_ _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_102_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24400__A2 _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21299_ _12222_ _02232_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_9_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23038_ _03763_ _03764_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_228_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15860_ _09463_ _09464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24164__A1 _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16641__A2 _10087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14811_ _07963_ _08615_ _08617_ _08364_ _08618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_153_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15791_ rbzero.spi_registers.buf_texadd3\[14\] _09409_ _09412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24989_ _05561_ _05565_ _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13455__A2 rbzero.spi_registers.vshift\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14652__B2 _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17530_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _10791_ _10792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14742_ rbzero.tex_b0\[35\] _08526_ _08548_ _08549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26728_ _00638_ clknet_leaf_36_i_clk rbzero.pov.ready_buffer\[58\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_216_i_clk_I clknet_5_6__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14673_ _07450_ _07465_ _08481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_17461_ rbzero.pov.spi_buffer\[70\] _10750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_212_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26659_ _00569_ clknet_leaf_158_i_clk rbzero.tex_b0\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_28_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18664__I _11650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19200_ _12037_ _12042_ _12043_ _12044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_16412_ rbzero.spi_registers.buf_texadd3\[21\] _09874_ _09879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13624_ rbzero.row_render.wall\[1\] _07435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14955__A2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17392_ rbzero.pov.spi_buffer\[52\] _10699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__22478__B2 _07433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19131_ _11958_ _11973_ _11974_ _11975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_41_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16343_ _08922_ _09820_ _09828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13555_ rbzero.row_render.size\[1\] _07366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21150__A1 _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25416__A1 _06037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_212_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19062_ _11909_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16274_ rbzero.spi_registers.buf_texadd2\[10\] _09769_ _09776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22914__I _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14707__A2 _07909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13486_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] rbzero.texV\[1\] rbzero.traced_texVinit\[1\]
+ _07297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_180_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18013_ _11156_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.trackDistY\[5\]
+ _11155_ _11157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_164_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15225_ _08989_ _08991_ _08988_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_180_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15156_ rbzero.spi_registers.spi_buffer\[5\] _08935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__20434__I _12912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14107_ _07520_ _07917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19964_ _12728_ _12733_ _12734_ _12735_ _12736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_15087_ _08878_ _08879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14432__I _07532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_240_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_186_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18915_ _07167_ _11825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_14038_ _07343_ _07848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19895_ _12666_ _12667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_129_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16787__C _10221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18846_ _11737_ _11769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_52_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_223_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25498__A4 _06012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18777_ _11720_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15989_ rbzero.spi_registers.buf_mapdx\[4\] _09560_ _09561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__18909__A1 _11779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23902__A1 _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22705__A2 rbzero.wall_tracer.stepDistX\[-5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17728_ _10913_ rbzero.pov.ready_buffer\[32\] _10917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20716__A1 _12433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20716__B2 _12426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17659_ _10865_ _10574_ _10868_ _10870_ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_161_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22096__I _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20670_ _01632_ _01761_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_58_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19329_ rbzero.tex_b1\[42\] rbzero.tex_b1\[41\] _12125_ _12127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16148__A1 _08915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19885__A2 _12006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13511__I _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22340_ _11148_ _03245_ _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22271_ _11193_ _03226_ _03235_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24010_ _04795_ _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_41_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21222_ _02171_ _02305_ _02303_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17139__B _10508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15438__I _08877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21153_ _02223_ _02240_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_243_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_243_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20104_ _12874_ _12649_ _12876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14331__B1 _08036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_165_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25961_ _06901_ _04928_ _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21084_ _02045_ _02165_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_208_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_238_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_208_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20035_ _12697_ _12807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24912_ _05320_ _05296_ _05696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_25892_ _06673_ _06674_ _06675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_226_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24843_ _05325_ _05341_ _05431_ _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__16269__I _09761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24774_ _05536_ _05539_ _05558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_87_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21986_ _03010_ _03011_ _03012_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_87_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23725_ rbzero.wall_tracer.trackDistY\[-6\] _03046_ _04564_ _04570_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26513_ _00423_ clknet_leaf_31_i_clk rbzero.debug_overlay.vplaneY\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_166_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20937_ _01990_ _02026_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__21380__A1 _12465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26444_ _00354_ clknet_5_25__leaf_i_clk rbzero.wall_tracer.rayAddendY\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23656_ _04404_ _04405_ _04452_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_139_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20868_ _01956_ _01437_ _01957_ _12790_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22607_ _07234_ _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26375_ _00285_ clknet_leaf_252_i_clk rbzero.spi_registers.buf_texadd1\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23587_ _04431_ _04439_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__19876__A2 _12647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20799_ _01785_ _01889_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_221_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25326_ _05493_ _06110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_153_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22538_ rbzero.wall_tracer.visualWallDist\[-6\] _03443_ _03444_ rbzero.traced_texa\[-6\]
+ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_153_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17887__A1 _08073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21683__A2 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25257_ _06040_ _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13271_ _06935_ _06977_ _07085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_118_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22469_ _08037_ _03403_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_134_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15010_ _07165_ _08809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_24208_ _04942_ _04967_ _04977_ _04987_ _04991_ _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_60_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18687__I0 rbzero.tex_r1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25188_ _05971_ _05910_ _05972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__17049__B _10436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_248_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24139_ _04825_ _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16311__A1 rbzero.spi_registers.buf_texadd2\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16961_ _10309_ _10372_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18700_ _11676_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22935__A2 _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15912_ _08957_ _09498_ _09503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19680_ _12449_ _12450_ _12451_ _12452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_16892_ _10309_ _10313_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_200_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18631_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _11634_ _11637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15843_ rbzero.spi_registers.buf_sky\[3\] _09438_ _09451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_189_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_243_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18562_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _11597_ _11598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_188_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23514__B _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15774_ _09397_ _09399_ _09395_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17513_ _10782_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14725_ _07935_ _08532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18493_ rbzero.tex_g1\[60\] rbzero.tex_g1\[59\] _11554_ _11558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17444_ rbzero.pov.spi_buffer\[66\] _10732_ _10729_ _10738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14656_ rbzero.tex_g1\[63\] _08448_ _08463_ _08464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14928__A2 _08728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23112__A2 _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13607_ _07339_ _07418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21123__A1 rbzero.wall_tracer.stepDistX\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17375_ _10684_ _10677_ _10686_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_156_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14587_ rbzero.tex_g1\[25\] _08317_ _08394_ _08395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19114_ _08153_ rbzero.wall_tracer.rayAddendY\[5\] _11958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_16326_ _09480_ _09669_ _09814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_13538_ _07348_ _07349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__18343__B _11444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17738__I _10915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19045_ rbzero.tex_g0\[54\] rbzero.tex_g0\[53\] _11898_ _11900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16257_ _08935_ _09759_ _09764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13469_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] _07280_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_140_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_188_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15208_ _08977_ _08969_ _08978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16188_ _09711_ _09712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15139_ _08920_ _08907_ _08921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16302__A1 _08994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_225_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19947_ _12718_ _12719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_226_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17473__I _10758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19878_ _12633_ _12635_ _12649_ _12650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_208_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24128__A1 _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18829_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] _11755_ _11756_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_65_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16089__I _09614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25623__C _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21840_ _02882_ _02885_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_223_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_203_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_203_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19555__A1 _08180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14092__A2 _07901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_1__f_i_clk_I clknet_3_0_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_206_i_clk clknet_5_18__leaf_i_clk clknet_leaf_206_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_21771_ rbzero.debug_overlay.vplaneX\[-3\] _12184_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20165__A2 _12936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25628__A1 _05880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23510_ _04268_ _04362_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20722_ _01692_ _01697_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24490_ _05273_ _05274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_148_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23441_ _04179_ _04059_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20653_ _12661_ _12448_ _01647_ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_18_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_91_i_clk_I clknet_5_26__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_26160_ _00070_ clknet_leaf_223_i_clk rbzero.mapdyw\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23372_ _04216_ _04226_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_144_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22554__I _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20584_ _01674_ _01675_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25111_ _05848_ _05849_ _05895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22323_ _03274_ _03277_ _03279_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26091_ _06846_ _03026_ _06844_ _06854_ _11825_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25042_ _05808_ _05814_ _05815_ _05826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_22254_ _11204_ _03221_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21417__A2 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21205_ _02292_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_22185_ _03108_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_113_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14005__C _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21136_ _02085_ _02103_ _02101_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_246_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_217_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26993_ _00903_ clknet_leaf_194_i_clk rbzero.tex_g0\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_100_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25944_ _06721_ _06724_ _06725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21067_ _02150_ _02155_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13844__C _07541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20018_ _12570_ _12790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_232_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25875_ rbzero.wall_tracer.rcp_fsm.state\[1\] _04928_ _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14607__B2 _07867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24826_ _05606_ _05608_ _05610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_240_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14083__A2 _07635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21969_ rbzero.wall_tracer.size\[3\] _02992_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20156__A2 _12223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24757_ _05501_ _05519_ _05540_ _05541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_201_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15631__I _09258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14510_ rbzero.tex_g0\[52\] _07617_ _08319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23708_ rbzero.wall_tracer.trackDistY\[-8\] _03041_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15490_ _09186_ _09187_ _09175_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24688_ _05356_ _05472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_194_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__25095__A2 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26427_ _00337_ clknet_leaf_249_i_clk rbzero.spi_registers.buf_texadd3\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14441_ _07532_ _08250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14247__I rbzero.debug_overlay.playerY\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23639_ _04476_ _04486_ _04490_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_154_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19849__A2 _12500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17160_ _10522_ _10524_ _10525_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_14372_ _08181_ _08182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_153_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26358_ _00268_ clknet_leaf_245_i_clk rbzero.spi_registers.buf_texadd1\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26044__A1 _06768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14691__B _08497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13323_ _07045_ _07122_ _07126_ _07136_ _07137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_16111_ _09651_ _09652_ _09648_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25309_ _06074_ _06078_ _06092_ _06093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_181_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26289_ _00199_ clknet_leaf_232_i_clk rbzero.spi_registers.buf_floor\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_17091_ rbzero.pov.ready_buffer\[18\] _10472_ _10473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16042_ _09591_ _09601_ _09602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13254_ _07007_ _07012_ _07068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__22456__I1 _07709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13185_ rbzero.spi_registers.texadd3\[17\] _06997_ _06992_ rbzero.spi_registers.texadd2\[17\]
+ _06998_ rbzero.spi_registers.texadd1\[17\] _06999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_248_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_202_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19801_ _12488_ _12571_ _12572_ _12573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__24358__A1 _05133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20712__I _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17993_ _11135_ _07234_ _11136_ _11137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__14846__A1 _08295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22908__A2 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19732_ _12488_ _12493_ _12503_ _12504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_16944_ rbzero.debug_overlay.playerY\[3\] _10358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_198_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19663_ _12335_ _12353_ _12370_ _12435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_205_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19722__B _12360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16875_ _10293_ _10294_ _10298_ _10299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_205_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_220_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18614_ rbzero.tex_r0\[48\] rbzero.tex_r0\[47\] _11623_ _11627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15826_ rbzero.spi_registers.spi_done _09437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19594_ rbzero.wall_tracer.stepDistY\[-9\] _12167_ _12365_ _12366_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_144_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15271__A1 rbzero.map_overlay.i_otherx\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24530__A1 _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18545_ _11588_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13770__B _07580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15757_ _09352_ _09387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_158_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14708_ rbzero.tex_b0\[57\] _08279_ _08514_ _08515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_113_i_clk_I clknet_5_31__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18476_ _11548_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15688_ rbzero.spi_registers.buf_texadd2\[12\] _09328_ _09335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17427_ _10723_ _10724_ _10725_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14639_ rbzero.tex_g1\[46\] _07645_ _08447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_192_i_clk clknet_5_9__leaf_i_clk clknet_leaf_192_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17358_ _10649_ _10674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23892__I0 rbzero.wall_tracer.rcp_fsm.o_data\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16309_ _09800_ _09801_ _09795_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17289_ _10621_ _10619_ _10622_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_153_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19028_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _11887_ _11890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17079__A2 _10443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_130_i_clk clknet_5_15__leaf_i_clk clknet_leaf_130_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_38_i_clk_I clknet_5_7__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_205_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23990_ rbzero.wall_tracer.rcp_fsm.operand\[5\] _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__24364__A4 _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22941_ _03785_ _03798_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_173_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19632__B _10317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25660_ _06399_ _06411_ _06444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22872_ _02624_ _02627_ _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_145_i_clk clknet_5_14__leaf_i_clk clknet_leaf_145_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14776__B _08497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24611_ _05376_ _05390_ _05395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_21823_ _10471_ _08127_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25591_ _06322_ _06369_ _06374_ _06375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_238_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_174_Right_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24542_ _05325_ _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_27330_ _01235_ clknet_leaf_188_i_clk rbzero.row_render.wall\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20069__I _12750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21754_ _10452_ _02697_ _09988_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20705_ _01794_ _01795_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24473_ _05246_ _05250_ _05257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_27261_ _01166_ clknet_leaf_116_i_clk rbzero.wall_tracer.visualWallDist\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21685_ _12046_ _02748_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23424_ _04036_ _04273_ _04277_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26212_ _00122_ clknet_leaf_240_i_clk rbzero.spi_registers.texadd1\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27192_ _01097_ clknet_leaf_77_i_clk rbzero.wall_tracer.size\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_20636_ rbzero.wall_tracer.stepDistX\[5\] _12444_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_202_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21638__A2 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_199_Left_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26143_ _00053_ clknet_leaf_216_i_clk rbzero.map_overlay.i_othery\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23355_ _04095_ _04103_ _04209_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__16282__I _09747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20567_ _01557_ _01659_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_132_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22306_ _03253_ _03263_ _03265_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_143_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26074_ _05008_ _05006_ _06842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_23286_ _04072_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20498_ _12480_ _12379_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13879__A2 rbzero.debug_overlay.playerY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25025_ _05637_ _05638_ _05683_ _05809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_22237_ _11240_ _03204_ _03207_ _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22168_ _11293_ _03104_ _03136_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_21119_ rbzero.wall_tracer.size_full\[10\] _02092_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__19067__I0 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24355__A4 _05111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22099_ _03092_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14990_ _08775_ net9 net8 _07230_ _08792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_26976_ _00886_ clknet_leaf_128_i_clk rbzero.texV\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__23563__A2 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25927_ _06686_ _06646_ _06708_ _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_31_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13941_ _07751_ rbzero.map_overlay.i_mapdy\[1\] rbzero.map_overlay.i_mapdy\[0\] _07752_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_191_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19542__B _12311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16660_ _10089_ _10020_ _10106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_161_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25858_ _06469_ _06512_ _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13872_ _07675_ _07679_ _07680_ _07682_ _07683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__14056__A2 _07821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15611_ _09241_ _09278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_126_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24363__I1 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24809_ _05558_ _05577_ _05592_ _05593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_16591_ _09923_ _10040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_25789_ _06572_ _06569_ _06573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13803__A2 _07579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18330_ _11461_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15542_ rbzero.spi_registers.buf_texadd0\[23\] _09220_ _09226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18261_ _11104_ _11404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15556__A2 _09230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15473_ _09173_ _09174_ _09175_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16753__A1 rbzero.pov.ready_buffer\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17212_ _10564_ _10565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_13_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14424_ _07484_ _08233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_182_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22826__A1 _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18192_ _11301_ _11303_ _11336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__21629__A2 _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17143_ rbzero.pov.ready_buffer\[10\] _10485_ _10511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_14355_ _08159_ _08016_ _08046_ _08160_ _08164_ _08165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_163_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13749__C _07496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13306_ rbzero.spi_registers.texadd2\[3\] _07108_ _07109_ rbzero.spi_registers.texadd1\[3\]
+ _07120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_14286_ _08095_ _08096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17074_ _10395_ _10460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16025_ rbzero.spi_registers.buf_mapdxw\[1\] _09583_ _09588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13237_ _07050_ _07024_ _07051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_110_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13168_ rbzero.spi_registers.texadd2\[13\] _06980_ _06981_ rbzero.spi_registers.texadd0\[13\]
+ _06930_ _06982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__21801__A2 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_181_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13099_ _06912_ _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17976_ _11109_ _11120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_146_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19715_ _12486_ _12487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__24751__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_62_i_clk clknet_5_21__leaf_i_clk clknet_leaf_62_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16927_ rbzero.pov.ready_buffer\[53\] _10288_ _10329_ _10343_ _10344_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__21565__A1 _12211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19646_ rbzero.wall_tracer.visualWallDist\[-5\] _12197_ _12244_ _12418_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16858_ _08049_ _10171_ _10284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_200_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15809_ rbzero.spi_registers.buf_texadd3\[19\] _09420_ _09425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19577_ _12255_ _12348_ _12349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_66_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16992__A1 _10345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16789_ _07699_ _08176_ _10203_ _10223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_172_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_77_i_clk clknet_5_29__leaf_i_clk clknet_leaf_77_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_196_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_196_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18528_ _11578_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18459_ rbzero.tex_g1\[45\] rbzero.tex_g1\[44\] _11538_ _11539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13558__A1 _07039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_233_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21470_ _02536_ _02555_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20421_ _01500_ _01514_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_160_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23140_ _03900_ _03902_ _03996_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_71_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20352_ _01372_ _01446_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_141_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18249__A1 rbzero.wall_tracer.rcp_done vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_i_clk clknet_5_5__leaf_i_clk clknet_leaf_15_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_23071_ _03919_ _03927_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_211_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20283_ _01377_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22022_ _02988_ _03031_ _03036_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26830_ _00740_ clknet_leaf_177_i_clk rbzero.tex_g1\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__19049__I0 rbzero.tex_g0\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_243_Right_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold47 _08773_ net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_26761_ _00671_ clknet_leaf_218_i_clk gpout0.vpos\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_243_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23973_ rbzero.wall_tracer.rcp_fsm.operand\[1\] _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__20359__A2 _10020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25712_ _06491_ _06492_ _06495_ _06496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_22924_ _03666_ _03780_ _03781_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_97_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_230_Left_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_26692_ _00602_ clknet_leaf_65_i_clk rbzero.pov.ready_buffer\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__21183__I _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25643_ _06381_ _06382_ _06427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_22855_ _01957_ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_149_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21806_ _08142_ rbzero.debug_overlay.vplaneX\[-7\] _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25574_ _05980_ _06046_ _06358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22786_ _02591_ _02605_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21911__I rbzero.wall_tracer.rayAddendX\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27313_ _01218_ clknet_leaf_110_i_clk rbzero.traced_texa\[-5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24525_ _05303_ _05308_ _05309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21737_ _11107_ _02782_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27244_ _01149_ clknet_leaf_78_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20527__I _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24456_ _05239_ _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_137_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21668_ _11360_ _02733_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20619_ _01611_ _01612_ _01710_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_23407_ _03772_ _04259_ _04207_ _04260_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_24387_ net70 _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_27175_ _01080_ clknet_5_17__leaf_i_clk rbzero.wall_tracer.rayAddendX\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14525__I _07541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21599_ _02580_ _02683_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14140_ _07945_ _07947_ _07949_ _07923_ _07464_ _07950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_34_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23338_ _04090_ _04105_ _04192_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26126_ _00036_ clknet_leaf_251_i_clk rbzero.spi_registers.spi_buffer\[18\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__26615__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14071_ rbzero.tex_r1\[1\] _07878_ _07881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26057_ _06823_ _06824_ _06827_ _06738_ _06743_ _06828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_23269_ rbzero.wall_tracer.trackDistX\[7\] _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_238_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25008_ _05774_ _05791_ _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_238_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13585__B _07044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17830_ _10980_ rbzero.pov.ready_buffer\[68\] _10983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_219_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_210_Right_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_128_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__26089__C _11825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17761_ _10935_ _10673_ _10930_ _10938_ _00623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_26959_ _00869_ clknet_leaf_114_i_clk rbzero.texV\[-11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14973_ net10 _08775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19500_ rbzero.wall_tracer.stepDistY\[-6\] _12271_ _12244_ _12272_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16712_ _10127_ _10140_ _10154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13924_ _07726_ _07728_ _07731_ _07734_ _07735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_88_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17692_ _10890_ rbzero.pov.ready_buffer\[20\] _10893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_233_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19431_ _12194_ _12196_ _12201_ _12202_ _12203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_18_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16643_ rbzero.wall_tracer.rayAddendY\[6\] _10089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_141_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13855_ _07573_ _07664_ _07665_ _07666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15091__I _08882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20770__A2 _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19362_ _12145_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16574_ _08102_ _10024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_13786_ _07576_ _07597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_202_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18313_ _11431_ _11448_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15525_ rbzero.spi_registers.buf_texadd0\[18\] _09209_ _09214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19293_ _12106_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16726__A1 _08875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18244_ _11387_ _11388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_215_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15456_ rbzero.spi_registers.vshift\[5\] _09163_ _09164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_215_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14407_ rbzero.tex_g0\[27\] _08202_ _08216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18175_ rbzero.map_overlay.i_othery\[2\] _11308_ rbzero.map_rom.i_row\[4\] _07732_
+ _11318_ _11319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_114_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15387_ _09109_ _09110_ _09112_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_154_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20286__A1 _12816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20286__B2 _12750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17126_ rbzero.pov.ready_buffer\[4\] _10379_ _10500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13960__A1 _07236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14338_ rbzero.debug_overlay.facingY\[10\] _08148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__17746__I _10905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17057_ _10427_ _10444_ _10446_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_94_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14269_ rbzero.debug_overlay.facingX\[-2\] _08079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15701__A2 _09340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20038__A1 _12666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19979__A1 _12750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16008_ _09564_ _09576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23775__A2 rbzero.wall_tracer.stepDistY\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14268__A2 _08033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17959_ rbzero.wall_tracer.mapX\[5\] _11103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_224_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20970_ _01943_ _01960_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_174_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15217__A1 _08983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19629_ _12399_ _12220_ _12400_ _12401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_189_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_235_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22640_ _03510_ _03514_ _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18167__B1 _11307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14440__A2 _08248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22571_ _03465_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16825__I _08805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24310_ _04933_ _04849_ _05094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21522_ _02489_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_25290_ _06073_ _06015_ _06074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24241_ _05024_ _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21453_ _02421_ _02537_ _02538_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_133_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15940__A2 _09494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20404_ _01421_ _01440_ _01497_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24172_ _04840_ _04921_ _04900_ _04955_ _04956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_21384_ _02466_ _02469_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_142_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23123_ _03727_ _03979_ _03872_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20335_ rbzero.wall_tracer.size_full\[3\] _13018_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_142_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18890__A1 rbzero.traced_texa\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput37 net37 o_rgb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_23054_ _03799_ _03804_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23766__A2 _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20266_ _12867_ _12940_ _13038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15176__I _08951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21777__A1 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22005_ rbzero.wall_tracer.rcp_fsm.o_data\[8\] _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_228_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14080__I _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20197_ _12968_ _12969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_216_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15456__A1 rbzero.spi_registers.vshift\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26813_ _00723_ clknet_leaf_186_i_clk rbzero.tex_g1\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_216_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19198__A2 _12039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24191__A2 _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26744_ _00654_ clknet_leaf_38_i_clk rbzero.pov.spi_done vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23956_ _04739_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_169_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15208__A1 _08977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22907_ rbzero.wall_tracer.trackDistX\[3\] _01699_ _03630_ _03765_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_168_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26675_ _00585_ clknet_leaf_28_i_clk rbzero.pov.ready_buffer\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23887_ _03008_ _04699_ _04705_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_223_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25626_ _06406_ _06409_ _06410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13640_ _07450_ rbzero.row_render.texu\[1\] _07451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22838_ _03688_ _03696_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14431__A2 _08227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25557_ _06154_ _06118_ _06341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_177_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_7_i_clk_I clknet_5_4__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13571_ _06866_ _07380_ _07361_ _06857_ _07382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_22769_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] _03622_
+ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15310_ _09052_ _09053_ _09055_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24508_ _05252_ net50 _05292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_136_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16290_ rbzero.spi_registers.spi_buffer\[14\] _09782_ _09788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_240_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25488_ _06079_ _06080_ _06081_ _05605_ _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_81_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24246__A3 _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27227_ _01132_ clknet_leaf_89_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15241_ rbzero.spi_registers.spi_buffer\[21\] _08992_ _09004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24439_ _05076_ _04961_ _05015_ _05223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_151_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20268__A1 _13037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15172_ rbzero.spi_registers.spi_buffer\[8\] _08948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_27158_ _01063_ clknet_leaf_199_i_clk rbzero.map_rom.i_row\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_50_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26109_ _00019_ clknet_leaf_232_i_clk rbzero.spi_registers.spi_buffer\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14123_ rbzero.tex_r1\[51\] _07632_ _07933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_19980_ _12725_ _12739_ _12751_ _12752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__16470__I _09926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27089_ _00999_ clknet_leaf_151_i_clk rbzero.tex_b1\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA_clkbuf_leaf_212_i_clk_I clknet_5_7__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18931_ _11829_ _11835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14054_ rbzero.tex_r1\[15\] _07818_ _07642_ _07864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19781__I _12476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15086__I _08877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18862_ _11781_ _11777_ _11782_ _11783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_246_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17813_ _10965_ _10728_ _10968_ _10971_ _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_18793_ _11713_ _11729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_175_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15814__I _09428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24182__A2 _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17744_ _10920_ _10657_ _10923_ _10926_ _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14956_ _08749_ _08753_ _08758_ _08759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_221_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13907_ _07227_ rbzero.map_overlay.i_othery\[2\] _07718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_17675_ _10872_ _10881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_187_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14887_ rbzero.tex_b1\[45\] _07561_ _08693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__16947__A1 _10359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19414_ _12183_ _12185_ _12186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16626_ rbzero.wall_tracer.rayAddendY\[5\] _10073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_217_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13838_ _07640_ _07643_ _07644_ _07647_ _07648_ _07649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_203_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19345_ _12135_ _12136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16557_ rbzero.debug_overlay.vplaneY\[10\] _10008_ _10009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13769_ _07421_ _07580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25958__I _05212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15508_ rbzero.spi_registers.buf_texadd0\[14\] _09194_ _09201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19276_ rbzero.tex_b1\[19\] rbzero.tex_b1\[18\] _12094_ _12097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_230_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16488_ _09896_ _09944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19956__I _12700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18227_ _09056_ _11343_ _11320_ _07736_ _07743_ _11259_ _11371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XANTENNA__14186__A1 _07991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15439_ _09150_ _09151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__25179__B _05943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20259__A1 _12982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18158_ _11252_ _11302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17109_ _10391_ _10487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16380__I _09855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18089_ _11189_ _11232_ _11233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20120_ _12889_ _12890_ _12891_ _12892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__23748__A2 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_228_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19416__A3 _12187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_245_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20051_ _12814_ _12821_ _12822_ _12823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_225_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15724__I _09349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23810_ _04004_ _04644_ _04625_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_225_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_225_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24790_ _05570_ _05571_ _05573_ _05574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__17144__C _10357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23741_ _11174_ _03053_ _04583_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_1_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20953_ _01911_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_178_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16938__A1 _08057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26460_ _00370_ clknet_leaf_207_i_clk rbzero.debug_overlay.playerX\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20884_ _01968_ _01973_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_177_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23672_ _04523_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15610__A1 rbzero.spi_registers.buf_texadd1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25411_ _06015_ _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_191_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22623_ _03474_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_26391_ _00301_ clknet_leaf_20_i_clk rbzero.spi_registers.buf_texadd2\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_193_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_161_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25342_ _06085_ _06086_ _06125_ _05337_ _06126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_22554_ _03435_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21505_ _02471_ _02476_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25273_ _06048_ _06055_ _06057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22485_ _03413_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_133_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27012_ _00922_ clknet_leaf_191_i_clk rbzero.tex_g0\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24224_ _04984_ _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21436_ _02373_ _02394_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_24155_ _04914_ _04928_ _04938_ _04939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_32_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17666__A2 rbzero.pov.ready_buffer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21367_ _02451_ _02452_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_248_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_20318_ _01410_ _01411_ _01412_ _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_23106_ _03810_ _03829_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24086_ _04869_ _04803_ _04795_ _04870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_247_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21298_ _12689_ _01917_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23037_ _03763_ _03764_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_9_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20249_ rbzero.wall_tracer.stepDistY\[2\] _12311_ _13017_ _13020_ _13021_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_219_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_86_i_clk_I clknet_5_25__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14810_ rbzero.row_render.wall\[1\] _08616_ _08617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15790_ rbzero.spi_registers.texadd3\[14\] _09407_ _09411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24988_ _05567_ _05575_ _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_98_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14741_ rbzero.tex_b0\[34\] _08206_ _08548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_54_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26727_ _00637_ clknet_leaf_36_i_clk rbzero.pov.ready_buffer\[57\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23939_ _04738_ _04741_ _04736_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_192_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21922__A1 _10040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19591__A2 _11994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25113__B2 _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17460_ _10748_ _10746_ _10749_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_196_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26658_ _00568_ clknet_leaf_157_i_clk rbzero.tex_b0\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14672_ _08357_ _08430_ _08479_ _08480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16411_ _09875_ _09877_ _09878_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25609_ _06336_ _06345_ _06393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13623_ rbzero.row_render.wall\[0\] _07434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17391_ _10695_ _10688_ _10698_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22478__A2 _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26589_ _00499_ clknet_leaf_36_i_clk rbzero.pov.spi_buffer\[58\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14955__A3 _07225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19130_ _11939_ _11974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16342_ rbzero.spi_registers.buf_texadd3\[3\] _09816_ _09827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23800__B _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13554_ rbzero.row_render.size\[2\] _07365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_137_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_212_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21150__A2 _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_212_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14168__A1 _06888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_171_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19061_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _11908_ _11909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16273_ _09774_ _09775_ _09773_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13485_ rbzero.traced_texVinit\[1\] rbzero.texV\[1\] rbzero.texV\[0\] rbzero.traced_texVinit\[0\]
+ _07296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_18012_ rbzero.wall_tracer.trackDistX\[6\] _11156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_136_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15224_ _08990_ _08984_ _08991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15155_ _08927_ _08930_ _08934_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22650__A2 _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13757__C _07551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20661__A1 _12236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14106_ _07513_ _07916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19963_ _12679_ _12680_ _12735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15086_ _08877_ _08878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__24350__C _05133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14340__A1 _08149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14037_ _07842_ _07844_ _07846_ _07847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_18914_ _11779_ _11824_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_186_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19894_ _12369_ _12666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_247_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14891__A2 _07592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18845_ _11752_ _11768_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24155__A2 _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14588__C _07589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_223_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18776_ rbzero.tex_r1\[53\] rbzero.tex_r1\[52\] _11719_ _11720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15988_ _09547_ _09560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22578__S _09900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14643__A2 _08291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17727_ _10915_ _10916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14939_ _08743_ _08744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17658_ _10866_ rbzero.pov.ready_buffer\[9\] _10870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22377__I _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16609_ _08104_ _08112_ _10057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_148_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16375__I _09815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17589_ _10825_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19328_ _12126_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_100_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19885__A3 _12169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19259_ rbzero.tex_b1\[12\] rbzero.tex_b1\[11\] _12083_ _12087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13906__A1 _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22270_ _11192_ _03221_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24630__A3 _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21221_ _09900_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13382__A2 _07191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21152_ _02225_ _02239_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_218_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19635__B _10208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_243_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20103_ _12874_ _12649_ _12875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13239__I _07052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_108_i_clk_I clknet_5_30__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25960_ _06739_ _06740_ _06741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21083_ _02037_ _02169_ _02170_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_229_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_208_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14882__A2 _08288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20034_ _12799_ _12804_ _12805_ _12806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_208_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24911_ _05320_ _05297_ _05695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13683__B _07493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25891_ _06631_ _06652_ _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25343__A1 _06003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24842_ _05604_ _05621_ _05622_ _05623_ _05625_ _05626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__14634__A2 _07810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24773_ _05519_ _05555_ _05556_ _05557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18765__I _11649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21985_ rbzero.wall_tracer.size\[8\] _03005_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20707__A2 _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26512_ _00422_ clknet_leaf_50_i_clk rbzero.debug_overlay.vplaneX\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_120_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23724_ rbzero.wall_tracer.trackDistY\[-6\] _03046_ _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20936_ _01991_ _02025_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_221_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26443_ _00353_ clknet_leaf_54_i_clk rbzero.wall_tracer.rayAddendY\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20867_ _01604_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23655_ _04394_ _04429_ _04506_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_8__f_i_clk clknet_3_2_0_i_clk clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_22606_ _03491_ _11391_ _03471_ _03482_ _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_36_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26374_ _00284_ clknet_leaf_252_i_clk rbzero.spi_registers.buf_texadd1\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23586_ _04435_ _04438_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20798_ _01788_ _01888_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_221_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_180_Left_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25325_ _06035_ _06014_ _06109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_153_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22537_ _03445_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__17887__A2 rbzero.wall_tracer.rayAddendX\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25256_ _06039_ _06040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_162_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13270_ _06988_ _07083_ _07084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22468_ _08008_ _03403_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_121_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15629__I _09254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24207_ _04950_ _04988_ _04989_ _04990_ _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_21419_ _02504_ _02120_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14533__I _07459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25187_ _05942_ _05944_ _05971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_22399_ _03344_ _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_24138_ _04875_ _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_248_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16960_ _08066_ _10368_ _10371_ _10286_ _10372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_24069_ _04753_ _04802_ _04803_ _04810_ _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_60_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15911_ rbzero.spi_registers.buf_otherx\[2\] _09495_ _09502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_200_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16891_ _08062_ _10301_ _10312_ _10313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_216_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_188_Right_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18630_ _11636_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_204_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15842_ _09140_ _09449_ _09450_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_34_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14625__A2 _07635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18561_ _11586_ _11597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_99_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15773_ rbzero.spi_registers.buf_texadd3\[9\] _09398_ _09399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_31__f_i_clk_I clknet_3_7_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17512_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _10781_ _10782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14724_ rbzero.tex_b0\[42\] _08528_ _08530_ _08531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18492_ _11557_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17443_ rbzero.pov.spi_buffer\[65\] _10737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_131_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14655_ rbzero.tex_g1\[62\] _07804_ _08463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_200_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13606_ _07323_ _07327_ _07417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_185_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17374_ rbzero.pov.spi_buffer\[48\] _10685_ _10682_ _10686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14586_ rbzero.tex_g1\[24\] _07563_ _08394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__21123__A2 _12231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19113_ rbzero.debug_overlay.facingY\[-2\] _11919_ _11957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_171_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16325_ _09812_ _09813_ _09807_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13537_ _07323_ _07347_ _07348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19044_ _11899_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16256_ rbzero.spi_registers.buf_texadd2\[5\] _09757_ _09763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13468_ rbzero.texV\[5\] _07279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16550__A2 rbzero.debug_overlay.vplaneY\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15207_ rbzero.spi_registers.spi_buffer\[13\] _08977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_188_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14443__I _07543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16187_ _09659_ _09711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__18678__I1 rbzero.tex_r1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13399_ _07209_ _07210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15138_ rbzero.spi_registers.spi_buffer\[1\] _08920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_54_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25573__A1 _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24376__A2 _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19946_ _12714_ _12717_ _12718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_225_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15069_ _08857_ _08859_ _08861_ _08862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22387__A1 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14599__B _07646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14864__A2 _07617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19877_ _12638_ _12648_ _12649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_155_Right_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18828_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] _11754_ _11755_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22139__A1 _11991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23705__B _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14616__A2 _07876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23887__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_203_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18759_ rbzero.tex_r1\[46\] rbzero.tex_r1\[45\] _11708_ _11710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_203_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21770_ _08128_ _02813_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_102_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25628__A2 _06328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20721_ _01709_ _01734_ _01811_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__21940__S _10125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20570__B1 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13522__I _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20652_ _01743_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23440_ _04062_ _02292_ _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_147_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22311__A1 _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_i_clk_I clknet_5_22__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23371_ _04218_ _04225_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20583_ _01627_ _01654_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25110_ _05847_ _05850_ _05894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22322_ _11290_ _03264_ _03278_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26090_ _06823_ _06819_ _06854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22253_ _03220_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25041_ _05805_ _05802_ _05803_ _05825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_170_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_3_0_i_clk_I clknet_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24271__B _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21204_ _02291_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22184_ _03163_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_113_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17664__I _10843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21135_ _02113_ _02116_ _02122_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__14304__A1 _07719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26992_ _00902_ clknet_leaf_194_i_clk rbzero.tex_g0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__22378__A1 _12577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14855__A2 _08568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25943_ _06722_ _06723_ _06697_ _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_21066_ _02151_ _02154_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_226_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16057__A1 _09525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20017_ _12706_ _12789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25874_ _05007_ _06657_ _06658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_198_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24825_ _05606_ _05608_ _05609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23878__A1 _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15280__A2 _09032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24756_ _05536_ _05539_ _05540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21968_ rbzero.wall_tracer.rcp_fsm.o_data\[-5\] _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__22550__A1 _11286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23707_ _04528_ _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20919_ _01683_ _01684_ _01879_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_24687_ _05364_ _05470_ _05410_ _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_21899_ _08123_ _11064_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_26426_ _00336_ clknet_leaf_249_i_clk rbzero.spi_registers.buf_texadd3\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14440_ rbzero.tex_g0\[0\] _08248_ _08249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23638_ _04487_ _04488_ _04489_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_230_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14240__B1 _08047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26357_ _00267_ clknet_leaf_246_i_clk rbzero.spi_registers.buf_texadd1\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14791__A1 _07601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14371_ rbzero.debug_overlay.playerX\[-9\] _08181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_153_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23569_ _04412_ _04421_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_64_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16110_ _08997_ _09646_ _09652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25308_ _06083_ _06090_ _06091_ _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_13322_ _07045_ _07131_ _07135_ _07136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_91_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17090_ _10395_ _10472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_133_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26288_ _00198_ clknet_leaf_227_i_clk rbzero.spi_registers.buf_floor\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16532__A2 rbzero.debug_overlay.vplaneY\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13346__A2 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16041_ _09600_ _09601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25239_ _06022_ _06023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14263__I rbzero.debug_overlay.facingX\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13253_ _07002_ _07006_ _07066_ _07067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22480__I _09972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13184_ _06918_ _06998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_36_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19800_ _12276_ _12570_ _12497_ _12502_ _12572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_20_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25555__A1 _06034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_248_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17992_ _11129_ _08374_ _11136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_236_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19731_ _12498_ _12502_ _12503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16943_ _10352_ _10328_ _10356_ _10357_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_224_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25307__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19662_ _12427_ _12428_ _12430_ _12433_ _12434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_205_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16874_ _10295_ _10297_ _10298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_220_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_220_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18613_ _11626_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15825_ _09435_ _09436_ _09430_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19593_ _12167_ _12363_ _12364_ _12365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_220_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23869__A1 _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_220_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18544_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _11587_ _11588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15756_ rbzero.spi_registers.texadd3\[5\] _09385_ _09386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13282__A1 _06906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14707_ rbzero.tex_b0\[56\] _07909_ _08514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_18475_ rbzero.tex_g1\[52\] rbzero.tex_g1\[51\] _11544_ _11548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14438__I _07511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15687_ rbzero.spi_registers.texadd2\[12\] _09326_ _09334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24356__B _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17426_ rbzero.pov.spi_buffer\[61\] _10721_ _10718_ _10725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14638_ _08442_ _08443_ _08445_ _07912_ _07913_ _08446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_7_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14882__B _08497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17749__I _10915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14782__A1 _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13585__A2 _07039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17357_ rbzero.pov.spi_buffer\[43\] _10673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14569_ reg_rgb\[2\] _08377_ _08195_ _08378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__23892__I1 rbzero.wall_tracer.stepDistX\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16308_ _09000_ _09793_ _09801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17288_ rbzero.pov.spi_buffer\[26\] _10615_ _10612_ _10622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19027_ _11889_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16239_ _09744_ _09749_ _09750_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13337__A2 _07147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_224_Right_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18276__A2 _11410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14837__A2 _08529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19929_ _12334_ _12697_ _12699_ _12700_ _12701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_205_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21032__A1 _12689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22940_ _03790_ _03797_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__21583__A2 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22871_ _02625_ _02626_ _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24610_ _05373_ _05375_ _05394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_84_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21822_ _08142_ _08129_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25590_ _06325_ _06368_ _06374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_222_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22532__A1 rbzero.wall_tracer.visualWallDist\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24541_ _05302_ _05324_ _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_5_26__f_i_clk clknet_3_6_0_i_clk clknet_5_26__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_21753_ _10466_ rbzero.wall_tracer.rayAddendX\[-4\] _02805_ _02806_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_47_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27260_ _01165_ clknet_leaf_95_i_clk rbzero.wall_tracer.visualWallDist\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20704_ _01738_ _01767_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24472_ _05241_ _05255_ _05256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22565__I _09939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21684_ _02744_ _12023_ _02745_ _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__24824__A3 _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26211_ _00121_ clknet_leaf_240_i_clk rbzero.spi_registers.texadd1\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23423_ _04273_ _04274_ _04276_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_163_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14773__A1 _08315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27191_ _01096_ clknet_leaf_78_i_clk rbzero.wall_tracer.size\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20635_ _12596_ _12593_ _01726_ _01619_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_19_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__26026__A2 rbzero.wall_tracer.rcp_fsm.o_data\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20846__A1 _12430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26142_ _00052_ clknet_leaf_216_i_clk rbzero.map_overlay.i_othery\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24037__A1 _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23354_ _04097_ _04102_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_150_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20566_ _01558_ _01658_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_34_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22305_ _11293_ _03264_ _03257_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26073_ _06839_ _06840_ _06841_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_20497_ _01588_ _01506_ _01589_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_23285_ _04137_ _04139_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22599__A1 _07241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25024_ _05545_ _05597_ _05808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_14_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22236_ _11213_ _03206_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_219_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16278__A1 rbzero.spi_registers.spi_buffer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22167_ _03140_ _03150_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21118_ _02076_ _02081_ _02077_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22098_ _03089_ _03091_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19067__I1 rbzero.tex_g0\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26975_ _00885_ clknet_leaf_203_i_clk rbzero.texV\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_245_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25926_ _06631_ _06642_ _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21049_ _12661_ _12594_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13940_ rbzero.map_overlay.i_mapdy\[2\] _07751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_31_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_252_i_clk clknet_5_0__leaf_i_clk clknet_leaf_252_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__14967__B net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25857_ _06548_ _06635_ _06641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13871_ gpout0.vpos\[6\] _07681_ _07682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15642__I _09289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19519__A2 _11073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15253__A2 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15610_ rbzero.spi_registers.buf_texadd1\[16\] _09270_ _09277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16450__A1 rbzero.debug_overlay.vplaneY\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24808_ _05587_ _05591_ _05592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_126_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16590_ _10038_ _10039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25788_ _06552_ _06572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_243_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15541_ rbzero.spi_registers.texadd0\[23\] _09218_ _09225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24739_ _05522_ _05523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16202__A1 _08990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_210_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18260_ rbzero.wall_tracer.mapX\[7\] _11403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15472_ _09111_ _09175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_194_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16753__A2 _10183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17211_ _08805_ _10564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_13_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14423_ rbzero.tex_g0\[16\] _08207_ _08232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26409_ _00319_ clknet_leaf_16_i_clk rbzero.spi_registers.buf_texadd3\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14764__A1 rbzero.tex_b0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18191_ _11332_ _11334_ _11335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22826__A2 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27389_ _01294_ clknet_leaf_97_i_clk rbzero.wall_tracer.trackDistY\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17142_ _10509_ _10510_ _10508_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14354_ _08163_ _08164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_123_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16505__A2 _09956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24418__I3 _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13305_ rbzero.spi_registers.texadd0\[3\] _07119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14516__A1 _08295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17073_ _08128_ _10458_ _10459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14285_ _08094_ _08095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16024_ _09584_ _09586_ _09587_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13236_ _07049_ _07050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__19455__A1 _07698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18502__I0 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_205_i_clk clknet_5_18__leaf_i_clk clknet_leaf_205_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13167_ _06927_ _06922_ _06981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_0_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_181_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13098_ _06911_ _06912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17975_ _11111_ _11100_ _11118_ _11119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_146_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22062__I0 rbzero.wall_tracer.rcp_fsm.o_data\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19714_ _12314_ _12317_ _12327_ _12486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_137_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16926_ _10341_ _10342_ _10275_ _10343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14877__B _08497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19645_ _08062_ _12013_ _12255_ _12416_ _12417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_16857_ _10282_ _10283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_232_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16441__A1 _09897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_200_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_200_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15808_ rbzero.spi_registers.texadd3\[19\] _09418_ _09424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19576_ rbzero.wall_tracer.size\[0\] _12246_ _12348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_189_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13255__A1 _07065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16788_ rbzero.debug_overlay.playerX\[-2\] _10222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__22514__A1 rbzero.wall_tracer.texu\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_220_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_196_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15739_ _09349_ _09373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18527_ rbzero.tex_r0\[10\] rbzero.tex_r0\[9\] _11576_ _11578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_207_i_clk_I clknet_5_18__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24086__B _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18458_ _11522_ _11538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17941__A1 _11070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16744__A2 _08181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17409_ _10546_ _10712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_233_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18389_ rbzero.tex_g1\[15\] rbzero.tex_g1\[14\] _11496_ _11499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_99_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20420_ _01508_ _01513_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_209_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20351_ _01374_ _01445_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23070_ _03790_ _03926_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__18249__A2 _11392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20282_ _01376_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_211_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22021_ rbzero.wall_tracer.stepDistY\[-10\] _03034_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_77_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25519__A1 _05889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold37 i_gpout0_sel[3] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__15483__A2 _09030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26760_ _00670_ clknet_leaf_218_i_clk gpout0.vpos\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23972_ _04765_ _04766_ _04767_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold48 i_gpout1_sel[2] net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_input25_I i_tex_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25711_ _06493_ _06494_ _06495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22923_ _03649_ _03665_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_194_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13691__B _07501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26691_ _00601_ clknet_leaf_64_i_clk rbzero.pov.ready_buffer\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_3_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_211_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25642_ _06376_ _06420_ _06425_ _06426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_223_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22854_ _02409_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21805_ _08133_ _08139_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25573_ _05234_ _06033_ _06304_ _06357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__14994__A1 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14078__I _07570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22785_ _02615_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14994__B2 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18185__A1 _11298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27312_ _01217_ clknet_leaf_111_i_clk rbzero.traced_texa\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24524_ _05307_ _05308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22295__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21736_ _08184_ _02773_ _02790_ _02791_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17932__A1 _08085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27243_ _01148_ clknet_leaf_82_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24455_ _05238_ _05239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21667_ _02732_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23406_ _04201_ _04206_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20618_ _01613_ _01621_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27174_ _01079_ clknet_leaf_50_i_clk rbzero.wall_tracer.rayAddendX\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24386_ _05085_ _05119_ _05169_ _05170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_191_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21598_ _02681_ _02682_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16499__A1 _09948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26125_ _00035_ clknet_leaf_252_i_clk rbzero.spi_registers.spi_buffer\[17\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Left_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23337_ _04093_ _04191_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20549_ _01641_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21639__I _09944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26056_ _06684_ _06664_ _06826_ _06670_ _06771_ _06663_ _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_14070_ _07842_ _07877_ _07879_ _07880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_23268_ _03618_ _04122_ _04123_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25007_ _05782_ _05790_ _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_22219_ _03176_ _03192_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23199_ _03726_ _04054_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_238_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22992__A1 _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_156_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16671__A1 _08096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_191_i_clk clknet_5_9__leaf_i_clk clknet_leaf_191_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_128_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14972_ _08744_ _08773_ _08774_ net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_17760_ _10937_ rbzero.pov.ready_buffer\[43\] _10938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26958_ _00868_ clknet_leaf_182_i_clk rbzero.tex_r1\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__21547__A2 _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16711_ _10143_ _10153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13923_ _07214_ _07732_ _07722_ _07102_ _07733_ _07734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_25909_ _05028_ _06685_ _06690_ _06691_ _06692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__16468__I _09896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17691_ _10884_ _10892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26889_ _00799_ clknet_leaf_176_i_clk rbzero.tex_r0\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_89_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15372__I _09074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19430_ _12162_ _12202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_16642_ _10072_ _10078_ _10085_ _10049_ _10088_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13854_ net18 _07665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13237__A1 _07050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24497__A1 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16573_ _08117_ _08107_ _10023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14985__A1 _07178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19361_ rbzero.tex_b1\[56\] rbzero.tex_b1\[55\] _12141_ _12145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_178_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13785_ rbzero.tex_r0\[6\] _07595_ _07462_ _07596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18312_ _11433_ _11446_ _11448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15524_ rbzero.spi_registers.texadd0\[18\] _09206_ _09213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19292_ rbzero.tex_b1\[26\] rbzero.tex_b1\[25\] _12104_ _12106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18243_ _11386_ _11387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_155_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15455_ _09150_ _09163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_215_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_215_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14406_ _08214_ _08215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18174_ rbzero.map_overlay.i_otherx\[0\] rbzero.map_rom.f4 _11318_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_167_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15386_ _09111_ _09112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17125_ _09902_ _10375_ _10499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14337_ _07205_ _08120_ _08146_ _08147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__21483__A1 _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_144_i_clk clknet_5_14__leaf_i_clk clknet_leaf_144_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17056_ rbzero.pov.ready_buffer\[32\] _10445_ _10446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_94_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14268_ _08003_ _08033_ _08077_ _08078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_40_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16007_ _08946_ _09574_ _09575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19979__A2 _12676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13219_ _06906_ _07024_ _07032_ _07033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_59_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14199_ _07975_ _08003_ _08008_ _08009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_148_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18858__I _11737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_159_i_clk clknet_5_10__leaf_i_clk clknet_leaf_159_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__17762__I _10915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13476__A1 rbzero.texV\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17958_ rbzero.wall_tracer.mapX\[6\] _11101_ _11102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_100_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16909_ _10327_ _10328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17889_ rbzero.wall_tracer.rayAddendX\[9\] _11033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15282__I _09034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19628_ rbzero.wall_tracer.stepDistX\[-10\] _11386_ _12400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_215_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19559_ rbzero.wall_tracer.size\[1\] _12247_ _12330_ _12166_ _12331_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_76_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18167__A1 _07757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18167__B2 rbzero.map_overlay.i_mapdy\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22570_ _11281_ _03461_ _03462_ rbzero.traced_texa\[7\] _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_158_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21710__A2 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21521_ _02591_ _02605_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_145_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13530__I _07340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24240_ _05023_ _05011_ _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__19667__A1 _07705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21452_ _02423_ _02428_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25359__C _06003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20403_ _01406_ _01420_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21383_ _02467_ _02468_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_24171_ _04922_ _04886_ _04825_ _04954_ _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_189_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13951__A2 _07757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17142__A2 _10510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23122_ _03868_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20334_ _12183_ _12005_ _12181_ _01428_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_248_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__23215__A2 _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23053_ _03799_ _03804_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_20265_ _12952_ _13034_ _13036_ _13037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xoutput38 net38 o_rgb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__14361__I rbzero.debug_overlay.playerX\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22004_ _03022_ _03011_ _03023_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20196_ _12553_ _12968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_228_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26812_ _00722_ clknet_leaf_186_i_clk rbzero.tex_g1\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_208_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13467__A1 rbzero.traced_texVinit\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22726__A1 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26743_ _00653_ clknet_leaf_42_i_clk rbzero.pov.ready_buffer\[73\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23955_ _04753_ _04743_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20201__A2 _12700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22906_ rbzero.wall_tracer.stepDistX\[4\] _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_224_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13219__A1 _06906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26674_ _00584_ clknet_leaf_28_i_clk rbzero.pov.ready_buffer\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_23886_ _01993_ _04704_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24479__A1 _05261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_123_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25625_ _06407_ _06339_ _06408_ _06409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_195_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22837_ _03690_ _03695_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14967__A1 _07175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23151__A1 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25556_ _05972_ _06110_ _06340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_52_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13570_ _07378_ _06863_ _06866_ _07380_ _07381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_22768_ _11163_ _01699_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_177_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20538__I _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21701__A2 _12051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24507_ _05279_ _05290_ _05291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_137_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21719_ _02768_ _02776_ _02777_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25487_ _06073_ _05968_ _06271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_109_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22699_ _11220_ _12243_ _03565_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_93_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_82_i_clk_I clknet_5_28__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_27226_ _01131_ clknet_leaf_81_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_156_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15240_ _08999_ _09002_ _09003_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24438_ _04932_ _05089_ _05222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_192_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_61_i_clk clknet_5_21__leaf_i_clk clknet_leaf_61_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15171_ _08945_ _08947_ _08934_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_27157_ _01062_ clknet_leaf_201_i_clk rbzero.map_rom.a6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24369_ _04806_ _04946_ _05046_ _05153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14122_ _07515_ _07932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26108_ _00018_ clknet_leaf_232_i_clk rbzero.spi_registers.spi_buffer\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27088_ _00998_ clknet_leaf_151_i_clk rbzero.tex_b1\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_104_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15695__A2 _09340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26039_ _06626_ _06733_ _06624_ _06621_ _06632_ _06667_ _06812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_18930_ _11834_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14053_ rbzero.tex_r1\[14\] _07805_ _07863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_76_i_clk clknet_5_30__leaf_i_clk clknet_leaf_76_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_162_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22965__A1 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21768__A2 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18861_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] _11782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_207_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15447__A2 _09157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Left_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__20440__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17812_ _10966_ rbzero.pov.ready_buffer\[62\] _10971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18792_ _11728_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__24182__A3 _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14955_ net5 net4 _07225_ _08757_ _08758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_17743_ _10921_ rbzero.pov.ready_buffer\[38\] _10926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_222_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23390__A1 _11410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13906_ _07697_ _07716_ _07257_ _07717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_14886_ rbzero.tex_b1\[47\] _07577_ _08603_ _08692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17674_ _10873_ _10587_ _10877_ _10880_ _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_19413_ _12184_ _12185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__25131__A2 _05889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14958__A1 _07050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13837_ _07526_ _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16625_ _10071_ _10072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_217_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14958__B2 _06892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_i_clk clknet_5_5__leaf_i_clk clknet_leaf_14_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_193_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15830__I _09113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16556_ _10007_ _10008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18346__C _11473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19344_ _12071_ _12135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19897__A1 _12667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13768_ _07420_ _07579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_75_Left_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15507_ rbzero.spi_registers.texadd0\[14\] _09192_ _09200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16487_ _09933_ _09915_ _09942_ _09943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14446__I _07601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19275_ _12096_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_210_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13699_ rbzero.tex_r0\[59\] _07509_ _07510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_230_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15438_ _08877_ _09150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18226_ _11107_ _11369_ _11370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14186__A2 _07995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15383__A1 rbzero.floor_leak\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_29_i_clk clknet_5_22__leaf_i_clk clknet_leaf_29_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_127_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_209_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15369_ rbzero.spi_registers.buf_leak\[1\] _09092_ _09099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18157_ _11269_ _11301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_170_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17108_ _10484_ _10393_ _10486_ _10357_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_18088_ _11224_ _11227_ _11231_ _11232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15277__I _09029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17039_ _08153_ _10432_ _10433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16883__A1 _10295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_228_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_84_Left_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_245_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20050_ _12794_ _12795_ _12822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_245_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20911__I _12300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22708__A1 _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13525__I _07335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23740_ _04581_ _04582_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20952_ _01904_ _01908_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_240_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21931__A2 _10087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25122__A2 _05905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14949__A1 _08750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23671_ _04522_ _11140_ _02767_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20883_ _12694_ _01969_ _01972_ _12693_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25410_ _05718_ _06194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_93_Left_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22622_ _03502_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26390_ _00300_ clknet_leaf_20_i_clk rbzero.spi_registers.buf_texadd2\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_220_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_104_i_clk_I clknet_5_30__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25341_ _05946_ _05961_ _05964_ _06125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__20498__A2 _12379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21695__A1 _12036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22553_ _03454_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__21898__B _10113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13260__I _07044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21504_ _02465_ _02470_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25272_ _06048_ _06055_ _06056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_63_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22484_ rbzero.wall_tracer.size\[0\] _03410_ _03412_ _07370_ _03413_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27011_ _00921_ clknet_leaf_189_i_clk rbzero.tex_g0\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24223_ _05006_ _05007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21435_ _02416_ _02431_ _02520_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_20_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16571__I _09944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21189__I _12383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25884__I _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24154_ _04923_ _04929_ _04937_ _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_161_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21366_ _02400_ _02433_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_169_Right_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23105_ _03959_ _03960_ _03961_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16874__A1 _10295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20317_ _12421_ _12380_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14091__I _07459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_248_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24085_ _04802_ _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21297_ _02234_ _02383_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_9_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23036_ rbzero.wall_tracer.stepDistX\[5\] _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_9_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20248_ _13018_ _13019_ _12277_ _13020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_229_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20422__A2 _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_29_i_clk_I clknet_5_22__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20179_ _12950_ _12728_ _12936_ _12951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__14101__A2 _07909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24164__A3 _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24987_ _05567_ _05575_ _05771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_231_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14740_ rbzero.tex_b0\[32\] _08541_ _07861_ _08547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23938_ rbzero.wall_tracer.rcp_fsm.i_data\[-7\] _04740_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26726_ _00636_ clknet_leaf_36_i_clk rbzero.pov.ready_buffer\[56\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_21__f_i_clk_I clknet_3_5_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_212_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25113__A2 _05333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26657_ _00567_ clknet_leaf_157_i_clk rbzero.tex_b0\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14671_ _07888_ _08454_ _08478_ _07477_ _08479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_86_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_23869_ _03539_ _04694_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_158_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16410_ _09855_ _09878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25608_ _06384_ _06391_ _06392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_157_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13622_ _07432_ _07433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_196_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17390_ rbzero.pov.spi_buffer\[52\] _10697_ _10693_ _10698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26588_ _00498_ clknet_leaf_35_i_clk rbzero.pov.spi_buffer\[57\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__23675__A2 _12043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16341_ _09825_ _09826_ _09822_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25539_ _06269_ _06169_ _06306_ _06323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21686__A1 _11300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13553_ rbzero.row_render.size\[3\] _07364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_212_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19060_ _11892_ _11908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_212_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16272_ _08955_ _09771_ _09775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22483__I _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13484_ _07293_ _07294_ _07295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_42_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27209_ _01114_ clknet_leaf_76_i_clk rbzero.wall_tracer.stepDistY\[-6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_18011_ rbzero.wall_tracer.trackDistX\[5\] _11155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_164_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15223_ rbzero.spi_registers.spi_buffer\[16\] _08990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_136_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__18303__A1 _07139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15154_ _08933_ _08934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_91_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14105_ rbzero.tex_r1\[46\] _07645_ _07915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16865__A1 rbzero.pov.ready_buffer\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20661__A2 _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19962_ _12679_ _12680_ _12734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_205_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15085_ _08876_ _08877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14036_ rbzero.tex_r1\[23\] _07845_ _07846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18913_ rbzero.traced_texa\[10\] rbzero.texV\[10\] _11823_ _11824_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__14340__A2 _08078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24203__I _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19893_ _12663_ _12664_ _12665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_18844_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] _11767_ _11768_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_59_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18775_ _11713_ _11719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_223_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15987_ _09558_ _09559_ _09553_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13345__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13300__B1 _07109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17726_ _09034_ _10915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14938_ net21 _08743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__19460__C _12231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13851__A1 _07555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17657_ _10865_ _10570_ _10868_ _10869_ _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14869_ _08316_ _08673_ _08674_ _08675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_188_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25969__I _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16608_ _08116_ _08110_ _10056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20178__I _12949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17588_ rbzero.tex_b0\[50\] rbzero.tex_b0\[49\] _10823_ _10825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19327_ rbzero.tex_b1\[41\] rbzero.tex_b1\[40\] _12125_ _12126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16539_ _09991_ _09992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_161_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19258_ _12086_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18209_ _11337_ _11303_ _11352_ _11353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16391__I _09814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13906__A2 _07716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19189_ _12031_ _12032_ _12033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__19342__I0 rbzero.tex_b1\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15001__S _07185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_247_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21220_ _02307_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21151_ _02230_ _02238_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20102_ _12635_ _12874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_229_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14331__A2 _08006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21082_ _02040_ _02166_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_229_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20033_ _12746_ _12748_ _12805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_208_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24910_ _05640_ _05530_ _05580_ _05298_ _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_clkbuf_leaf_30_i_clk_I clknet_5_22__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14779__C _08565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25890_ _06630_ _06647_ _06673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_176_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23952__I _10491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24841_ _05604_ _05624_ _05625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_225_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24772_ _05501_ _05540_ _05556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21984_ _02983_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_87_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26511_ _00421_ clknet_leaf_60_i_clk rbzero.debug_overlay.vplaneX\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23723_ _02750_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20935_ _01992_ _02024_ _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_194_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25879__I _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26442_ _00352_ clknet_leaf_54_i_clk rbzero.wall_tracer.rayAddendY\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23654_ _04367_ _04393_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_25_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20866_ _12498_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_166_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_238_Right_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22605_ _02732_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__21668__A1 _11360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26373_ _00283_ clknet_leaf_252_i_clk rbzero.spi_registers.buf_texadd1\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23585_ _04436_ _04316_ _04437_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20797_ _01793_ _01887_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25324_ _06066_ _06106_ _06107_ _06108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_148_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22536_ rbzero.wall_tracer.visualWallDist\[-7\] _03443_ _03444_ rbzero.traced_texa\[-7\]
+ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25255_ _06038_ _05811_ _06032_ _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_107_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22467_ _08012_ _03403_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24206_ _04975_ _04990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_21418_ _02016_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25186_ _05969_ _05970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_22398_ _03342_ _11405_ _03343_ _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24137_ _04884_ _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_103_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21349_ _02327_ _02435_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_124_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_248_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24068_ _04806_ _04827_ _04840_ _04851_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23593__A1 _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15645__I _09302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23019_ _03841_ _03876_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15910_ _09500_ _09501_ _09491_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_235_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16890_ _10288_ _10310_ _10311_ _10282_ _10312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_246_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15841_ _08924_ _09446_ _09450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20159__A1 _12398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18560_ _11596_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15772_ _09117_ _09398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__17024__A1 rbzero.pov.ready_buffer\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17511_ _10780_ _10781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14723_ rbzero.tex_b0\[43\] _08529_ _08530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_86_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26709_ _00619_ clknet_leaf_61_i_clk rbzero.pov.ready_buffer\[39\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_18491_ rbzero.tex_g1\[59\] rbzero.tex_g1\[58\] _11554_ _11557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16476__I _08099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14654_ rbzero.tex_g1\[60\] _07940_ _07907_ _08462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17442_ _10734_ _10735_ _10736_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_157_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13605_ _07354_ _07389_ rbzero.row_render.size\[10\] _07353_ _07416_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_205_Right_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_200_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14585_ rbzero.tex_g1\[26\] _07872_ _07580_ _08393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__18691__I _11649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17373_ _10649_ _10685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19112_ _08151_ _10107_ _11956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__22427__B _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16324_ _09667_ _09804_ _09813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13536_ _07272_ _07276_ _07310_ _07347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__20331__A1 _12283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16255_ _09758_ _09760_ _09762_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19043_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _11898_ _11899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14936__I1 _08741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13467_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] _07278_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15206_ rbzero.spi_registers.spi_buffer\[14\] _08975_ _08976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_211_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_188_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16186_ _08973_ _09709_ _09710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_188_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13398_ gpout0.hpos\[5\] gpout0.hpos\[4\] _07208_ gpout0.hpos\[6\] _07209_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__23820__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15137_ _08915_ _08918_ _08919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_199_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19945_ _12715_ _12716_ _12717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_15068_ rbzero.spi_registers.spi_counter\[2\] _08859_ _08860_ _08861_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_239_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_225_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14019_ _07804_ _07829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19876_ _12523_ _12647_ _12648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18827_ _11753_ _11754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__18866__I _08753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18758_ _11709_ _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_203_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17015__A1 rbzero.pov.ready_buffer\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_203_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17709_ _10847_ _10903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18689_ rbzero.tex_r1\[16\] rbzero.tex_r1\[15\] _11666_ _11670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_102_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20720_ _01690_ _01708_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_172_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20570__B2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20651_ _12590_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23370_ _04221_ _04224_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20582_ _01572_ _01626_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22321_ _09926_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18106__I rbzero.map_rom.i_row\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25261__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__22075__A1 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25040_ _05807_ _05816_ _05823_ _05824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_22252_ _11248_ _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24271__C _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21203_ _11296_ _12229_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22183_ _11094_ _03092_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21134_ _02185_ _02221_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_113_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26991_ _00901_ clknet_leaf_131_i_clk rbzero.tex_g0\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA_clkbuf_3_7_0_i_clk_I clknet_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22378__A2 _08041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25942_ _05995_ _06614_ _06723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_21065_ _02152_ _02153_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__23682__I _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20016_ _12787_ _12788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_25873_ _05022_ _05028_ _06633_ _06656_ _06657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_214_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_213_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17680__I _10884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23327__A1 _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24824_ _05351_ _05607_ _05354_ _05608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_216_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17006__A1 rbzero.pov.ready_buffer\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24755_ _05460_ _05537_ _05538_ _05539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__21889__A1 _10113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21967_ _02997_ _02998_ _02999_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23706_ _11203_ _04529_ _04553_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20918_ _01873_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_194_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24686_ _05374_ _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_167_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21898_ _02936_ _02938_ _10113_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_193_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26425_ _00335_ clknet_leaf_249_i_clk rbzero.spi_registers.buf_texadd3\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23637_ _04397_ _04391_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20849_ _12413_ _01607_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13043__A2 _06859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14240__A1 _08042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19400__I _12171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14240__B2 _08049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26356_ _00266_ clknet_leaf_248_i_clk rbzero.spi_registers.buf_texadd1\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14370_ rbzero.debug_overlay.playerX\[-8\] _08180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__20313__A1 _12885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23568_ _04415_ _04420_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_30_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25307_ _06024_ _06007_ _06091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13321_ rbzero.spi_registers.texadd0\[1\] _07127_ _07134_ _06905_ _07135_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_181_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22519_ _03433_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_26287_ _00197_ clknet_leaf_228_i_clk rbzero.spi_registers.buf_floor\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23499_ _04245_ _04246_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16040_ _09599_ _09600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25238_ _06009_ _06007_ _06022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13252_ _07065_ _07007_ _07066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25169_ _05896_ _05952_ _05953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13183_ _06922_ _06997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_36_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24358__A3 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17991_ _07774_ _11135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_236_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_183_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19730_ _12501_ _12502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16942_ _10220_ _10357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_198_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19661_ _12432_ _12433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_245_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_205_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16873_ rbzero.debug_overlay.playerY\[-7\] _10296_ _10297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__14059__B2 _07867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18612_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _11623_ _11626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_220_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15824_ rbzero.spi_registers.buf_texadd3\[23\] _09118_ _09436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19592_ rbzero.wall_tracer.size_full\[-9\] _12172_ _12364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18543_ _11586_ _11587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14719__I _07537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15755_ _09349_ _09385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14706_ rbzero.tex_b0\[58\] _08506_ _08280_ _08513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18474_ _11547_ _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15686_ _09332_ _09333_ _09325_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23033__S _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17425_ _10712_ _10724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14637_ rbzero.tex_g1\[42\] _07909_ _08444_ _08445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_16_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14568_ _07770_ _08376_ _07231_ _08377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_17356_ _10670_ _10666_ _10672_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16307_ rbzero.spi_registers.buf_texadd2\[19\] _09791_ _09800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13519_ _07295_ _07303_ _07304_ _07330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_17287_ rbzero.pov.spi_buffer\[25\] _10621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14499_ _07493_ _08308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22057__A1 _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19026_ rbzero.tex_g0\[46\] rbzero.tex_g0\[45\] _11887_ _11889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16238_ _09711_ _09750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16169_ rbzero.spi_registers.buf_texadd1\[8\] _09696_ _09697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24429__S0 _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_203_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20191__I _12334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25546__A2 _06329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14298__A1 _08106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14403__B _08211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15285__I _09028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14298__B2 _08107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19928_ _12352_ _12700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_205_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21032__A2 _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19859_ _12625_ _12627_ _12630_ _12631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_214_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22870_ _02668_ _02669_ _03728_ _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__25931__B _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21821_ _02811_ _02867_ _02868_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_84_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24540_ _05309_ _05318_ _05323_ _05324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_21752_ _02803_ _02804_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20703_ _01679_ _01737_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24471_ _05254_ _05255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16844__I _07167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21683_ _08057_ _02746_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26210_ _00120_ clknet_leaf_240_i_clk rbzero.spi_registers.texadd1\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23422_ _04036_ _04275_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27190_ _01095_ clknet_leaf_77_i_clk rbzero.wall_tracer.size\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_20634_ rbzero.wall_tracer.stepDistX\[4\] _12444_ _01725_ _01726_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__22296__A1 _11287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_150_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26141_ _00051_ clknet_leaf_216_i_clk rbzero.map_overlay.i_othery\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20846__A2 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23353_ _04198_ _04207_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20565_ _01561_ _01657_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_144_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23677__I _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22304_ _03209_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26072_ _04799_ rbzero.wall_tracer.rcp_fsm.o_data\[4\] _09113_ _06841_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_23284_ _03772_ _04080_ _04089_ _04138_ _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_33_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13328__A3 _06879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20496_ _01504_ _01505_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__23796__A1 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25023_ _05598_ _05757_ _05806_ _05807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__22599__A2 _08752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17675__I _10872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22235_ _03205_ _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22166_ rbzero.wall_tracer.rcp_fsm.i_data\[-1\] _03144_ _03149_ _03150_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__26697__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__19890__I _12661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21117_ _02089_ _02099_ _02204_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_22097_ _03090_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_26974_ _00884_ clknet_leaf_123_i_clk rbzero.texV\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_227_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25925_ _05076_ _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21048_ _02000_ _12383_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17624__B _10256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13870_ rbzero.debug_overlay.playerY\[3\] _07681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_25856_ _06639_ _06640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_161_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24807_ _05589_ _05590_ _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14997__C1 _07178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25787_ _06549_ _06570_ _06571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_22999_ _03732_ _03739_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14461__A1 _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23720__A1 _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15540_ _07025_ _09180_ _09224_ _09182_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_24738_ _05520_ _05521_ _05467_ _05522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_97_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15471_ rbzero.spi_registers.buf_texadd0\[4\] _09165_ _09174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27457_ _01362_ clknet_leaf_71_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24669_ _05392_ _05405_ _05453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_166_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_152_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14422_ _08225_ _08228_ _08230_ _08215_ _07465_ _08231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_17210_ rbzero.pov.spi_buffer\[6\] _10563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_194_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26408_ _00318_ clknet_leaf_13_i_clk rbzero.spi_registers.buf_texadd3\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14764__A2 _08518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15961__A1 _09525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18190_ _11333_ _11334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_27388_ _01293_ clknet_leaf_99_i_clk rbzero.wall_tracer.trackDistY\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__19152__A1 _11990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14353_ _08161_ _08064_ _08060_ _08162_ _08163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_17141_ rbzero.pov.ready_buffer\[9\] _10472_ _10510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_182_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26339_ _00249_ clknet_leaf_238_i_clk rbzero.spi_registers.buf_texadd0\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13304_ _07062_ _07117_ _07118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__22039__A1 _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17072_ _10391_ _10458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14284_ rbzero.debug_overlay.vplaneY\[10\] _08094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16023_ _09564_ _09587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13235_ _07040_ _07049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19455__A2 _12007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_237_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25528__A2 _06311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13166_ _06927_ rbzero.wall_hot\[1\] _06980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13097_ _06910_ _06911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17974_ _11113_ _11115_ _11117_ _11118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19713_ _12473_ _12478_ _12484_ _12485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_TAPCELL_ROW_146_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22062__I1 rbzero.wall_tracer.stepDistY\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16925_ _08018_ _10337_ _10342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_77_i_clk_I clknet_5_29__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16929__I _09139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19644_ _11953_ _11998_ _12415_ _12004_ _12416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_16856_ _10281_ _10282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_189_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_200_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15807_ _09422_ _09423_ _09417_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_200_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19575_ _12180_ _12344_ _12346_ _12347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__14449__I _08226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16787_ _07700_ _10215_ _10219_ _10221_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_13999_ rbzero.tex_r1\[31\] _07807_ _07808_ _07809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13353__I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16992__A3 _10398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18526_ _11577_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15738_ _09370_ _09371_ _09372_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_237_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_201_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18457_ _11537_ _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15669_ rbzero.spi_registers.texadd2\[7\] _09315_ _09321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24267__A2 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__17941__A2 _11071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22278__A1 rbzero.wall_tracer.visualWallDist\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17408_ rbzero.pov.spi_buffer\[56\] _10711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_248_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_18388_ _11498_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_99_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17339_ rbzero.pov.spi_buffer\[39\] _10650_ _10659_ _10660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19908__C _12222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20350_ _01396_ _01444_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_144_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23778__A1 _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19009_ _11879_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20281_ rbzero.wall_tracer.visualWallDist\[3\] _12199_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__19446__A2 rbzero.wall_tracer.rayAddendY\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22020_ _02980_ _03031_ _03035_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22450__A1 rbzero.wall_tracer.texu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23971_ _08810_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold38 net7 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_199_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25710_ _06453_ _06400_ _06494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22922_ _03674_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_26690_ _00600_ clknet_leaf_64_i_clk rbzero.pov.ready_buffer\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20764__A1 _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input18_I i_mode[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25641_ _06377_ _06419_ _06425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22853_ _02651_ _02652_ _03711_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21804_ _02840_ _02842_ _02851_ _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25572_ _06351_ _06352_ _06292_ _06353_ _06355_ _06356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_79_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22784_ _03641_ _03642_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20516__A1 _12706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27311_ _01216_ clknet_leaf_111_i_clk rbzero.traced_texa\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24523_ _05304_ _05306_ _05307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21735_ _02779_ _11123_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_27242_ _01147_ clknet_leaf_82_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24454_ _05116_ _05128_ _05238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_176_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21666_ _11138_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14746__A2 _08528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23405_ _03792_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20617_ _01690_ _01708_ _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_152_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27173_ _01078_ clknet_leaf_50_i_clk rbzero.wall_tracer.rayAddendX\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24385_ _05167_ _05168_ _05126_ _05169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_21597_ _02582_ _02680_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26124_ _00034_ clknet_leaf_252_i_clk rbzero.spi_registers.spi_buffer\[16\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23336_ _04104_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_20548_ _12527_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_132_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Left_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26055_ _06683_ _06622_ _06825_ _06826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_23267_ _04008_ _04006_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20479_ _01496_ _01540_ _01571_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25006_ _05784_ _05789_ _05790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_219_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22218_ _03182_ _03183_ _03191_ _03180_ rbzero.wall_tracer.rcp_fsm.i_data\[9\] _03192_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_23198_ _03817_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_246_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22992__A2 _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22149_ _03114_ _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_238_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_163_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26957_ _00867_ clknet_leaf_182_i_clk rbzero.tex_r1\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14971_ _08743_ reg_gpout\[0\] _08774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_128_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14682__A1 _08379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16710_ _10093_ _10140_ _10152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25908_ _05020_ _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13922_ rbzero.map_overlay.i_otherx\[2\] _06874_ _07733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20755__A1 _12835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17690_ _10889_ _10601_ _10885_ _10891_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_26888_ _00798_ clknet_leaf_176_i_clk rbzero.tex_r0\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XPHY_EDGE_ROW_113_Left_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16641_ _10073_ _10087_ _10088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25839_ _05995_ _06614_ _06623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__14269__I rbzero.debug_overlay.facingX\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13853_ _07607_ _07623_ _07663_ _07477_ _07664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_241_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19360_ _12144_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_187_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16572_ _10022_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_13784_ _07594_ _07595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_202_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_178_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18311_ _11431_ _11447_ _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15523_ _09211_ _09212_ _09202_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19291_ _12105_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_18242_ _11385_ _11386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_44_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15454_ _09160_ _09161_ _09162_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14737__A2 _08526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_215_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_191_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14405_ _07448_ _08214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18173_ _07722_ _11315_ _11251_ rbzero.map_overlay.i_othery\[4\] _11316_ _11317_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_25_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15385_ _08986_ _09111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_122_Left_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_170_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17124_ _10447_ _10497_ _10498_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_52_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14336_ _08124_ _08137_ _08141_ _08145_ _08146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__21483__A2 _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17055_ _10396_ _10445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14267_ _08053_ _08058_ _08026_ _08055_ _08077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_150_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13218_ _07025_ _07026_ _07029_ _07031_ _07032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16006_ _09550_ _09574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22432__A1 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14198_ _07100_ _07988_ _08008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_209_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13348__I _06892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13149_ rbzero.spi_registers.texadd1\[6\] _06916_ _06963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17957_ _11100_ _11101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_131_Left_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16908_ net17 _10177_ _09257_ _10327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17888_ _10997_ _11030_ _11031_ _11032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_164_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19627_ _12316_ _12399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16839_ _10266_ _10261_ _10264_ _10267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13228__A2 _07035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13083__I _06897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19558_ _12176_ _11992_ _12246_ _12329_ _12330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_220_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18167__A2 _11306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18509_ rbzero.tex_r0\[2\] rbzero.tex_r0\[1\] _11566_ _11568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16178__A1 _08959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19489_ _12260_ _12261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__21171__A1 _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21520_ _02599_ _02604_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__15925__A1 rbzero.spi_registers.buf_othery\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13936__B1 _07678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21451_ _02429_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_161_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20402_ _01423_ _01494_ _01495_ _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_24170_ _04904_ _04907_ _04953_ _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21382_ _02068_ _01535_ _02078_ _02066_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_181_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_251_i_clk clknet_5_0__leaf_i_clk clknet_leaf_251_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23121_ _03976_ _03977_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20333_ _12177_ _12325_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13686__C _07496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23052_ _03835_ _03878_ _03833_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20264_ _12867_ _12940_ _13035_ _13036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_45_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14900__A2 _07561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput39 net39 o_rgb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_22003_ rbzero.wall_tracer.size_full\[7\] _03020_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_100_i_clk_I clknet_5_26__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20195_ _12659_ _12967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16653__A2 _08118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26811_ _00721_ clknet_leaf_186_i_clk rbzero.tex_g1\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13467__A2 rbzero.spi_registers.vshift\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26742_ _00652_ clknet_leaf_40_i_clk rbzero.pov.ready_buffer\[72\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23954_ rbzero.wall_tracer.rcp_fsm.operand\[-3\] _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_5_11__f_i_clk_I clknet_3_2_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22905_ rbzero.wall_tracer.trackDistX\[4\] _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23885_ _04684_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18784__I _11713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26673_ _00583_ clknet_leaf_28_i_clk rbzero.pov.ready_buffer\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_168_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25624_ _06050_ _06087_ _06408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22836_ _03691_ _03694_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_224_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_204_i_clk clknet_5_13__leaf_i_clk clknet_leaf_204_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_22767_ _03618_ _03625_ _03626_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25555_ _06034_ _05966_ _06339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_5_10__f_i_clk clknet_3_2_0_i_clk clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24506_ _05284_ _05285_ _05289_ _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_21718_ _11338_ _11424_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25486_ _06269_ _06169_ _06270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22698_ _03231_ _12266_ _03564_ _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_25_i_clk_I clknet_5_20__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_27225_ _01130_ clknet_leaf_110_i_clk rbzero.wall_tracer.stepDistY\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_156_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24437_ _04993_ _04994_ _05214_ _05221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_173_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21649_ _10019_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_23_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15170_ _08946_ _08929_ _08947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_219_i_clk clknet_5_6__leaf_i_clk clknet_leaf_219_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_24368_ _05146_ _05151_ _05075_ _05152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_151_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27156_ _01061_ clknet_leaf_199_i_clk rbzero.map_rom.b6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_105_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14121_ rbzero.tex_r1\[49\] _07930_ _07907_ _07931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23319_ _03860_ _03817_ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26107_ _00017_ clknet_leaf_244_i_clk rbzero.spi_registers.spi_counter\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_27087_ _00997_ clknet_leaf_151_i_clk rbzero.tex_b1\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24299_ _05082_ _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_14052_ _07856_ _07858_ _07860_ _07861_ _07827_ _07862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_104_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26038_ _05027_ _06811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_162_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19564__B _10297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18959__I _11850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22965__A2 _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18860_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] _11781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_246_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24167__A1 _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_219_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17811_ _10965_ _10726_ _10968_ _10970_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__24167__B2 _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17841__A1 _10845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18791_ rbzero.tex_r1\[60\] rbzero.tex_r1\[59\] _11724_ _11728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_246_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13458__A2 rbzero.spi_registers.vshift\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17742_ _10920_ _10655_ _10923_ _10925_ _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_27_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14954_ _07164_ _08755_ _08756_ gpout0.clk_div\[1\] _08757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_234_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13905_ _07703_ _07711_ _07715_ _07716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_17673_ _10875_ rbzero.pov.ready_buffer\[14\] _10880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14885_ rbzero.tex_b1\[46\] _08506_ _08691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_242_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19412_ rbzero.wall_tracer.rayAddendX\[-3\] _12184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_203_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16624_ _09972_ _10071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13836_ rbzero.tex_r0\[28\] _07645_ _07646_ _07647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_217_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15080__A1 _08869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_193_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19343_ _12134_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16555_ rbzero.wall_tracer.rayAddendY\[1\] _10007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13767_ rbzero.tex_r0\[3\] _07577_ _07578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19897__A2 _12668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15506_ _09198_ _09199_ _09191_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19274_ rbzero.tex_b1\[18\] rbzero.tex_b1\[17\] _12094_ _12096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16486_ _08107_ _09942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__26092__A1 rbzero.wall_tracer.rcp_fsm.o_data\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13698_ _07508_ _07509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_230_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18225_ rbzero.map_overlay.i_mapdx\[4\] _07742_ _11369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_96_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15437_ _09147_ _09148_ _09149_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_96_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24642__A2 _05425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18156_ _11255_ _11300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_15368_ rbzero.floor_leak\[1\] _09090_ _09098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17107_ rbzero.pov.ready_buffer\[21\] _10485_ _10486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14319_ rbzero.debug_overlay.vplaneX\[-7\] _08129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_124_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18087_ _11180_ _11228_ _11230_ _11231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_41_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15299_ rbzero.spi_registers.buf_othery\[3\] _09045_ _09048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17038_ _10374_ _10432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16883__A2 _10305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22405__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17773__I _09034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22612__C _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_245_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18085__B2 _11175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20967__A1 _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25990__I _06768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16635__A2 _09928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_209_Left_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18989_ rbzero.tex_g0\[30\] rbzero.tex_g0\[29\] _11866_ _11868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14646__A1 _07889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23905__A1 _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22708__A2 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20719__A1 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_219_Right_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__19585__A1 rbzero.wall_tracer.visualWallDist\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_178_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20951_ _01899_ _02038_ _02039_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_1_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23670_ _04514_ _04521_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20882_ _01971_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14949__A2 _08751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15071__A1 _08809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22621_ rbzero.wall_tracer.texu\[1\] rbzero.texu_hot\[1\] _03476_ _03502_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25340_ _06025_ _06089_ _06123_ _06124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_146_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22552_ _11293_ _03449_ _03450_ rbzero.traced_texa\[0\] _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_218_Left_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__22854__I _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21503_ _02586_ _02493_ _02587_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25271_ _06053_ _06054_ _06055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_199_i_clk_I clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22483_ _03411_ _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_190_i_clk clknet_5_12__leaf_i_clk clknet_leaf_190_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_185_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24222_ _05005_ _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_27010_ _00920_ clknet_leaf_189_i_clk rbzero.tex_g0\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_21434_ _02419_ _02430_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_20_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24153_ _04930_ _04932_ _04934_ _04917_ _04936_ _04937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__14372__I _08181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16323__A1 rbzero.spi_registers.buf_texadd2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21365_ _02402_ _02432_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24397__A1 _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23104_ _03858_ _03875_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20316_ _12410_ _12296_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14305__C _08114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24084_ _04867_ _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16874__A2 _10297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21296_ _02231_ _02236_ _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_251_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23035_ rbzero.wall_tracer.trackDistX\[5\] _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_219_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20247_ rbzero.wall_tracer.size\[10\] _12911_ _12912_ _13019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_9_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_227_Left_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_219_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20178_ _12949_ _12950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16299__I _09761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25897__A1 _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_216_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_204_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24986_ net51 _05768_ _05769_ _05770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19576__A1 rbzero.wall_tracer.size\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26725_ _00635_ clknet_leaf_34_i_clk rbzero.pov.ready_buffer\[55\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23937_ _04739_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19403__I rbzero.wall_tracer.side vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20549__I _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26656_ _00566_ clknet_leaf_156_i_clk rbzero.tex_b0\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14670_ _07928_ _08466_ _08477_ _08478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xclkbuf_leaf_143_i_clk clknet_5_15__leaf_i_clk clknet_leaf_143_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_23868_ _04693_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_169_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25607_ _06386_ _06390_ _06391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_212_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13621_ rbzero.row_render.side _07432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22819_ _02631_ _02637_ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21135__A1 _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_236_Left_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_200_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26587_ _00497_ clknet_leaf_34_i_clk rbzero.pov.spi_buffer\[56\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23799_ _11162_ _03065_ _04634_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_39_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16340_ _08915_ _09820_ _09826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25538_ _06161_ _06164_ _06311_ _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_54_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13552_ rbzero.row_render.size\[4\] _07363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19559__B _12330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26074__A1 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_212_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_171_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_158_i_clk clknet_5_10__leaf_i_clk clknet_leaf_158_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13483_ rbzero.texV\[4\] _07285_ _07294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16271_ rbzero.spi_registers.buf_texadd2\[9\] _09769_ _09774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25469_ _06019_ _06251_ _06253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_212_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14168__A3 _07195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18010_ _11149_ _11153_ _11154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27208_ _01113_ clknet_leaf_79_i_clk rbzero.wall_tracer.stepDistY\[-7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15222_ rbzero.spi_registers.spi_buffer\[17\] _08975_ _08989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18303__A2 _07160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15153_ _08932_ _08933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_105_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27139_ _01049_ clknet_leaf_43_i_clk rbzero.wall_tracer.rayAddendY\[-9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_91_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14104_ _07905_ _07908_ _07911_ _07912_ _07913_ _07914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_91_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19961_ _12732_ _12733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15084_ _08875_ _08876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_245_Left_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14035_ _07483_ _07845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18912_ _11819_ _11821_ _11822_ _11823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_19892_ _12211_ _12224_ _12664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_120_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19803__A2 _12271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18843_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] _11766_ _11767_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__15327__B _09066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13626__I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18774_ _11718_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15986_ _08977_ _09551_ _09559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_223_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_240_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19567__A1 rbzero.wall_tracer.visualWallDist\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17725_ _10912_ _10637_ _10908_ _10914_ _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_240_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14937_ _08742_ net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16937__I rbzero.debug_overlay.playerY\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17656_ _10866_ rbzero.pov.ready_buffer\[8\] _10869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14868_ rbzero.tex_b1\[4\] _07595_ _08674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_230_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24312__A1 _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16607_ _10039_ _10040_ _10047_ _10049_ _10055_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_13819_ _07520_ _07630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21126__A1 _12685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17587_ _10824_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14799_ _08603_ _08604_ _08605_ _08606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_86_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24863__A2 _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19326_ _12114_ _12125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16538_ rbzero.wall_tracer.rayAddendY\[0\] _09991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__26065__A1 _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19257_ rbzero.tex_b1\[11\] rbzero.tex_b1\[10\] _12083_ _12086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16469_ _09925_ _09926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15356__A2 _09088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18208_ _11332_ _11333_ _11302_ _11112_ _11352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_171_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19188_ rbzero.wall_tracer.mapY\[6\] _12016_ _12032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_247_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18139_ rbzero.wall_tracer.visualWallDist\[5\] _11283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__16305__A1 _08997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21150_ _02113_ _02237_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20101_ _12654_ _12871_ _12872_ _12873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_22_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21081_ _02040_ _02166_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13340__1 clknet_leaf_225_i_clk net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_6_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20032_ _12802_ _12803_ _12804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_226_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16608__A2 _08110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14619__A1 _07868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24840_ _05621_ _05622_ _05624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14095__A2 _07641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25225__I _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_i_clk clknet_5_23__leaf_i_clk clknet_leaf_60_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_21983_ rbzero.wall_tracer.rcp_fsm.o_data\[0\] _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_24771_ _05501_ _05540_ _05555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_241_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13842__A2 _07583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26510_ _00420_ clknet_leaf_60_i_clk rbzero.debug_overlay.vplaneX\[-1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23722_ _11196_ _04554_ _04567_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18230__A1 _09056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20934_ _02007_ _02010_ _02023_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_120_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15044__A1 _08831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23106__A2 _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26441_ _00351_ clknet_leaf_54_i_clk rbzero.wall_tracer.rayAddendY\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20865_ _01948_ _01952_ _01953_ _01954_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_138_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23653_ _04377_ _04380_ _04504_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16792__A1 rbzero.pov.ready_buffer\[66\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23657__A3 _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_75_i_clk clknet_5_31__leaf_i_clk clknet_leaf_75_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22604_ _03489_ _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23584_ _04400_ _04317_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26372_ _00282_ clknet_leaf_252_i_clk rbzero.spi_registers.buf_texadd1\[16\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__21668__A2 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20796_ _01796_ _01886_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22535_ _03437_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25323_ _06067_ _06068_ _06107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_193_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20340__A2 _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25254_ _05809_ _05810_ _06038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22466_ _03402_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24205_ _04974_ _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_21417_ _02501_ _02502_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25185_ _05237_ _05968_ _05969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22093__A2 _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22397_ _03342_ _12056_ _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24136_ _04881_ _04920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_60_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21348_ _02397_ _02434_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__24304__I _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14858__B2 _08294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_13_i_clk clknet_5_5__leaf_i_clk clknet_leaf_13_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_131_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24067_ _04850_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_102_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23042__A1 _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21279_ _02359_ _02365_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__18302__I rbzero.hsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23018_ _03856_ _03858_ _03875_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_168_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23593__A2 _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15840_ rbzero.spi_registers.buf_sky\[2\] _09439_ _09449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_28_i_clk clknet_5_20__leaf_i_clk clknet_leaf_28_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_204_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15771_ rbzero.spi_registers.texadd3\[9\] _09396_ _09397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24969_ _05637_ _05685_ _05748_ _05752_ _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__13833__A2 _07626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15661__I _09302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17510_ _10758_ _10780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14722_ _07509_ _08529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26708_ _00618_ clknet_leaf_61_i_clk rbzero.pov.ready_buffer\[38\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_18490_ _11556_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22695__S _11400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17441_ rbzero.pov.spi_buffer\[65\] _10732_ _10729_ _10736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_200_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14653_ rbzero.tex_g1\[61\] _07807_ _08461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26639_ _00549_ clknet_leaf_171_i_clk rbzero.tex_b0\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_197_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13604_ rbzero.row_render.size\[10\] _07360_ _07384_ _07414_ _06883_ _07415_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__19021__I0 rbzero.tex_g0\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17372_ rbzero.pov.spi_buffer\[47\] _10684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14584_ rbzero.tex_g1\[27\] _07597_ _08392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19721__A1 _12489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19111_ _08159_ rbzero.wall_tracer.rayAddendY\[8\] _11955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16323_ rbzero.spi_registers.buf_texadd2\[23\] _09802_ _09812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16492__I rbzero.wall_tracer.rayAddendY\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13535_ rbzero.floor_leak\[3\] _07329_ _07333_ rbzero.floor_leak\[2\] _07345_ _07346_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_40_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19042_ _11892_ _11898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_180_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16254_ _09761_ _09762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_180_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13466_ _07272_ _07276_ _07277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14010__A2 _07818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15205_ _08916_ _08975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_188_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16185_ _09675_ _09709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_188_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13397_ _06877_ _07188_ _07208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20095__A1 _12665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15136_ _08917_ _08918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21831__A2 _09921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__26613__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19944_ _12502_ _12284_ _12716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15067_ rbzero.spi_registers.spi_counter\[0\] _08853_ _08860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_71_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_225_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24376__A4 _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_225_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_242_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14018_ _07817_ _07820_ _07824_ _07826_ _07827_ _07828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_clkbuf_leaf_147_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19875_ _12646_ _12647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18826_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] _11750_ _11753_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18757_ rbzero.tex_r1\[45\] rbzero.tex_r1\[44\] _11708_ _11709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15969_ rbzero.spi_registers.buf_vinf _09545_ _09478_ _09546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_203_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17708_ _10896_ _10623_ _10899_ _10902_ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_72_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18688_ _11669_ _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_102_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_216_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17639_ _10856_ _10857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13588__A1 _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20650_ _01574_ _01575_ _01581_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__19012__I0 rbzero.tex_g0\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19712__A1 _12402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19309_ rbzero.tex_b1\[33\] rbzero.tex_b1\[32\] _12115_ _12116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15520__B _09202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20581_ _01669_ _01672_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__20322__A2 _12584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22320_ _11164_ _03275_ _03276_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22251_ _03202_ _03217_ _03219_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_182_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20086__A1 _12761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21202_ _02179_ _02289_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13760__A1 _07555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22182_ _03161_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_223_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_21133_ _02203_ _02220_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_218_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13694__C _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26990_ _00900_ clknet_leaf_131_i_clk rbzero.tex_g0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_100_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25941_ _05995_ _06614_ _06722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21064_ _12713_ _01466_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20015_ _12431_ _12787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25872_ _06634_ _06644_ _06655_ _05021_ _06656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_24823_ _05420_ _05607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__21338__A1 _12299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15481__I _09067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24754_ _05463_ _05481_ _05482_ _05538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_154_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15017__A1 _08807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21966_ rbzero.wall_tracer.size\[2\] _02992_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19951__A1 _12721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23705_ _03544_ _04552_ _04533_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20917_ _01995_ _02006_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14097__I _07492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13215__B _07028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24288__B1 _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24685_ _05385_ _05372_ _05469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_166_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21897_ _02936_ _02938_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26424_ _00334_ clknet_leaf_249_i_clk rbzero.spi_registers.buf_texadd3\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20848_ _12483_ _12647_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23636_ _04397_ _04391_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20827__I _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14240__A2 _08045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26355_ _00265_ clknet_leaf_245_i_clk rbzero.spi_registers.buf_texadd0\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14825__I _07563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23567_ _04416_ _04419_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20779_ _01760_ _01762_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25306_ _06010_ _06089_ _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13320_ _07127_ _07132_ _07133_ _07134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_22518_ rbzero.wall_tracer.texu\[3\] _03429_ _03430_ _07452_ _03433_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_23498_ rbzero.wall_tracer.stepDistX\[9\] _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26286_ _00196_ clknet_leaf_230_i_clk rbzero.spi_registers.buf_sky\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17190__A1 _10538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24055__A3 _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25237_ _06020_ _05974_ _06021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13251_ _07040_ _07065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22449_ _03351_ _03389_ _03390_ _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15740__A2 _09373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13182_ _06990_ _06995_ _06996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_25168_ _05951_ _05920_ _05840_ _05952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24119_ _04730_ _04724_ _04718_ _04819_ _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_20_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25099_ _05882_ _05883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17990_ _11133_ _11134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_183_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16941_ rbzero.pov.ready_buffer\[55\] _10288_ _10329_ _10355_ _10356_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_159_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19660_ _12431_ _12432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_148_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16872_ _08028_ rbzero.debug_overlay.playerY\[-9\] _10296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18611_ _11625_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_220_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15823_ rbzero.spi_registers.texadd3\[23\] _09032_ _09435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19591_ _12289_ _11994_ _12290_ _12362_ _12363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_220_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18542_ _11564_ _11586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_220_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15754_ _09381_ _09382_ _09384_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15008__A1 _08807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__19942__A1 _12713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14705_ rbzero.tex_b0\[59\] _08252_ _08512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_197_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18473_ rbzero.tex_g1\[51\] rbzero.tex_g1\[50\] _11544_ _11547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_158_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14936__S _07185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15559__A2 _09230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15685_ rbzero.spi_registers.buf_texadd2\[11\] _09328_ _09333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17424_ rbzero.pov.spi_buffer\[60\] _10723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__22438__B _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14636_ rbzero.tex_g1\[43\] _07625_ _08444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17355_ rbzero.pov.spi_buffer\[43\] _10662_ _10671_ _10672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16508__A1 _09927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14567_ _08370_ _08372_ _08375_ _08376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13779__C _07589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_73_i_clk_I clknet_5_29__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16306_ _09798_ _09799_ _09795_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13518_ _07328_ _07329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17286_ _10617_ _10619_ _10620_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14498_ _07814_ _08305_ _08306_ _08307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__17181__A1 _10538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19025_ _11888_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_153_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16237_ _09591_ _09748_ _09749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13449_ rbzero.traced_texVinit\[9\] _07259_ _07260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_23_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16168_ _09671_ _09696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18130__B1 _11249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24429__S1 _05212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15119_ rbzero.spi_registers.mosi _08903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14470__I _07835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16099_ _09642_ _09643_ _09637_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19927_ _12698_ _12699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_205_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19858_ _12628_ _12629_ _12630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_138_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18809_ _11738_ _11739_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19789_ _12560_ _12561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_183_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16995__A1 _10345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_21820_ _11077_ _02696_ _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21751_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.wall_tracer.rayAddendX\[-5\] _02800_
+ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_159_Left_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__22348__B _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20702_ _01791_ _01792_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24470_ _05253_ _05205_ _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_21682_ _11133_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_191_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20633_ _11387_ _01532_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23421_ _04151_ _04157_ _04159_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__22296__A2 _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23352_ _04201_ _04206_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_26140_ _00050_ clknet_leaf_215_i_clk rbzero.map_overlay.i_othery\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20564_ _01567_ _01656_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_33_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22303_ rbzero.wall_tracer.trackDistY\[0\] _03254_ _03262_ _03263_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__17956__I _11099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26071_ _06823_ _06789_ _06756_ _06840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23283_ _04083_ _04088_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_115_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24442__B1 _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20495_ _01504_ _01505_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_61_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23894__S _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22234_ _11248_ _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25022_ _05802_ _05803_ _05805_ _05806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_132_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_168_Left_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22165_ _11985_ _03121_ _03093_ _11068_ _03148_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_100_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23693__I _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21116_ _02087_ _02088_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22096_ _03082_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26973_ _00883_ clknet_leaf_123_i_clk rbzero.texV\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_234_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17691__I _10884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25924_ _06696_ _06701_ _06705_ _06706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_21047_ _12210_ _01994_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_245_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15238__A1 _09000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25855_ _06514_ _06545_ _06639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_226_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24806_ _05523_ _05535_ _05590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__16100__I _09595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25786_ _06552_ _06569_ _06570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22998_ _03843_ _03847_ _03855_ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_126_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_177_Left_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24737_ _05464_ _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21949_ rbzero.wall_tracer.size_full\[-11\] _02986_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16738__A1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21731__A1 _11344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27456_ _01361_ clknet_leaf_72_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15470_ rbzero.spi_registers.texadd0\[4\] _09163_ _09173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24668_ _05434_ _05451_ _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_194_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26407_ _00317_ clknet_leaf_245_i_clk rbzero.spi_registers.buf_texadd3\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14421_ rbzero.tex_g0\[22\] _08227_ _08229_ _08230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23619_ _04368_ _04370_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27387_ _01292_ clknet_leaf_100_i_clk rbzero.wall_tracer.trackDistY\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24599_ _05370_ _05381_ _05383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23868__I _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19152__A2 _11991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17140_ _10145_ _10485_ _10509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14352_ rbzero.debug_overlay.facingY\[-4\] _08162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26338_ _00248_ clknet_leaf_238_i_clk rbzero.spi_registers.buf_texadd0\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__19567__B _12245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13303_ _07049_ _07113_ _07116_ _07057_ _07117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_108_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17071_ _10456_ _10457_ _10436_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14283_ _08074_ _08092_ _08093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_26269_ _00179_ clknet_leaf_17_i_clk rbzero.spi_registers.texadd3\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_186_Left_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16022_ _09518_ _09585_ _09586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13234_ _07019_ _07023_ _07048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_0__f_i_clk_I clknet_3_0_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21798__A1 _10477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15386__I _09111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14290__I rbzero.debug_overlay.vplaneY\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17466__A2 _10544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13165_ _06934_ _06978_ _06979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13096_ _06909_ _06910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17973_ _11116_ _11099_ _11117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_237_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19712_ _12402_ _12483_ _12484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16924_ _08018_ _10337_ _10341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__15229__A1 _08994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23108__I _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19643_ _10310_ _12415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16855_ _10280_ _10163_ _09028_ _10281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_233_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21970__A1 _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20773__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_195_Left_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_189_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15806_ rbzero.spi_registers.buf_texadd3\[18\] _09420_ _09423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_220_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19574_ _12345_ _11993_ _12346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_200_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16786_ _10220_ _10221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_232_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_200_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13998_ _07520_ _07808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__19915__A1 _12684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14452__A2 _08258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23711__A2 _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18525_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _11576_ _11577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15737_ _09336_ _09372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_237_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16945__I _07681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_237_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20525__A2 _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18456_ rbzero.tex_g1\[44\] rbzero.tex_g1\[43\] _11533_ _11537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15668_ _09319_ _09320_ _09314_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_185_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24267__A3 _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17407_ _10708_ _10700_ _10710_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17941__A3 _11073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14619_ _07868_ _08423_ _08426_ _08427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__22278__A2 _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18387_ rbzero.tex_g1\[14\] rbzero.tex_g1\[13\] _11496_ _11498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15599_ rbzero.spi_registers.texadd1\[13\] _09268_ _09269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20289__A1 _12235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17338_ _10658_ _10659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_248_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17269_ _10605_ _10606_ _10607_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15704__A2 _09340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16901__A1 rbzero.pov.ready_buffer\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19008_ rbzero.tex_g0\[38\] rbzero.tex_g0\[37\] _11877_ _11879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20280_ _12962_ _12976_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21789__B2 _09918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14414__B _08222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14133__C _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22202__A2 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23970_ rbzero.wall_tracer.rcp_fsm.i_data\[0\] _04755_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_194_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold39 net97 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_209_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_208_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14691__A2 _08496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22921_ _03777_ _03778_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23950__A2 _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21961__A1 _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25640_ _06373_ _06422_ _06423_ _06424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_22852_ _02650_ _02653_ _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_211_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23702__A2 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21803_ _08132_ _08144_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25571_ _06157_ _06354_ _06293_ _06355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_196_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22783_ _02617_ _02640_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20516__A2 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21713__A1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27310_ _01215_ clknet_leaf_112_i_clk rbzero.traced_texa\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24522_ _05129_ _05305_ net77 _05306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_38_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21734_ _11108_ _11122_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_213_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27241_ _01146_ clknet_leaf_82_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24453_ _05236_ _05237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21665_ _02730_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_136_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23404_ _04256_ _04257_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20616_ _01698_ _01707_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_164_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27172_ _01077_ clknet_leaf_50_i_clk rbzero.wall_tracer.rayAddendX\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24384_ _04720_ _05047_ _05168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17145__A1 _09035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21596_ _02582_ _02680_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_35_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26123_ _00033_ clknet_leaf_4_i_clk rbzero.spi_registers.spi_buffer\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23335_ _04146_ _04189_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20547_ _01629_ _01639_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17696__A2 rbzero.pov.ready_buffer\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18893__A1 rbzero.traced_texa\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26054_ _06697_ _06723_ _06825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23266_ _03491_ _04013_ _04121_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_20478_ _01498_ _01539_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25005_ _05787_ _05788_ _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22217_ _03177_ _03190_ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23197_ _03811_ _04052_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22441__A2 _07704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22148_ _03090_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_163_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15934__I _09504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_21_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22079_ _03024_ _03034_ _03075_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26956_ _00866_ clknet_leaf_182_i_clk rbzero.tex_r1\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14970_ _08747_ net96 _08772_ _08773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_128_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14682__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25907_ _06686_ _06687_ _06689_ _06667_ _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13921_ rbzero.map_overlay.i_othery\[4\] _07732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_96_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26887_ _00797_ clknet_leaf_175_i_clk rbzero.tex_r0\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_107_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20755__A2 _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16640_ _10086_ _10087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25838_ _06621_ _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13852_ _07624_ _07650_ _07662_ _07663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_202_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25694__A2 _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14434__A2 _08206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16571_ _09944_ _10022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25769_ _06526_ _06537_ _06553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13783_ _07419_ _07594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16765__I _10178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14985__A3 _07712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18310_ _07181_ _11445_ _11446_ _11447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_186_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15522_ rbzero.spi_registers.buf_texadd0\[17\] _09209_ _09212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19290_ rbzero.tex_b1\[25\] rbzero.tex_b1\[24\] _12104_ _12105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_246_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18241_ _11384_ _11385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_27439_ _01344_ clknet_leaf_72_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15453_ _09111_ _09162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_61_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22716__B _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14404_ _08208_ _08212_ _07465_ _08213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_191_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18172_ rbzero.map_overlay.i_othery\[3\] _11256_ _11316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_182_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15384_ rbzero.spi_registers.buf_leak\[5\] _09103_ _09110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17123_ rbzero.pov.ready_buffer\[3\] _10379_ _10498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14335_ _08143_ _08022_ _08046_ _08144_ _08145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__23209__A1 _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22680__A2 _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24957__A1 _05696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17054_ _08149_ _10443_ _10444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14266_ _08075_ _08076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16005_ rbzero.spi_registers.buf_mapdy\[2\] _09572_ _09573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13217_ rbzero.spi_registers.texadd2\[22\] _07027_ _07030_ rbzero.spi_registers.texadd1\[22\]
+ _07031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14197_ _08006_ _08007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_210_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24222__I _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13148_ rbzero.spi_registers.texadd0\[6\] _06962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_57_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24185__A2 _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13079_ _06894_ net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17956_ _11099_ _11100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16907_ _10309_ _10326_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17887_ _08073_ rbzero.wall_tracer.rayAddendX\[8\] _11031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__21943__A1 rbzero.wall_tracer.rcp_done vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13364__I _07175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_221_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19626_ _12397_ _12398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_189_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16838_ _10166_ _10266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_205_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14425__A2 _08233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19557_ _12249_ _11078_ _12329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23696__A1 _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16769_ _10194_ _10205_ _10206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__19051__I _11892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18508_ _11567_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19488_ _12259_ _12260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_186_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23448__A1 _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18439_ _11527_ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21450_ _02525_ _02535_ _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__17127__A1 _06900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20401_ _01425_ _01439_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21381_ _02340_ _02343_ _01726_ _01620_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_32_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22671__A2 _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20332_ _12525_ _13024_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23120_ _03864_ _03874_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23051_ _03904_ _03907_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20263_ _12870_ _12939_ _13035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_101_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22002_ rbzero.wall_tracer.rcp_fsm.o_data\[7\] _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_228_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20194_ _12932_ _12934_ _12965_ _12966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_179_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26810_ _00720_ clknet_leaf_179_i_clk rbzero.tex_g1\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_110_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22187__A1 _11290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_195_i_clk_I clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23971__I _08810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14664__A2 _07460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23923__A2 _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26741_ _00651_ clknet_leaf_40_i_clk rbzero.pov.ready_buffer\[71\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23953_ _04750_ _04751_ _04752_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25125__A1 _05908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22904_ _03618_ _03761_ _03762_ _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_4_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22587__I _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26672_ _00582_ clknet_leaf_34_i_clk rbzero.pov.ready_buffer\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23884_ _12511_ _04686_ _04703_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14416__A2 _08202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25623_ _06084_ _05971_ _06125_ _05720_ _06407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_123_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22835_ _03692_ _03693_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_123_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25554_ _06299_ _06300_ _06337_ _06338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_196_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22766_ rbzero.wall_tracer.trackDistX\[2\] _03605_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24505_ _05286_ _05288_ _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_177_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19896__I _12237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21717_ _10243_ _02773_ _02774_ _02775_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_25485_ _06161_ _06164_ _06269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_52_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22697_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] _03558_
+ _03564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_192_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27224_ _01129_ clknet_leaf_107_i_clk rbzero.wall_tracer.stepDistY\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24436_ _05197_ _05157_ _05162_ _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_156_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13927__B2 _07736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20835__I _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21648_ _08106_ rbzero.wall_tracer.rayAddendY\[-6\] _09910_ _02721_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_35_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22111__A1 _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27155_ _01060_ clknet_leaf_202_i_clk rbzero.map_rom.c6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24367_ _05088_ _05147_ _05150_ _05151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_50_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21579_ _02503_ _02505_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14120_ _07498_ _07930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26106_ _00016_ clknet_leaf_244_i_clk rbzero.spi_registers.spi_counter\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23318_ _03725_ _03815_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27086_ _00996_ clknet_leaf_151_i_clk rbzero.tex_b1\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24298_ _05017_ _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14054__B _07642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26037_ _06802_ _03008_ _06808_ _06809_ _06810_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_14051_ _07825_ _07861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_123_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23249_ _04093_ _04104_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_247_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_203_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14104__B2 _07912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17810_ _10966_ rbzero.pov.ready_buffer\[61\] _10970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18790_ _11727_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22178__A1 _11039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14655__A2 _07804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17741_ _10921_ rbzero.pov.ready_buffer\[37\] _10925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26939_ _00849_ clknet_leaf_184_i_clk rbzero.tex_r1\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14953_ _08754_ _08748_ _08756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_238_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13184__I _06918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13904_ _07709_ _07060_ _07052_ _07699_ _07714_ _07715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_203_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17672_ _10873_ _10585_ _10877_ _10879_ _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14884_ _08684_ _08689_ _08690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14407__A2 _08202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19411_ _12177_ _12183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16623_ _01029_ _10061_ _10070_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13835_ _07524_ _07646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16554_ _09945_ _10005_ _10006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19342_ rbzero.tex_b1\[48\] rbzero.tex_b1\[47\] _12130_ _12134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13766_ _07576_ _07577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_186_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15505_ rbzero.spi_registers.buf_texadd0\[13\] _09194_ _09199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19273_ _12095_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_195_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16485_ _09924_ _09937_ _09941_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_223_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13697_ _07481_ _07508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18224_ _11359_ _11367_ _11299_ _11368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_230_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15436_ _09111_ _09149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_96_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18155_ _11298_ _11299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__14591__A1 _07848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15367_ _09096_ _09097_ _09089_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__18857__A1 _08750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22653__A2 _12214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23850__A1 rbzero.wall_tracer.stepDistY\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_230_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17106_ _10391_ _10485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14318_ _08127_ _08128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18086_ _11166_ _11185_ _11229_ _11230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_15298_ rbzero.map_overlay.i_othery\[3\] _09043_ _09047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13359__I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24380__C _05163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17037_ _10430_ _10431_ _10414_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14249_ _08025_ _08030_ _08059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_7_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14899__B _08214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14894__A2 _08698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_245_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20967__A2 _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18988_ _11867_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22169__B2 _11067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_183_Right_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17939_ rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.rayAddendX\[-2\] _11079_
+ _11082_ _11083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__21916__A1 _10477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25107__A1 _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20950_ _01901_ _02028_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19609_ _12380_ _12381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__23669__A1 rbzero.wall_tracer.stepDistX\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15523__B _09202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20881_ _11389_ _01843_ _01970_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_95_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13822__I _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22620_ _03501_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22551_ _03453_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21502_ _02464_ _02477_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_192_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25270_ _06049_ _06052_ _06054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22482_ _09938_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24221_ _05004_ _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_17_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18848__A1 rbzero.traced_texa\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21433_ _02460_ _02518_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_185_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23841__A1 _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24152_ _04930_ _04836_ _04935_ _04936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_21364_ _02325_ _02438_ _02436_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19665__B _12408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20315_ _12480_ _12258_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23103_ _03858_ _03875_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24083_ _04866_ _04858_ _04859_ _04861_ _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_21295_ _02378_ _02381_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14885__A2 _08506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20246_ rbzero.wall_tracer.size\[10\] _12911_ _13018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_23034_ _03891_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_244_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21080__A1 _09901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20177_ _12760_ _12949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__17823__A2 rbzero.pov.ready_buffer\[66\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14637__A2 _07909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24985_ _05558_ _05592_ _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_150_Right_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26724_ _00634_ clknet_leaf_34_i_clk rbzero.pov.ready_buffer\[54\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23936_ _04727_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_197_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22580__A1 rbzero.wall_tracer.wall\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23206__I _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26655_ _00565_ clknet_leaf_157_i_clk rbzero.tex_b0\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23867_ _04683_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_150_Left_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17204__I _10544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25606_ _06387_ _06388_ _06389_ _06390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_158_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13620_ _07430_ _07431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_22818_ _02628_ _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_175_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26586_ _00496_ clknet_leaf_34_i_clk rbzero.pov.spi_buffer\[55\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23798_ _11164_ rbzero.wall_tracer.stepDistY\[3\] _04631_ _04634_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__21135__A2 _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18387__I0 rbzero.tex_g1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25537_ _06265_ _06314_ _06320_ _06321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13551_ rbzero.row_render.size\[5\] _07362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22749_ _03608_ _03601_ _03609_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26074__A2 _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16011__A1 _08950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16270_ _09770_ _09772_ _09773_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25468_ _06019_ _06251_ _06252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_212_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13482_ rbzero.texV\[3\] _07291_ _07292_ _07293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_212_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27207_ _01112_ clknet_leaf_77_i_clk rbzero.wall_tracer.stepDistY\[-8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15221_ _08982_ _08985_ _08988_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15659__I _09289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24419_ net62 _05202_ _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_136_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25399_ _06181_ _06182_ _06183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__19500__A2 _12271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20646__A1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18303__A3 _06859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15152_ _08931_ _08932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_27138_ _01048_ clknet_leaf_31_i_clk rbzero.wall_tracer.rayAddendX\[-6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14103_ _07495_ _07913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_239_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19960_ _12731_ _12732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15083_ _07204_ _08872_ _08873_ _08874_ _08875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_27069_ _00979_ clknet_leaf_144_i_clk rbzero.tex_b1\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_22_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14876__A2 _08496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14034_ rbzero.tex_r1\[22\] _07843_ _07844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18911_ rbzero.traced_texa\[9\] _07259_ _11822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19891_ _12662_ _12192_ _12663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15394__I _09118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_227_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18842_ _11763_ _11765_ _11766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14628__A2 _07834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23899__A1 _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18773_ rbzero.tex_r1\[52\] rbzero.tex_r1\[51\] _11714_ _11718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15985_ rbzero.spi_registers.buf_mapdx\[3\] _09548_ _09558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_145_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13300__A2 _07111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17724_ _10913_ rbzero.pov.ready_buffer\[31\] _10914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14936_ reg_rgb\[5\] _08741_ _07185_ _08742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_145_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_250_i_clk clknet_5_0__leaf_i_clk clknet_leaf_250_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_188_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14867_ rbzero.tex_b1\[5\] _07890_ _08673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17655_ _10850_ _10868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__17114__I _10491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16606_ _10053_ _10054_ _09899_ _10055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13818_ _07628_ _07629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17586_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _10823_ _10824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14798_ rbzero.tex_b0\[4\] _08247_ _08605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16537_ _08104_ _09990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19325_ _12124_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13749_ _07556_ _07557_ _07558_ _07559_ _07496_ _07560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_57_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16002__A1 _09542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_143_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16468_ _09896_ _09925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_19256_ _12085_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15419_ _09114_ _09135_ _09136_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_18207_ _11347_ _11348_ _11350_ _11334_ _11351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_182_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19187_ _11913_ _12009_ _12030_ _12031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16399_ _09868_ _09869_ _09867_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18138_ rbzero.wall_tracer.visualWallDist\[6\] _11282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_247_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25576__A1 _05949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18069_ rbzero.wall_tracer.trackDistX\[-11\] _11213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20100_ _12615_ _12651_ _12872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14867__A2 _07890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21080_ _09901_ _02167_ _02168_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_186_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13817__I _07340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_203_i_clk clknet_5_13__leaf_i_clk clknet_leaf_203_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_20031_ _12682_ _12797_ _12796_ _12803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__21062__A1 _12300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23735__B _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17805__A2 rbzero.pov.ready_buffer\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__19558__A2 _11992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_9_i_clk clknet_5_1__leaf_i_clk clknet_leaf_9_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_225_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24770_ _05550_ _05553_ _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_21982_ _03008_ _02998_ _03009_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_218_i_clk clknet_5_3__leaf_i_clk clknet_leaf_218_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__22562__A1 _11284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22562__B2 rbzero.traced_texa\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23721_ _04542_ _04566_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20933_ _02013_ _02022_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__18230__A2 _11343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16241__A1 _08913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26440_ _00350_ clknet_leaf_55_i_clk rbzero.wall_tracer.rayAddendY\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23652_ _04378_ _04379_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_20864_ _01726_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_194_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25241__I _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22603_ _03486_ _03488_ _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_49_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26371_ _00281_ clknet_leaf_6_i_clk rbzero.spi_registers.buf_texadd1\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23583_ _04311_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19030__I1 rbzero.tex_g0\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20795_ _01854_ _01885_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25322_ _06069_ _06106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22534_ _03435_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_162_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15479__I _09064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25253_ _06036_ _06037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22465_ _10255_ _11444_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24204_ _04973_ _04988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_162_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21416_ _01925_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_122_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25184_ _05967_ _05968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22396_ _03341_ _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__25567__A1 _06328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24135_ _04918_ _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21347_ _02400_ _02433_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24066_ _04843_ _04849_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_131_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21278_ _02360_ _02364_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_130_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23017_ _03864_ _03874_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20229_ _12999_ _12381_ _12520_ _12491_ _13001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_200_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16480__A1 _09927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19549__A2 _11067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15770_ _09037_ _09396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24968_ _05686_ _05717_ _05751_ _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_169_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14721_ _08276_ _08528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_23919_ _08813_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26707_ _00617_ clknet_leaf_61_i_clk rbzero.pov.ready_buffer\[37\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24899_ _05651_ _05680_ _05682_ _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_169_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17440_ _10712_ _10735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14652_ _08455_ _08456_ _08458_ _08459_ _07935_ _08460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_26638_ _00548_ clknet_leaf_149_i_clk rbzero.tex_b0\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__22305__A1 _11293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17980__A1 _11107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16783__A2 _10217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13603_ _07408_ _07410_ _07413_ _07414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14794__A1 _07462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17371_ _10681_ _10677_ _10683_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_156_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14583_ _08387_ _08388_ _08390_ _07826_ _07827_ _08391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26569_ _00479_ clknet_leaf_64_i_clk rbzero.pov.spi_buffer\[38\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19110_ _11953_ _11954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16322_ _09810_ _09811_ _09807_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13534_ _07342_ _07344_ _07345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15389__I _09113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19041_ _11897_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13349__A2 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16253_ _09659_ _09761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_125_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13465_ _07273_ _07274_ _07275_ _07276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_153_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22724__B _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15204_ _08972_ _08974_ _08971_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_211_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16184_ rbzero.spi_registers.buf_texadd1\[12\] _09707_ _09708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13396_ gpout0.hpos\[8\] _07207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_188_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21292__A1 _12691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15135_ _08916_ _08917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19943_ _12276_ _12692_ _12715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15066_ _08853_ _08858_ _08859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24431__S _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24230__A1 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_242_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21044__A1 _12668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13637__I _07443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14017_ _07449_ _07827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_120_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_242_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19874_ _12645_ _12646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__25326__I _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18825_ _11737_ _11752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_207_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18756_ _11692_ _11708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_223_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15968_ _09458_ _09544_ _09545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_175_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17707_ _10897_ rbzero.pov.ready_buffer\[26\] _10902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_188_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14919_ _07624_ _08719_ _08724_ _08725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_69_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15899_ _08942_ _09476_ _09493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18687_ rbzero.tex_r1\[15\] rbzero.tex_r1\[14\] _11666_ _11669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_102_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17638_ rbzero.pov.spi_done _10856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17971__A1 rbzero.map_rom.f4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14785__A1 _07912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17569_ rbzero.tex_b0\[42\] rbzero.tex_b0\[41\] _10812_ _10814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_147_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19308_ _12114_ _12115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20580_ _01643_ _01670_ _01671_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19239_ rbzero.tex_b1\[3\] rbzero.tex_b1\[2\] _12073_ _12076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22250_ rbzero.wall_tracer.visualWallDist\[-9\] _03218_ _03211_ _03219_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23272__A2 _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21283__A1 _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21201_ _02243_ _02288_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22181_ _12005_ _03120_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_142_i_clk clknet_5_14__leaf_i_clk clknet_leaf_142_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_21132_ _02205_ _02219_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_113_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21035__A1 _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22083__I0 rbzero.wall_tracer.rcp_fsm.o_data\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25940_ _06702_ _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21063_ _12683_ _01631_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20014_ _12778_ _12784_ _12785_ _12786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25871_ _05027_ _06654_ _06655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__17463__B _10751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_157_i_clk clknet_5_10__leaf_i_clk clknet_leaf_157_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__19234__I _12072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24822_ _05413_ _05605_ _05606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_216_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24753_ _05481_ _05482_ _05463_ _05537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_240_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21965_ _02983_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_167_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23704_ _04549_ _04550_ _04551_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19951__A2 _12722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_20916_ _01998_ _02005_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24684_ _05465_ _05467_ _05468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24288__B2 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21896_ _02920_ _08138_ _02937_ _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_26423_ _00333_ clknet_leaf_251_i_clk rbzero.spi_registers.buf_texadd3\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23635_ _04376_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_193_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20847_ _01817_ _01818_ _01936_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26354_ _00264_ clknet_leaf_249_i_clk rbzero.spi_registers.buf_texadd0\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23566_ _04417_ _04418_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20778_ _01860_ _01868_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16517__A2 _08869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25305_ _06088_ _06089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_147_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14528__A1 rbzero.tex_g0\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22517_ _03432_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26285_ _00195_ clknet_leaf_227_i_clk rbzero.spi_registers.buf_sky\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23497_ _11410_ _04349_ _04350_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25236_ _05728_ _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_190_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13250_ _07063_ _07064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__19467__A1 _12224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22448_ _03345_ _03389_ _03347_ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__24460__A1 _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24315__I _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24460__B2 _05133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20077__A2 _12224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25167_ _05336_ _05951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_150_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13751__A2 _07561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13181_ _06991_ _06993_ _06994_ _06995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22379_ _03320_ _10193_ _03324_ _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24118_ _04806_ _04901_ _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_237_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25098_ _05879_ _05881_ _05882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24049_ rbzero.wall_tracer.rcp_fsm.operand\[6\] _04832_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_16940_ _10353_ _10354_ _10275_ _10355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_183_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16871_ _10170_ _10295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_148_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18610_ rbzero.tex_r0\[46\] rbzero.tex_r0\[45\] _11623_ _11625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15822_ _09433_ _09434_ _09430_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_220_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19590_ _12248_ _11081_ _12362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17092__C _09441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22526__A1 _12834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18541_ _11585_ _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15753_ _09383_ _09384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14288__I rbzero.debug_overlay.vplaneY\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14704_ _08264_ _08503_ _08510_ _08511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_158_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18472_ _11546_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15684_ rbzero.spi_registers.texadd2\[11\] _09326_ _09332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14635_ rbzero.tex_g1\[41\] _07906_ _07907_ _08443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17423_ _10720_ _10713_ _10722_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14566_ _08374_ net2 _08375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17354_ _10658_ _10671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_16_i_clk_I clknet_5_4__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16305_ _08997_ _09793_ _09799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13517_ _07323_ _07327_ _07328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__14519__A1 _08316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17285_ rbzero.pov.spi_buffer\[25\] _10615_ _10612_ _10620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16008__I _09564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14497_ rbzero.tex_g0\[41\] _07898_ _08306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16236_ _09747_ _09748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19024_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _11887_ _11888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13448_ rbzero.texV\[9\] _07259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_153_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14751__I _07917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16167_ _09694_ _09695_ _09689_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13379_ gpout0.vpos\[2\] _07190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15118_ _08894_ _08902_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_239_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16098_ _08983_ _09635_ _09643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21017__A1 _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13367__I _07178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22065__I0 rbzero.wall_tracer.rcp_fsm.o_data\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19926_ _12593_ _12698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15049_ _08839_ _08841_ _08842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_74_i_clk clknet_5_29__leaf_i_clk clknet_leaf_74_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19857_ _12260_ _12496_ _12527_ _12569_ _12629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_18808_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] _11735_ _11739_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_208_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19788_ _12479_ _12560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_223_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_89_i_clk clknet_5_24__leaf_i_clk clknet_leaf_89_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_211_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18739_ rbzero.tex_r1\[37\] rbzero.tex_r1\[36\] _11698_ _11699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_84_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21750_ _08131_ rbzero.wall_tracer.rayAddendX\[-5\] _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__17944__A1 _08073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20701_ _01746_ _01751_ _01753_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12_i_clk clknet_5_6__leaf_i_clk clknet_leaf_12_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_21681_ _12019_ _12021_ _12022_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__13830__I _07341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23420_ _04155_ _04163_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_20632_ _12303_ _01723_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23351_ _04202_ _04205_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20563_ _01570_ _01655_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22364__B rbzero.wall_tracer.wall\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22302_ _11181_ _03239_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26070_ _06785_ _06836_ _06838_ _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15183__A1 _08957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_27_i_clk clknet_5_20__leaf_i_clk clknet_leaf_27_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_116_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23282_ _04135_ _04136_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_115_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24293__I1 _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24442__A1 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20494_ _01585_ _01586_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24442__B2 _05225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25021_ _05546_ _05596_ _05804_ _05805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__15757__I _09352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22233_ _03203_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13733__A2 _07543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_30__f_i_clk_I clknet_3_7_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18121__A1 _07694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22164_ _11286_ _03104_ _03136_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__17972__I rbzero.map_rom.f2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21115_ _02187_ _02202_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_246_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__25942__A1 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22095_ _08374_ _12164_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26972_ _00882_ clknet_leaf_124_i_clk rbzero.texV\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_165_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25923_ _06703_ _06704_ _06705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21046_ _01999_ _02004_ _02134_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_214_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25854_ _06637_ _06638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22508__A1 rbzero.wall_tracer.size\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24805_ net61 _05585_ _05588_ _05589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_199_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25785_ _06553_ _06556_ _06568_ _06569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_202_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14997__B2 _07180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22997_ _03848_ _03854_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_186_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24736_ _04919_ _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21948_ _02985_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17935__A1 _08084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27455_ _01360_ clknet_leaf_71_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24667_ _05438_ _05450_ _05451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__26612__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21879_ _02921_ _02904_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13740__I _07331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17212__I _10564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26406_ _00316_ clknet_leaf_246_i_clk rbzero.spi_registers.buf_texadd3\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14420_ rbzero.tex_g0\[23\] _07832_ _08229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_154_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23618_ _04435_ _04438_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19688__A1 _12425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27386_ _01291_ clknet_leaf_101_i_clk rbzero.wall_tracer.trackDistY\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__24681__A1 _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24598_ _05381_ _05370_ _05382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_37_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19152__A3 _11992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14351_ rbzero.debug_overlay.facingY\[-5\] _08161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26337_ _00247_ clknet_leaf_238_i_clk rbzero.spi_registers.buf_texadd0\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23549_ _04312_ _04315_ _04401_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13302_ _07114_ _07115_ _07049_ _07116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17070_ rbzero.pov.ready_buffer\[13\] _10434_ _10457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14282_ _08076_ _08078_ _08091_ _08092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26268_ _00178_ clknet_leaf_21_i_clk rbzero.spi_registers.texadd3\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24433__A1 _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13185__B1 _06992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16021_ _09550_ _09585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25219_ _05388_ _06003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_33_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13233_ _07033_ _07043_ _07046_ _07047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14921__A1 _08201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26199_ _00109_ clknet_leaf_10_i_clk rbzero.spi_registers.texadd0\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22995__B2 _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13164_ _06936_ _06977_ _06978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19583__B _12310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_1__f_i_clk clknet_3_0_0_i_clk clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_242_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13095_ _06908_ rbzero.wall_hot\[1\] _06909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17972_ rbzero.map_rom.f2 _11116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__20522__B _12182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19711_ _12482_ _12483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16923_ _10236_ _10334_ _10340_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__19612__A1 _12383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20222__A2 _12273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19642_ _12413_ _12414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__23833__B _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16854_ net17 _10280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_232_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15805_ rbzero.spi_registers.texadd3\[18\] _09418_ _09422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19573_ rbzero.wall_tracer.side _12345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__14988__A1 _07164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_200_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13997_ _07518_ _07807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16785_ _07166_ _10220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_204_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19602__I rbzero.wall_tracer.stepDistX\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_200_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18524_ _11565_ _11576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15736_ rbzero.spi_registers.buf_texadd3\[0\] _09364_ _09371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13660__A1 rbzero.row_render.texu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_237_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17926__A1 _08079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18455_ _11536_ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15667_ rbzero.spi_registers.buf_texadd2\[6\] _09317_ _09320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13650__I _07460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17406_ rbzero.pov.spi_buffer\[56\] _10709_ _10706_ _10710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_233_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14618_ _07842_ _08424_ _08425_ _08426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__19679__A1 _12355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15598_ _09254_ _09268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13412__A1 _07195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18386_ _11497_ _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__18726__I0 rbzero.tex_r1\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20289__A2 _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13963__A2 _07772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14549_ _08201_ _08314_ _08356_ _08357_ _08358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_56_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17337_ _06897_ _10658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15165__A1 _08942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24424__A1 _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17268_ rbzero.pov.spi_buffer\[21\] _10603_ _10599_ _10607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19007_ _11878_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16219_ _09731_ _09733_ _09734_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17199_ _10546_ _10555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21789__A2 _09977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19909_ _12678_ _12679_ _12680_ _12681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_227_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15526__B _09202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13825__I _07524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22920_ _03676_ _03699_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_242_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_22851_ _12760_ _03709_ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19512__I _12283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21802_ _02811_ _02849_ _02850_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25570_ _06290_ _06354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22782_ _02588_ _02616_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24521_ _05182_ _05305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21733_ _11409_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27240_ _01145_ clknet_leaf_82_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24452_ _05029_ _05236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21664_ _11138_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19668__B _11382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23403_ _04193_ _04230_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17967__I rbzero.map_rom.f2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20615_ _01702_ _01706_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_163_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27171_ _01076_ clknet_leaf_51_i_clk rbzero.wall_tracer.rayAddendX\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_191_i_clk_I clknet_5_9__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24383_ _05131_ _05122_ _05166_ _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21595_ _02642_ _02679_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__18342__A1 _07176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17145__A2 rbzero.pov.ss_buffer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26122_ _00032_ clknet_leaf_4_i_clk rbzero.spi_registers.spi_buffer\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23334_ _04167_ _04188_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_160_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20546_ _01637_ _01638_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26053_ _06772_ _06680_ _06824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23265_ _03898_ _04120_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20477_ _01568_ _01569_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25004_ _05393_ _05288_ _05255_ _05476_ _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_131_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_197_Right_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22216_ _11278_ _03096_ _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23196_ _03815_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_18_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22147_ _03120_ _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22992__A4 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14131__A2 _07920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22078_ _03074_ _03070_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26955_ _00865_ clknet_leaf_182_i_clk rbzero.tex_r1\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_128_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25906_ _06688_ _06624_ _06689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_156_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21029_ _12777_ _01579_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13920_ _07729_ _07730_ _07731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26886_ _00796_ clknet_5_10__leaf_i_clk rbzero.tex_r0\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_13851_ _07555_ _07661_ _07570_ _07662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25837_ _06606_ _06620_ _06621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19422__I _12169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16570_ _09998_ _10018_ _10021_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_48_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13782_ rbzero.tex_r0\[7\] _07592_ _07593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25768_ _06550_ _06542_ _06551_ _06552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_27_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__22901__A1 _12036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14985__A4 _07191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15521_ rbzero.spi_registers.texadd0\[17\] _09206_ _09211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24719_ _05258_ _05276_ _05233_ _05300_ _05503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_25699_ _06478_ _06482_ _06483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_195_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18240_ _11383_ _11384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_155_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15452_ rbzero.spi_registers.buf_vshift\[4\] _09154_ _09161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27438_ _01343_ clknet_leaf_72_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14403_ rbzero.tex_g0\[31\] _08210_ _08211_ _08212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_215_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15383_ rbzero.floor_leak\[5\] _09101_ _09109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18171_ _11112_ _11315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_232_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27369_ _01274_ clknet_leaf_98_i_clk rbzero.wall_tracer.trackDistY\[-11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17136__A2 _10485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17122_ _08106_ _10375_ _10497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15147__A1 _08926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14334_ rbzero.debug_overlay.vplaneX\[-9\] _08144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_170_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24406__A1 _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17053_ _10392_ _10443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15698__A2 _09340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14265_ rbzero.debug_overlay.facingX\[10\] _08075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_36_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16004_ _09547_ _09572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_94_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13216_ _07015_ _07030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_164_Right_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14196_ _07998_ _08005_ _08006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_210_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_210_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20443__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13147_ _06958_ _06953_ _06959_ _06960_ _06961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_148_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13078_ _06883_ _06888_ _06891_ _06893_ _06894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_17955_ _11098_ _11099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22196__A2 _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16906_ _07706_ _10301_ _10325_ _10326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16021__I _09550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17886_ _11000_ _11029_ _10998_ _11030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__21943__A2 _11392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19625_ _12206_ _12189_ _12396_ _12397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__24378__C _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16837_ _10236_ _10259_ _10265_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_220_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Left_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_19556_ _12327_ _12328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13633__A1 _07305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16768_ _10203_ _10204_ _10205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_221_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18507_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _11566_ _11567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15719_ _09357_ _09358_ _09348_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14476__I _07551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19487_ _12258_ _12259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16699_ _10092_ _10128_ _10142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13380__I gpout0.vpos\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18438_ rbzero.tex_g1\[36\] rbzero.tex_g1\[35\] _11523_ _11527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14189__A2 _07189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21459__A1 _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13936__A2 _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18369_ rbzero.tex_g1\[6\] rbzero.tex_g1\[5\] _11486_ _11488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20400_ _01425_ _01439_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21380_ _12465_ _01966_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14425__B _08220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20331_ _12283_ _12918_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25070__A1 _05838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_23050_ _03772_ _03842_ _03905_ _03906_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__19824__A1 _12595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20262_ _12955_ _13033_ _13034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_141_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24413__I _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22001_ _03019_ _03011_ _03021_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20193_ _12662_ _12223_ _12931_ _12965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_11_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_138_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23952_ _10491_ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26740_ _00650_ clknet_leaf_40_i_clk rbzero.pov.ready_buffer\[70\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input23_I i_reset vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22903_ rbzero.wall_tracer.trackDistX\[3\] _03605_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25125__A2 _05871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26671_ _00581_ clknet_leaf_34_i_clk rbzero.pov.ready_buffer\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_212_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23883_ rbzero.wall_tracer.rcp_fsm.o_data\[-2\] _04689_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_169_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15770__I _09037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25622_ _06404_ _06361_ _06405_ _06406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22834_ _12684_ _02112_ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_123_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23687__A2 rbzero.wall_tracer.stepDistY\[-10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25553_ _06302_ _06303_ _06337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21698__A1 _11307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22765_ _03621_ _03623_ _03624_ _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_177_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24504_ _05287_ _05271_ _05288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_137_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21716_ _02769_ _11114_ _02740_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25484_ _06178_ _06266_ _06267_ _06268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_192_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22696_ _03563_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27223_ _01128_ clknet_leaf_107_i_clk rbzero.wall_tracer.stepDistY\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24435_ _05218_ _05219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_137_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13927__A2 _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21647_ _02720_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_173_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20337__B _12311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27154_ _01059_ clknet_leaf_201_i_clk rbzero.map_rom.d6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24366_ _05063_ _05064_ _05148_ _05149_ _05150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_21578_ _02500_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26105_ _00015_ clknet_leaf_244_i_clk rbzero.spi_registers.spi_counter\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23317_ _03868_ _04050_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20529_ _01613_ _01621_ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27085_ _00995_ clknet_leaf_151_i_clk rbzero.tex_b1\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24297_ _05077_ _05078_ _05080_ _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__21947__I _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26036_ _10987_ _06810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14050_ rbzero.tex_r1\[10\] _07810_ _07859_ _07860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23248_ _04095_ _04103_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__24323__I _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23179_ _03922_ _03925_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17740_ _10920_ _10652_ _10923_ _10924_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_26938_ _00848_ clknet_leaf_185_i_clk rbzero.tex_r1\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14952_ _08754_ net4 _08755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__17054__A1 _08149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13903_ _07712_ _07713_ _07714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16776__I _10178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17671_ _10875_ rbzero.pov.ready_buffer\[13\] _10879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26869_ _00779_ clknet_leaf_166_i_clk rbzero.tex_r0\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14883_ _08685_ _08686_ _08687_ _08688_ _08334_ _08689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_19410_ _12181_ _12182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16622_ _10063_ _09977_ _10069_ _10036_ _10070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_199_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13834_ _07341_ _07645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_230_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13615__A1 _07325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_217_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19341_ _12133_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21689__A1 _11260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16553_ _10000_ _10003_ _10005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__14296__I _08105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13765_ _07575_ _07576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_210_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22350__A2 _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15504_ rbzero.spi_registers.texadd0\[13\] _09192_ _09198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19272_ rbzero.tex_b1\[17\] rbzero.tex_b1\[16\] _12094_ _12095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16484_ rbzero.wall_tracer.rayAddendY\[-4\] _09940_ _09941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13696_ _07479_ _07507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_210_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_233_Right_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18223_ _11362_ _11364_ _11366_ _11367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15435_ rbzero.spi_registers.buf_vshift\[0\] _09131_ _09148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13918__A2 rbzero.map_overlay.i_othery\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20247__B _12912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17400__I _06897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15366_ rbzero.spi_registers.buf_leak\[0\] _09092_ _09097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18154_ _11266_ _11277_ _11295_ _11297_ _11298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__18857__A2 _08751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17105_ _10483_ _10484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__20664__A2 _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14317_ rbzero.debug_overlay.vplaneX\[-6\] _08127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18085_ _11160_ _11161_ rbzero.wall_tracer.trackDistY\[-3\] _11175_ _11187_ _11229_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_15297_ _09044_ _09046_ _09042_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_151_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17036_ rbzero.pov.ready_buffer\[27\] _10412_ _10431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14248_ _07997_ _08038_ _08058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_123_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19806__A1 _12577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14179_ _06871_ _06886_ gpout0.hpos\[6\] _07988_ _07989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_110_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_245_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25355__A2 _06100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18987_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _11866_ _11867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13375__I _07185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17938_ _11081_ _11082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13308__C _07041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_53_Left_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__25107__A2 _05889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17869_ _11010_ _11011_ _11012_ _11013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15804__B _09417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19608_ _12379_ _12380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_233_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20880_ rbzero.wall_tracer.stepDistX\[7\] _12445_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19539_ _12310_ _12311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_159_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22550_ _11286_ _03449_ _03450_ rbzero.traced_texa\[-1\] _03453_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24618__A1 _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_200_Right_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21501_ _02478_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22481_ _03409_ _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_185_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17310__I _10602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Left_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24220_ _05002_ _05003_ _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_64_i_clk_I clknet_5_21__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21432_ _02495_ _02517_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_134_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14582__A2 _07821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16859__A1 rbzero.pov.ready_buffer\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24151_ _04781_ _04837_ _04935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__20655__A2 _12489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21363_ _02447_ _02448_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_142_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19665__C _12222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23102_ _03856_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__22372__B _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20314_ _01407_ _12995_ _01408_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24082_ _04757_ _04853_ _04866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_141_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21294_ _02379_ _02380_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_141_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17466__B _10751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23033_ _03890_ _03763_ _02767_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_229_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20245_ _12178_ _12011_ _12182_ _13016_ _13017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_247_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14602__C _07638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21080__A2 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20176_ _12663_ _12664_ _12935_ _12948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_71_Left_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24984_ _05558_ _05592_ _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_192_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26723_ _00633_ clknet_leaf_34_i_clk rbzero.pov.ready_buffer\[53\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23935_ _04737_ _04725_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__22580__A2 _09974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23866_ _02990_ _04690_ _04692_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_212_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26654_ _00564_ clknet_leaf_156_i_clk rbzero.tex_b0\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__20591__A1 _12398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25605_ _05977_ _06005_ _06389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_197_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22817_ _03646_ _03675_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_157_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23797_ _04627_ _04619_ _04633_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_175_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14270__A1 _08079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26585_ _00495_ clknet_leaf_34_i_clk rbzero.pov.spi_buffer\[54\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_200_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19700__I _12471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22332__A2 _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13550_ rbzero.row_render.size\[8\] _07357_ _07361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25536_ _06268_ _06313_ _06320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_22748_ rbzero.wall_tracer.trackDistX\[0\] _03599_ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_177_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25467_ _06028_ _06251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_192_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13481_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] _07292_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22679_ _02730_ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_212_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_212_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15220_ _08987_ _08988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17220__I _10543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27206_ _01111_ clknet_leaf_77_i_clk rbzero.wall_tracer.stepDistY\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24418_ _05042_ _05121_ _05130_ _05136_ _05038_ _05059_ _05202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_30_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25398_ _06041_ _06182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15151_ _07165_ _08931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_24349_ _05016_ _05133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_35_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18303__A4 _07149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27137_ _01047_ clknet_leaf_31_i_clk rbzero.wall_tracer.rayAddendX\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14102_ _07539_ _07912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15082_ gpout0.vpos\[7\] gpout0.vpos\[6\] _07216_ _08874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_27068_ _00978_ clknet_leaf_144_i_clk rbzero.tex_b1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_91_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26019_ _06745_ _06746_ _06794_ _05242_ _06795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__13533__B1 _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14033_ _07486_ _07843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18910_ rbzero.traced_texa\[9\] _07259_ _11821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_56_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19890_ _12661_ _12662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18841_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] _11765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_227_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18986__I _11850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13195__I _06992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18772_ _11717_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_209_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15984_ _09556_ _09557_ _09553_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__17027__A1 _08155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22020__A1 _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17723_ _10905_ _10913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14935_ _07770_ _08740_ _08192_ _08741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_240_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17654_ _10865_ _10567_ _10861_ _10867_ _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14866_ _08321_ _08670_ _08671_ _08672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_212_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16605_ _10050_ _10052_ _10054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_98_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13817_ _07340_ _07628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17585_ _10822_ _10823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14797_ rbzero.tex_b0\[5\] _08209_ _08604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22323__A2 _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19324_ rbzero.tex_b1\[40\] rbzero.tex_b1\[39\] _12120_ _12124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16536_ _09988_ _09989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13748_ rbzero.tex_r0\[40\] _07545_ _07539_ _07559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19255_ rbzero.tex_b1\[10\] rbzero.tex_b1\[9\] _12083_ _12085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16467_ _09923_ _09924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13679_ rbzero.tex_r0\[50\] _07487_ _07489_ _07490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_116_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18206_ _11349_ _11340_ _11306_ rbzero.map_rom.i_row\[4\] _11350_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_15418_ rbzero.spi_registers.buf_floor\[1\] _09119_ _09136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19186_ _12029_ _12030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16398_ rbzero.spi_registers.spi_buffer\[17\] _09865_ _09869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_207_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20637__A2 _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18137_ rbzero.wall_tracer.visualWallDist\[7\] _11281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15349_ _09083_ _09084_ _09073_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_247_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18068_ rbzero.wall_tracer.trackDistX\[-10\] _11212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_41_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15585__I _09258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17019_ _10407_ _10417_ _10418_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_10_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20030_ _12792_ _12793_ _12801_ _12802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_226_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17018__A1 rbzero.pov.ready_buffer\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21981_ rbzero.wall_tracer.size\[7\] _03005_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23720_ _02751_ _04565_ _03561_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20932_ _02015_ _02021_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_87_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23651_ _04358_ _04501_ _04502_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20863_ _01701_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22602_ _03483_ _03487_ _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_25_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26370_ _00280_ clknet_leaf_4_i_clk rbzero.spi_registers.buf_texadd1\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23582_ _04305_ _04433_ _04434_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_20794_ _01857_ _01884_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclkbuf_5_29__f_i_clk clknet_3_7_0_i_clk clknet_5_29__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_147_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25321_ _06063_ _06094_ _06105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_14_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22533_ _03442_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22078__A1 _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25252_ _06035_ _06036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_153_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22464_ _11462_ _07981_ _03401_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_161_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__23814__A2 _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24203_ _04986_ _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_228_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21415_ _12684_ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_118_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25183_ _05966_ _05967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22395_ _03327_ _03341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24134_ _04844_ _04915_ _04917_ _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_5_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21346_ _02402_ _02432_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__25567__A2 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24065_ rbzero.wall_tracer.rcp_fsm.operand\[9\] net75 _04847_ _04848_ _04849_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_131_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21277_ _02357_ _02363_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23016_ _03867_ _03873_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20228_ _12568_ _12999_ _12380_ _12520_ _13000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__22250__A1 rbzero.wall_tracer.visualWallDist\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20159_ _12398_ _12930_ _12931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17009__A1 _08073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19549__A3 _11068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24967_ _05650_ _05749_ _05638_ _05750_ _05751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_222_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14720_ rbzero.tex_b0\[41\] _08526_ _08308_ _08527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26706_ _00616_ clknet_leaf_61_i_clk rbzero.pov.ready_buffer\[36\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_231_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23918_ rbzero.wall_tracer.rcp_fsm.operand\[-10\] _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__23661__B _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18221__A3 _11306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24898_ _05678_ _05681_ _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_87_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14651_ _07337_ _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26637_ _00547_ clknet_leaf_148_i_clk rbzero.tex_b0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23849_ rbzero.wall_tracer.stepDistY\[10\] _04678_ _02760_ _04679_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_240_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13602_ _06857_ _07409_ _07412_ _07413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17370_ rbzero.pov.spi_buffer\[47\] _10674_ _10682_ _10683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_200_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15991__A1 _08980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14582_ rbzero.tex_g1\[18\] _07821_ _08389_ _08390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26568_ _00478_ clknet_leaf_64_i_clk rbzero.pov.spi_buffer\[37\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16321_ _09011_ _09804_ _09811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25519_ _05889_ _05999_ _06303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13533_ rbzero.floor_leak\[1\] _07343_ _07332_ rbzero.floor_leak\[2\] _07344_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26499_ _00409_ clknet_leaf_56_i_clk rbzero.debug_overlay.facingY\[-1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22069__A1 _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19040_ rbzero.tex_g0\[52\] rbzero.tex_g0\[51\] _11893_ _11897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_180_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16252_ _08926_ _09759_ _09760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13464_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] _07275_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__23805__A2 _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15203_ _08973_ _08969_ _08974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13395_ _07198_ _07202_ _07205_ _07206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_16183_ _09671_ _09707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_152_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_229_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15134_ rbzero.spi_registers.ss_buffer\[1\] _08867_ _08904_ _08916_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_129_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19942_ _12713_ _12304_ _12714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15065_ _08839_ _08824_ _08851_ _08858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_49_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14016_ _07825_ _07826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_242_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22241__A1 _12834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21044__A2 _13012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19873_ _12644_ _12645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__17799__A2 rbzero.pov.ready_buffer\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_18824_ _11738_ _11751_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_12_i_clk_I clknet_5_6__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_207_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18755_ _11707_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15967_ rbzero.spi_registers.spi_done _08842_ _09544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13653__I _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17706_ _10896_ _10621_ _10899_ _10901_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14918_ _08720_ _08721_ _08723_ _08564_ _08334_ _08724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_76_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18686_ _11668_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15898_ rbzero.spi_registers.buf_leak\[5\] _09481_ _09492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17637_ _10849_ _10551_ _10851_ _10855_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14849_ rbzero.tex_b1\[14\] _08277_ _08655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__20486__I _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17568_ _10813_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_237_i_clk_I clknet_5_6__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19173__A1 _11251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19307_ _12071_ _12114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16519_ _09972_ _09973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17499_ rbzero.tex_b0\[12\] rbzero.tex_b0\[11\] _10770_ _10774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19238_ _12075_ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_147_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13321__C _06905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19169_ _11949_ _12010_ _12011_ _12012_ _12013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA_clkbuf_5_20__f_i_clk_I clknet_3_5_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21200_ _02246_ _02287_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22180_ _03158_ _03115_ _03159_ _03160_ _09918_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__21283__A2 _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14433__B _07867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21131_ _02206_ _02218_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_113_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22083__I1 rbzero.wall_tracer.stepDistY\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21062_ _12300_ _01474_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_20013_ _12781_ _12783_ _12785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_25870_ _06645_ _06648_ _06653_ _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24821_ _05348_ _05605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_240_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21964_ rbzero.wall_tracer.rcp_fsm.o_data\[-6\] _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_24752_ _05523_ _05535_ _05536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__20546__A1 _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23703_ _04549_ _04550_ _12036_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20915_ _01999_ _02004_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_234_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24683_ _05334_ _05466_ _05467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21895_ _02920_ _08125_ _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24288__A2 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26422_ _00332_ clknet_leaf_251_i_clk rbzero.spi_registers.buf_texadd3\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23634_ _04478_ _04484_ _04485_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20846_ _12430_ _01608_ _01819_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14776__A2 _08554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23565_ _04222_ _04327_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26353_ _00263_ clknet_leaf_249_i_clk rbzero.spi_registers.buf_texadd0\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20777_ _01862_ _01867_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18911__A1 rbzero.traced_texa\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25304_ _06087_ _06088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_22516_ rbzero.wall_tracer.texu\[2\] _03429_ _03430_ _07450_ _03432_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14528__A2 _07894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26284_ _00194_ clknet_leaf_231_i_clk rbzero.spi_registers.buf_sky\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23496_ _04245_ _04006_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16823__B _10252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25235_ _06004_ _06017_ _06018_ _06019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_134_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22447_ _03385_ _03388_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__19467__A2 _12238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21274__A2 _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25166_ _05783_ _05948_ _05949_ _05236_ _05950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_13180_ rbzero.spi_registers.texadd0\[16\] _06913_ _06994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22471__A1 _08033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22116__I _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22378_ _12577_ _08041_ _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13738__I _07443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24117_ _04900_ _04901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21329_ _02405_ _02415_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25097_ _05880_ _05719_ _05844_ _05881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_36_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24212__A2 _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21955__I _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24048_ _04781_ _04830_ _04831_ _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_198_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22223__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14700__A2 _07938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_183_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19425__I _11381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16870_ rbzero.pov.ready_buffer\[46\] _10252_ _10294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20785__A1 _12501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_186_i_clk_I clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15821_ rbzero.spi_registers.buf_texadd3\[22\] _09118_ _09434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25999_ _06672_ _06777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_220_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18540_ rbzero.tex_r0\[16\] rbzero.tex_r0\[15\] _11581_ _11585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15752_ _09240_ _09383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_206_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14703_ _08504_ _08505_ _08508_ _08294_ _08509_ _08510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_18471_ rbzero.tex_g1\[50\] rbzero.tex_g1\[49\] _11544_ _11546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_231_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15683_ _09330_ _09331_ _09325_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_158_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17422_ rbzero.pov.spi_buffer\[60\] _10721_ _10718_ _10722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14634_ rbzero.tex_g1\[40\] _07810_ _08442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_184_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_202_i_clk clknet_5_13__leaf_i_clk clknet_leaf_202_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17353_ rbzero.pov.spi_buffer\[42\] _10670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14565_ _08373_ _08374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16304_ rbzero.spi_registers.buf_texadd2\[18\] _09791_ _09798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13516_ _07306_ _07308_ _07327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_222_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17284_ _10618_ _10619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14496_ rbzero.tex_g0\[40\] _07600_ _08305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19023_ _11871_ _11887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_141_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16235_ _09746_ _09747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13447_ _07257_ _07258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_8_i_clk clknet_5_1__leaf_i_clk clknet_leaf_8_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__18504__I _10757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19458__A2 _12229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_217_i_clk clknet_5_3__leaf_i_clk clknet_leaf_217_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_246_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__21265__A2 _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22462__A1 _11462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16166_ _08944_ _09687_ _09695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13378_ _07188_ _07189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15117_ rbzero.spi_registers.spi_counter\[6\] _08901_ _08902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16141__A1 _09591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16097_ rbzero.spi_registers.buf_texadd0\[15\] _09633_ _09642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21017__A2 _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22065__I1 _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19925_ _12696_ _12697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15048_ rbzero.spi_registers.spi_cmd\[2\] _08841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_19856_ _12548_ _12569_ _12496_ _12298_ _12628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_207_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18807_ _11737_ _11738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19787_ _12471_ _12411_ _12559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14479__I _07537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16999_ rbzero.pov.ready_buffer\[39\] _10403_ _10404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16995__A3 _10400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18738_ _11692_ _11698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__20528__A1 _12836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16908__B _09257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18669_ rbzero.tex_r1\[7\] rbzero.tex_r1\[6\] _11656_ _11659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17944__A2 rbzero.wall_tracer.rayAddendX\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20700_ _01789_ _01790_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21680_ _02739_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_164_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20631_ _01722_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_178_Right_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23350_ _04203_ _04204_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_46_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20562_ _01627_ _01654_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22301_ _03253_ _03260_ _03261_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_132_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23281_ _04076_ _04107_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20493_ _01508_ _01513_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_115_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25020_ _05549_ _05595_ _05804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22232_ _11248_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22163_ _03140_ _03147_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21114_ _02196_ _02201_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_112_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22094_ _03087_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26971_ _00881_ clknet_leaf_120_i_clk rbzero.texV\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_165_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25922_ _06688_ _06615_ _05880_ _06704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_21045_ _01996_ _01743_ _02002_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__20767__A1 _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25853_ _06590_ _06636_ _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_199_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24804_ _05388_ _05534_ _05588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25784_ _06559_ _06567_ _06568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22996_ _03850_ _03853_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24735_ _05518_ _05502_ _05519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_143_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21947_ _02982_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__21192__A1 _12299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27454_ _01359_ clknet_leaf_71_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_189_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24666_ _05441_ _05444_ _05449_ _05450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_16_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21878_ _02920_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__24130__A1 _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26405_ _00315_ clknet_leaf_245_i_clk rbzero.spi_registers.buf_texadd3\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20829_ _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23617_ _04412_ _04421_ _04468_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_27385_ _01290_ clknet_leaf_102_i_clk rbzero.wall_tracer.trackDistY\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19688__A2 _12447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24597_ _05373_ _05375_ _05380_ _05381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_154_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14350_ rbzero.debug_overlay.facingY\[-9\] _08160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_145_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_26336_ _00246_ clknet_leaf_238_i_clk rbzero.spi_registers.buf_texadd0\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21495__A2 _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23548_ _04313_ _04314_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_163_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13301_ rbzero.spi_registers.texadd2\[5\] _07108_ _07026_ rbzero.spi_registers.texadd0\[5\]
+ _07115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_14281_ _08080_ _08083_ _08086_ _08090_ _08091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_23479_ _04326_ _04332_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26267_ _00177_ clknet_leaf_15_i_clk rbzero.spi_registers.texadd3\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24433__A2 _05216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16020_ rbzero.spi_registers.buf_mapdxw\[0\] _09583_ _09584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13232_ _07045_ _07046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_25218_ _05996_ _06001_ _06002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__22444__A1 _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14921__A2 _08703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26198_ _00108_ clknet_leaf_12_i_clk rbzero.spi_registers.texadd0\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22995__A2 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13163_ _06940_ _06976_ _06977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25149_ _05287_ _05892_ _05933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__16123__A1 rbzero.spi_registers.buf_texadd0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13094_ rbzero.wall_hot\[0\] _06908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_17971_ rbzero.map_rom.f4 _11114_ _11115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_236_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19710_ _12481_ _12482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19155__I _11998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16922_ rbzero.pov.ready_buffer\[52\] _10169_ _10286_ _10339_ _10340_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_218_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19641_ _12412_ _12413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18671__I0 rbzero.tex_r1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16853_ _10272_ _10279_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_233_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25697__A1 _05949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14437__B2 _07463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25697__B2 _05951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15804_ _09419_ _09421_ _09417_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_232_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19572_ _12249_ _11079_ _12344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16784_ rbzero.pov.ready_buffer\[65\] _10201_ _10202_ _10218_ _10219_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_220_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13996_ rbzero.tex_r1\[30\] _07805_ _07806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_204_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_200_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23405__I _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18523_ _11575_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15735_ rbzero.spi_registers.texadd3\[0\] _09362_ _09370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_66_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25449__A1 _06037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_237_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17926__A2 _11069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_196_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18454_ rbzero.tex_g1\[43\] rbzero.tex_g1\[42\] _11533_ _11536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_141_i_clk clknet_5_14__leaf_i_clk clknet_leaf_141_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15666_ rbzero.spi_registers.texadd2\[6\] _09315_ _09319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19128__A1 _08162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17405_ _10696_ _10709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14617_ rbzero.tex_g1\[3\] _07878_ _08425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16019__I _09547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18385_ rbzero.tex_g1\[13\] rbzero.tex_g1\[12\] _11496_ _11497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__19679__A2 _12357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15597_ _09265_ _09266_ _09267_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17336_ rbzero.pov.spi_buffer\[38\] _10657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14548_ _07326_ _08357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_99_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15858__I _09139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_156_i_clk clknet_5_10__leaf_i_clk clknet_leaf_156_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17267_ _10571_ _10606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14479_ _07537_ _08288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19006_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _11877_ _11878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16218_ _09711_ _09734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13176__B2 _06926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14373__B1 _08047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14912__A2 _07592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17198_ rbzero.pov.spi_buffer\[3\] _10554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_178_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16149_ _09681_ _09682_ _09678_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_178_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15807__B _09417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22738__A2 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19908_ _12356_ _12358_ _12361_ _12222_ _12680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__19603__A2 _11071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18662__I0 rbzero.tex_r1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19839_ _12604_ _12609_ _12610_ _12611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_224_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22850_ _01945_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_247_Right_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_223_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21801_ _02845_ _02722_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22781_ _02642_ _02679_ _03639_ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_210_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_109_i_clk clknet_5_31__leaf_i_clk clknet_leaf_109_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_24520_ net90 _05304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21732_ _02768_ _02787_ _02788_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19119__A1 _08160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24451_ _05234_ _05235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_191_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21663_ _02728_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14873__S _08355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_134_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20614_ _01703_ _01705_ _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23402_ _04197_ _04229_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24382_ _04953_ _05122_ _05166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22674__A1 _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27170_ _01075_ clknet_leaf_51_i_clk rbzero.wall_tracer.rayAddendX\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_191_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21594_ _02644_ _02678_ _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17469__B _10751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23333_ _04170_ _04187_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_26121_ _00031_ clknet_leaf_5_i_clk rbzero.spi_registers.spi_buffer\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20685__B1 _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20545_ _01471_ _01630_ _01636_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_132_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18144__I rbzero.wall_tracer.visualWallDist\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13167__A1 _06927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26052_ _06816_ _06823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23264_ _04015_ _04119_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_131_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20476_ _01491_ _01542_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14903__A2 _08506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13288__I _07101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22215_ _03176_ _03189_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25003_ _05570_ _05785_ _05786_ _05787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23195_ _03860_ _04050_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20988__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__26560__CLK clknet_5_21__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22146_ _03119_ _03133_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__17853__A1 rbzero.debug_overlay.facingX\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16599__I _09988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22077_ rbzero.wall_tracer.stepDistY\[8\] _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_26954_ _00864_ clknet_leaf_182_i_clk rbzero.tex_r1\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25905_ _06630_ _06688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_145_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21028_ _02113_ _02116_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26885_ _00795_ clknet_leaf_165_i_clk rbzero.tex_r0\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA_clkbuf_leaf_59_i_clk_I clknet_5_23__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_242_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_199_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25836_ _06618_ _06601_ _06619_ _06620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13850_ _07655_ _07660_ _07661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_92_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_214_Right_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23154__A2 _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25767_ _06538_ _06539_ _06551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_230_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_48_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13781_ _07591_ _07592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22979_ _03724_ _03741_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_178_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15520_ _09207_ _09210_ _09202_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_219_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24718_ _05438_ _05450_ _05502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__15919__A1 _08962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25698_ _06480_ _06481_ _05979_ _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_195_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_27437_ _01342_ clknet_leaf_72_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15451_ rbzero.spi_registers.vshift\[4\] _09151_ _09160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24649_ _05346_ _05431_ _05432_ _05433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_i_clk clknet_5_29__leaf_i_clk clknet_leaf_73_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_61_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14402_ _07946_ _08211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_61_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22665__A1 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18170_ _11305_ _11311_ _11313_ _11314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27368_ _01273_ clknet_leaf_97_i_clk rbzero.wall_tracer.trackDistX\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15382_ _09107_ _09108_ _09100_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_232_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19530__A1 rbzero.wall_tracer.visualWallDist\[-11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17121_ _10495_ _10496_ _10492_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26319_ _00229_ clknet_leaf_214_i_clk rbzero.spi_registers.buf_mapdx\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14333_ _08142_ _08143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_135_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25603__A1 _05951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27299_ _01204_ clknet_leaf_209_i_clk rbzero.row_render.size\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14355__B1 _08046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17052_ _10427_ _10441_ _10442_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__22417__A1 rbzero.wall_tracer.texu\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14264_ _08071_ _08007_ _08023_ _08072_ _08017_ _08073_ _08074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_52_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_88_i_clk clknet_5_24__leaf_i_clk clknet_leaf_88_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16003_ _09570_ _09571_ _09565_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13215_ rbzero.spi_registers.texadd3\[22\] _07027_ _07028_ _07029_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_94_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23090__A1 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14195_ _08001_ _08004_ _08005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_210_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_210_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20443__A3 _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13146_ rbzero.spi_registers.texadd3\[7\] _06914_ _06923_ rbzero.spi_registers.texadd2\[7\]
+ _06909_ _06960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__21640__A2 _09971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14658__A1 _07841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23917__A1 _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13926__I rbzero.map_overlay.i_mapdx\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_11_i_clk clknet_5_4__leaf_i_clk clknet_leaf_11_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17954_ _11097_ _11098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13077_ _06892_ _06881_ _06893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__23393__A2 _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16905_ _10314_ _10321_ _10324_ _10325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17885_ _11002_ _11027_ _11028_ _11029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_245_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19624_ _12395_ _11388_ _12396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16836_ rbzero.pov.ready_buffer\[71\] _10260_ _10261_ _10263_ _10264_ _10265_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_178_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_i_clk clknet_5_20__leaf_i_clk clknet_leaf_26_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19555_ _08180_ _11097_ _12326_ _12159_ _12327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__14757__I _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16767_ rbzero.debug_overlay.playerX\[-5\] _10195_ _10204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13979_ _07760_ _06884_ _07778_ _07788_ _07789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_232_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18506_ _11565_ _11566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_220_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15718_ rbzero.spi_registers.buf_texadd2\[19\] _09353_ _09358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19486_ _12243_ _12245_ _12253_ _12257_ _12258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_75_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16698_ _10093_ _10128_ _10141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18437_ _11526_ _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15649_ rbzero.spi_registers.buf_texadd2\[1\] _09306_ _09307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__22656__A1 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18368_ _11487_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19521__A1 rbzero.wall_tracer.size\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14706__B _08280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18324__A2 _08753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17319_ _10643_ _10641_ _10644_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18299_ _11432_ _07228_ _11435_ _11437_ _11438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_79_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20330_ _12998_ _01424_ _13000_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_160_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14897__A1 _07609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20261_ _12977_ _13032_ _13033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19824__A2 _12199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22000_ rbzero.wall_tracer.size_full\[6\] _03020_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20192_ _12236_ _12963_ _12964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23908__A1 _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23951_ rbzero.wall_tracer.rcp_fsm.i_data\[-4\] _04740_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_60_i_clk_I clknet_5_23__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22902_ _03629_ _03631_ _03760_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26670_ _00580_ clknet_leaf_34_i_clk rbzero.pov.ready_buffer\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23882_ _03004_ _04699_ _04702_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input16_I i_mode[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25621_ _06359_ _06360_ _06405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22833_ _12691_ _02291_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_123_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21147__B2 _12192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25552_ _06332_ _06289_ _06335_ _06336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_79_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19679__B _12360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22764_ _03586_ _02688_ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_63_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_220_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24503_ net76 _05287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21715_ _02769_ _11114_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_25483_ _06170_ _06171_ _06135_ _06267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_22695_ _03562_ _11195_ _11400_ _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27222_ _01127_ clknet_leaf_113_i_clk rbzero.wall_tracer.stepDistY\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_43_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22647__A1 _12775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24434_ _05208_ _05213_ _05215_ _05217_ _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_47_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21646_ rbzero.wall_tracer.rayAddendY\[-7\] _01778_ _02719_ _02034_ _02720_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27153_ _01058_ clknet_leaf_225_i_clk reg_rgb\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24365_ _05065_ _05067_ _05069_ _04877_ _05149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_21577_ _02545_ _02551_ _02549_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_23_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26104_ _00014_ clknet_leaf_244_i_clk rbzero.spi_registers.spi_counter\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20528_ _12836_ _01620_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23316_ _04049_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24296_ _05079_ _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27084_ _00994_ clknet_leaf_151_i_clk rbzero.tex_b1\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_90_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24604__I _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18079__A1 _11200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26035_ _06769_ _06706_ _06742_ _06809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__23072__A1 _12733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23247_ _04097_ _04102_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20459_ _09901_ _01550_ _01552_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23178_ _03921_ _03925_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_246_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22129_ _09982_ _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_207_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_26937_ _00847_ clknet_leaf_185_i_clk rbzero.tex_r1\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14951_ net5 _08754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__22060__S _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17054__A2 _10443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13902_ rbzero.debug_overlay.playerY\[-1\] _07713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17670_ _10873_ _10582_ _10877_ _10878_ _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_26868_ _00778_ clknet_leaf_166_i_clk rbzero.tex_r0\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14882_ rbzero.tex_b1\[36\] _08288_ _08497_ _08688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__23127__A2 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16621_ _10064_ _10068_ _10069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_242_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25819_ _05951_ _05990_ _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13833_ rbzero.tex_r0\[29\] _07626_ _07644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21138__A1 _12684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26799_ _00709_ clknet_leaf_173_i_clk rbzero.tex_g1\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13615__A2 _07348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19340_ rbzero.tex_b1\[47\] rbzero.tex_b1\[46\] _12130_ _12133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16552_ _10000_ _10003_ _10004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_193_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13764_ _07482_ _07575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21689__A2 _12051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15503_ _09196_ _09197_ _09191_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19271_ _12093_ _12094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16565__A1 _10015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16483_ _09939_ _09940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15910__B _09491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13695_ _07497_ _07505_ _07506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_210_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18222_ _11345_ _11357_ _11365_ _11366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_15434_ rbzero.spi_registers.vshift\[0\] _09129_ _09147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_96_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14040__A2 _07843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18153_ _11296_ _11297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_15365_ rbzero.floor_leak\[0\] _09090_ _09096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17104_ _10482_ _10483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14316_ rbzero.debug_overlay.vplaneX\[0\] _08126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18084_ _11171_ _11182_ _11176_ _11228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15296_ rbzero.spi_registers.buf_othery\[2\] _09045_ _09046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19608__I _12379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17035_ _08162_ _10410_ _10430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14247_ rbzero.debug_overlay.playerY\[2\] _08057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19806__A2 _11068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14178_ _07208_ _07988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_245_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13129_ _06911_ _06941_ _06942_ _06943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18986_ _11850_ _11866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_175_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input8_I i_gpout1_sel[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17937_ _08082_ _11080_ _11081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16967__I _10377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_206_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17868_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] _11012_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_139_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25512__B1 _06148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19607_ _12374_ _12288_ _12377_ _12378_ _12379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16819_ _07694_ _10249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_191_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14264__C1 _08017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17799_ _10959_ rbzero.pov.ready_buffer\[57\] _10963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_220_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14803__A1 _07839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13606__A2 _07327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19538_ _12255_ _12310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_75_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19469_ _12213_ _12239_ _12241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21500_ _02583_ _02584_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22480_ _09972_ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__24094__A3 _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21431_ _02496_ _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_155_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16308__A1 _09000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24150_ _04933_ net66 _04934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21362_ _02314_ _02440_ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20313_ _12885_ _12481_ _12259_ _12988_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_23101_ _03912_ _03957_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__19518__I _12179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24081_ _04749_ _04864_ _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__14950__I _08752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21293_ _12683_ _01803_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23032_ _02761_ _03766_ _03889_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20244_ _12183_ _11039_ _13016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_219_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20175_ _12866_ _12945_ _12946_ _12947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__25346__A3 _06129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__26498__D _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14098__A2 _07906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24983_ _05763_ _05766_ _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13845__A2 _07591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26722_ _00632_ clknet_leaf_33_i_clk rbzero.pov.ready_buffer\[52\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_231_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23934_ rbzero.wall_tracer.rcp_fsm.operand\[-7\] _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_197_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20040__A1 _12667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26653_ _00563_ clknet_leaf_156_i_clk rbzero.tex_b0\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23865_ _03533_ _04687_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20591__A2 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25604_ _05983_ _06014_ _06388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22816_ _03666_ _03674_ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_197_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26584_ _00494_ clknet_leaf_34_i_clk rbzero.pov.spi_buffer\[53\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23796_ _03760_ _04632_ _04625_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19733__A1 _12468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14270__A2 _08011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25535_ _06264_ _06315_ _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__26019__C _05242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22747_ rbzero.wall_tracer.trackDistX\[0\] _03599_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__16547__A1 _08110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20343__A2 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25466_ _06203_ _06209_ _06249_ _06250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__22119__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13480_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] _07291_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22678_ _11409_ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_165_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_212_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21023__I _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27205_ _01110_ clknet_leaf_108_i_clk rbzero.wall_tracer.stepDistY\[-10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_212_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24417_ _05197_ _05198_ _05199_ _05200_ _05201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_205_Left_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16117__I _09599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21629_ rbzero.wall_tracer.rayAddendX\[-7\] _02689_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25397_ _06073_ _06181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_124_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14065__C _07604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15150_ _08928_ _08929_ _08930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27136_ _01046_ clknet_leaf_43_i_clk rbzero.wall_tracer.rayAddendX\[-8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24348_ _05121_ _05130_ _05131_ _04910_ _05038_ _05080_ _05132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_63_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14101_ rbzero.tex_r1\[42\] _07909_ _07910_ _07911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19428__I _12199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15081_ gpout0.vpos\[9\] _08786_ _08873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_27067_ _00977_ clknet_leaf_148_i_clk rbzero.tex_b1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24279_ _04977_ _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_91_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26018_ _06721_ _06704_ _06749_ _06794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14032_ _07586_ _07842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_121_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_227_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18840_ _11752_ _11764_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_227_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14089__A2 _07898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23348__A2 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18771_ rbzero.tex_r1\[51\] rbzero.tex_r1\[50\] _11714_ _11717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_214_Left_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15983_ _08973_ _09551_ _09557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_207_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19163__I _12006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17722_ _10903_ _10912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14934_ _07971_ _08738_ _08739_ _07242_ _08740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_240_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17653_ _10866_ rbzero.pov.ready_buffer\[7\] _10867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14865_ rbzero.tex_b1\[7\] _07633_ _08671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16604_ _10050_ _10052_ _10053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13816_ rbzero.tex_r0\[27\] _07626_ _07627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19024__I0 rbzero.tex_g0\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17584_ _10758_ _10822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14796_ _07337_ _08603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_85_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19323_ _12123_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_187_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16535_ _09916_ _09988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13747_ rbzero.tex_r0\[41\] _07537_ _07558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20334__A2 _12005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19254_ _12084_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_223_Left_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16466_ _09920_ _09923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13678_ _07488_ _07489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15210__A1 rbzero.spi_registers.spi_buffer\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14013__A2 _07822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18205_ _11302_ _11349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15417_ rbzero.color_floor\[1\] _09115_ _09135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23284__A1 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22087__A2 _12163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19185_ _11913_ _12009_ _12028_ _12029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_183_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16397_ rbzero.spi_registers.buf_texadd3\[17\] _09863_ _09868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_5_10__f_i_clk_I clknet_3_2_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18136_ _11278_ _11279_ _11280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_53_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15348_ rbzero.spi_registers.buf_mapdy\[5\] _09078_ _09084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24244__I _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_247_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18067_ rbzero.wall_tracer.trackDistX\[-10\] _11210_ _11211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15279_ _09029_ _09032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17018_ rbzero.pov.ready_buffer\[22\] _10403_ _10418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_238_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13386__I gpout0.vpos\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_233_i_clk_I clknet_5_3__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_232_Left_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18969_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _11856_ _11857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_225_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21980_ rbzero.wall_tracer.rcp_fsm.o_data\[-1\] _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_20931_ _02017_ _02020_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_179_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21770__A1 _08128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__22648__B _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20862_ _01951_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23650_ _04441_ _04444_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22601_ _07236_ _03472_ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_25_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_241_Left_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23581_ _04307_ _04432_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14945__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20793_ _01858_ _01883_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__17321__I _10611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25320_ _05977_ _06103_ _06104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_187_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22532_ rbzero.wall_tracer.visualWallDist\[-8\] _03436_ _03438_ rbzero.traced_texa\[-8\]
+ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25251_ _06034_ _06035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_170_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22463_ _07064_ _07187_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24202_ _04873_ _04979_ _04982_ _04985_ _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_21414_ _02001_ _02377_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25182_ _05910_ _05945_ _05965_ _05966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_135_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22394_ _03326_ _03339_ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24133_ _04916_ _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21345_ _02416_ _02431_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_32_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16701__A1 _10067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21276_ _02361_ _02362_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_24064_ _04844_ _04834_ _04845_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_103_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20227_ _12494_ _12999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23015_ _03869_ _03872_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_168_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20158_ _12929_ _12930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20089_ _12859_ _12860_ _12861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24966_ _05678_ _05681_ _05750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_222_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19954__A1 _12714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_222_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26705_ _00615_ clknet_leaf_61_i_clk rbzero.pov.ready_buffer\[35\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23917_ _04720_ _08814_ _04723_ _11473_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_99_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24897_ _05679_ _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__21761__A1 _10455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18221__A4 _11307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14650_ rbzero.tex_g1\[57\] _07906_ _08457_ _08458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26636_ _00546_ clknet_leaf_164_i_clk rbzero.tex_b0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_185_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23848_ rbzero.wall_tracer.trackDistY\[10\] _04677_ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19706__A1 _12476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15440__A1 rbzero.spi_registers.vshift\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23502__A2 _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13601_ rbzero.row_render.size\[9\] _07411_ _07412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_184_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14581_ rbzero.tex_g1\[19\] _07822_ _08389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_26567_ _00477_ clknet_leaf_63_i_clk rbzero.pov.spi_buffer\[36\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20316__A2 _12296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23779_ _03615_ _04617_ _04560_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16320_ rbzero.spi_registers.buf_texadd2\[22\] _09802_ _09810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25518_ _06301_ _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_184_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13532_ _07336_ _07343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_149_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26498_ _00408_ clknet_leaf_55_i_clk rbzero.debug_overlay.facingY\[-2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16251_ _09747_ _09759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25449_ _06037_ _06103_ _06233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23266__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_182_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13463_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] _07274_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_192_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21688__I _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15202_ rbzero.spi_registers.spi_buffer\[12\] _08973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16182_ _09705_ _09706_ _09700_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13394_ _07203_ _07204_ _07205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_63_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_229_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15133_ rbzero.spi_registers.spi_buffer\[2\] _08915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_27119_ _01029_ clknet_leaf_229_i_clk reg_vsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_211_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19941_ _12261_ _12713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15064_ rbzero.spi_registers.spi_counter\[2\] _08857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14015_ _07492_ _07825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_208_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_242_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19872_ rbzero.wall_tracer.stepDistX\[0\] _12643_ _12159_ _12644_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_242_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15259__A1 rbzero.map_overlay.i_otherx\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24518__A1 _05298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18823_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] _11750_ _11751_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__24369__I1 _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_207_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13809__A2 _07600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15966_ _09541_ _09543_ _09536_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18754_ rbzero.tex_r1\[44\] rbzero.tex_r1\[43\] _11703_ _11707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16310__I _09741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23741__A2 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17705_ _10897_ rbzero.pov.ready_buffer\[25\] _10901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14917_ rbzero.tex_b1\[59\] _08554_ _08722_ _08723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15897_ _09489_ _09490_ _09491_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18685_ rbzero.tex_r1\[14\] rbzero.tex_r1\[13\] _11666_ _11668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__20555__A2 _12448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_159_Right_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_69_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Left_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_172_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14848_ _07889_ _08635_ _08640_ _08645_ _08653_ _08654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_17636_ _10852_ rbzero.pov.ready_buffer\[2\] _10855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_102_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17567_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _10812_ _10813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14779_ _08582_ _08583_ _08585_ _08502_ _08565_ _08586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_59_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16518_ _09916_ _09971_ _09972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_19306_ _12113_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__19173__A2 _12015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17498_ _10773_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19237_ rbzero.tex_b1\[2\] rbzero.tex_b1\[1\] _12073_ _12075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16449_ _09904_ _09905_ _09906_ _09907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16931__A1 _10346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19168_ _11981_ _11983_ _11985_ _11997_ _12012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_26_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18119_ _11116_ _11263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_19099_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] _11943_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21130_ _02214_ _02217_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_197_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_113_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21061_ _01923_ _02149_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_245_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20012_ _12781_ _12783_ _12784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_225_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24820_ _05428_ _05429_ _05604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_226_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23762__B _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14473__A2 _07909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_129_Left_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__23732__A2 _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24751_ _05387_ _05525_ _05534_ _05535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_21963_ _02996_ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21743__A1 _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23702_ _11202_ _03041_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_234_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20914_ _02002_ _02003_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_96_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24682_ _05350_ _05354_ _05466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15422__A1 _08197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21894_ _02935_ _02931_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26421_ _00331_ clknet_leaf_252_i_clk rbzero.spi_registers.buf_texadd3\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23633_ _03861_ _04382_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20845_ _01822_ _01827_ _01934_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_232_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26352_ _00262_ clknet_leaf_249_i_clk rbzero.spi_registers.buf_texadd0\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23564_ _04220_ _04217_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20776_ _01865_ _01866_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_181_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25303_ _06085_ _06086_ _06087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_135_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22515_ _03431_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26283_ _00193_ clknet_leaf_227_i_clk rbzero.spi_registers.buf_sky\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23495_ _03491_ _04250_ _04348_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16922__A1 rbzero.pov.ready_buffer\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_138_Left_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25234_ _06008_ _06016_ _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23799__A2 _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22446_ _03386_ _03387_ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14624__B _07613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25165_ _05288_ _05949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22377_ _03322_ _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_161_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24116_ _04895_ _04867_ _04871_ _04899_ _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_21328_ _02408_ _02414_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25096_ _05520_ _05880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_53_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21259_ _02344_ _02345_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24047_ _04810_ _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_236_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_224_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20234__A1 _12986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_129_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21982__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_147_Left_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15820_ rbzero.spi_registers.texadd3\[22\] _09032_ _09433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25998_ _06720_ _06715_ _06775_ _06769_ _06776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_217_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15751_ rbzero.spi_registers.buf_texadd3\[4\] _09375_ _09382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24949_ _05730_ _05731_ _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_35_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_202_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14702_ _07496_ _08509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18470_ _11545_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15682_ rbzero.spi_registers.buf_texadd2\[10\] _09328_ _09331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17421_ _10696_ _10721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_185_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26619_ _00529_ clknet_leaf_163_i_clk rbzero.tex_b0\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14633_ _08435_ _08440_ _08441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17352_ _10668_ _10666_ _10669_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14564_ rbzero.trace_state\[2\] _08373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_56_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16303_ _09796_ _09797_ _09795_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_126_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_235_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13515_ _07325_ _07326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17283_ _10543_ _10618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14495_ _07479_ _08304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_246_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19022_ _11886_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16234_ _09458_ _09745_ _09746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_125_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13446_ gpout0.vpos\[8\] _07248_ _07250_ _07256_ _07257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_2_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16165_ rbzero.spi_registers.buf_texadd1\[7\] _09685_ _09694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17469__A2 _10544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13377_ gpout0.hpos\[2\] _07187_ _07188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15116_ rbzero.spi_registers.spi_counter\[5\] _08899_ _08901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16096_ _09640_ _09641_ _09637_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19924_ _12596_ _12696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15047_ _08839_ _08824_ _08840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_228_Right_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_239_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19855_ _12626_ _12382_ _12627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_247_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_235_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18806_ _08752_ _11737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16040__I _09599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19786_ _12422_ _12557_ _12558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16998_ _10396_ _10403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_222_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24397__C _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18737_ _11697_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15949_ _09530_ _09531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16975__I _08932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21725__A1 _11343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18668_ _11658_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_153_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17619_ net26 rbzero.tex_b0\[63\] _10838_ _10842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14495__I _07479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18599_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _11618_ _11619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14428__C _08222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20630_ _01715_ _01720_ _01721_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13332__C _06879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22150__A1 rbzero.wall_tracer.visualWallDist\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22150__B2 _11073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20561_ _01628_ _01653_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16904__A1 _10168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22300_ _11286_ _03237_ _03257_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13718__A1 _07507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13179__C1 _06918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20492_ _01503_ _01507_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23280_ _04079_ _04106_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22231_ _03201_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14391__A1 _08197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22162_ rbzero.wall_tracer.rcp_fsm.i_data\[-2\] _03144_ _03146_ _03147_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21113_ _02197_ _02200_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_160_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22093_ _03084_ _03086_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__18430__I _11479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26970_ _00880_ clknet_leaf_117_i_clk rbzero.texV\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_239_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25921_ _06702_ _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_165_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21044_ _12668_ _13012_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_165_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_130_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25852_ _06548_ _06635_ _06608_ _06636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_226_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24803_ _05584_ _05586_ _05587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25783_ _06560_ _06566_ _06567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__20519__A2 _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22995_ _03851_ _03852_ _03714_ _02260_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__19261__I _12072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24734_ net64 _05517_ _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_21946_ _02983_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_143_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18432__I1 rbzero.tex_g1\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27453_ _01358_ clknet_leaf_71_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24665_ _05445_ _05448_ _05449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_166_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21877_ _08122_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26404_ _00314_ clknet_leaf_244_i_clk rbzero.spi_registers.buf_texadd3\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23616_ _04415_ _04420_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_27384_ _01289_ clknet_leaf_104_i_clk rbzero.wall_tracer.trackDistY\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20828_ _01917_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24596_ _05376_ _05378_ _05379_ _05380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xclkbuf_5_13__f_i_clk clknet_3_3_0_i_clk clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26335_ _00245_ clknet_leaf_241_i_clk rbzero.spi_registers.buf_texadd0\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24269__I0 _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23547_ _04309_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20759_ _01848_ _01849_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13300_ rbzero.spi_registers.texadd3\[5\] _07111_ _07109_ rbzero.spi_registers.texadd1\[5\]
+ _07114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_55_i_clk_I clknet_5_25__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14280_ _08087_ _08064_ _08060_ _08088_ _08089_ _08090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_18_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26266_ _00176_ clknet_leaf_15_i_clk rbzero.spi_registers.texadd3\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23478_ _04328_ _04331_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25217_ _06000_ _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14382__A1 _07225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13231_ _07044_ _07045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22429_ _03321_ _07705_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26197_ _00107_ clknet_leaf_12_i_clk rbzero.spi_registers.texadd0\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25148_ _05931_ _05932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13162_ _06944_ _06974_ _06975_ _06976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14134__A1 _07507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25079_ _05827_ _05802_ _05862_ _05863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_13093_ rbzero.spi_registers.texadd0\[15\] _06907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_17970_ rbzero.map_rom.f3 _11099_ _11114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_155_Left_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14685__A2 _08491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19073__A1 _08159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16921_ _10238_ _10337_ _10338_ _10339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_217_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19640_ _12411_ _12412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_245_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16852_ _08175_ _10273_ _10278_ _10229_ _10279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_102_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15803_ rbzero.spi_registers.buf_texadd3\[17\] _09420_ _09421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19571_ _12342_ _12343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_137_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16783_ _10194_ _10217_ _10218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_189_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13995_ _07804_ _07805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_233_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15734_ _09368_ _09369_ _09361_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_66_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18522_ rbzero.tex_r0\[8\] rbzero.tex_r0\[7\] _11571_ _11575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_66_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22380__A1 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_237_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18453_ _11535_ _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15665_ _09316_ _09318_ _09314_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_158_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_164_Left_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_201_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17404_ rbzero.pov.spi_buffer\[55\] _10708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14616_ rbzero.tex_g1\[2\] _07876_ _08424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_233_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18384_ _11480_ _11496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15596_ _09241_ _09267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22132__A1 rbzero.wall_tracer.visualWallDist\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22132__B2 _11078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17335_ _10655_ _10653_ _10656_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14547_ _08333_ _08354_ _08355_ _08356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__18887__A1 rbzero.traced_texa\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20143__B1 _12910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22683__A2 _12499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17266_ rbzero.pov.spi_buffer\[20\] _10605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14478_ rbzero.tex_g0\[32\] _08258_ _08287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16217_ _09005_ _09732_ _09733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19005_ _11871_ _11877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13429_ _07238_ _07239_ _07240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13176__A2 _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14373__A1 _07708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17197_ _10551_ _10545_ _10553_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14373__B2 _08182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16148_ _08915_ _09676_ _09682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_173_Left_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_77_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24188__A2 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18250__I _11393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16079_ rbzero.spi_registers.buf_texadd0\[10\] _09622_ _09629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19907_ _12338_ _12340_ _12343_ _12369_ _12679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_19838_ _12543_ _12602_ _12610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 i_debug_map_overlay net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19769_ _12461_ _12505_ _12541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_160_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21800_ _09982_ _02844_ _02848_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_190_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22780_ _02585_ _02641_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22371__A1 _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_182_Left_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_125_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21731_ _11344_ _02782_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24450_ _05233_ _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21662_ _12044_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14600__A2 _07591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23401_ _04140_ _04233_ _04254_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_20613_ _12497_ _01607_ _01704_ _12492_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__22375__C _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24381_ _05082_ _05152_ _05164_ _05165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_129_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21593_ _02676_ _02677_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22674__A2 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26120_ _00030_ clknet_leaf_5_i_clk rbzero.spi_registers.spi_buffer\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20685__A1 rbzero.traced_texVinit\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21987__S _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23332_ _04171_ _04186_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_172_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20544_ _01471_ _01630_ _01636_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_144_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20685__B2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26051_ _06821_ _06822_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_172_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13167__A2 _06922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23263_ _04115_ _04118_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__23623__A1 _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20475_ _01493_ _01541_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_191_Left_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25002_ _05571_ _05573_ _05786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22214_ _03182_ _03183_ _03188_ _03180_ rbzero.wall_tracer.rcp_fsm.i_data\[8\] _03189_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_23194_ _03812_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_219_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14116__A1 _07555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22145_ rbzero.wall_tracer.rcp_fsm.i_data\[-5\] _03126_ _03132_ _03133_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17853__A2 rbzero.wall_tracer.rayAddendX\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14667__A2 _07919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22076_ _03022_ _03060_ _03073_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26953_ _00863_ clknet_leaf_183_i_clk rbzero.tex_r1\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
Xclkbuf_leaf_201_i_clk clknet_5_12__leaf_i_clk clknet_leaf_201_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25904_ _06606_ _06620_ _06687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_233_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21027_ _12816_ _01918_ _02115_ _12675_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_145_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26884_ _00794_ clknet_leaf_165_i_clk rbzero.tex_r0\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14419__A2 _08227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25835_ _06592_ _06600_ _06619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_7_i_clk clknet_5_4__leaf_i_clk clknet_leaf_7_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25766_ _06538_ _06539_ _06550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13780_ _07575_ _07591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_236_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_22978_ _03724_ _03741_ _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_216_i_clk clknet_5_6__leaf_i_clk clknet_leaf_216_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_48_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24717_ _05456_ _05500_ _05484_ _05501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_219_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_178_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21929_ _02951_ _02968_ _02959_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_219_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25697_ _05949_ _05975_ _06118_ _05951_ _06481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_178_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20912__A2 _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27436_ _01341_ clknet_leaf_72_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__25300__A1 _05869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15450_ _09158_ _09159_ _09149_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24648_ _05406_ _05430_ _05432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__22058__S _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22114__A1 _11081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16592__A2 _08105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14401_ _08209_ _08210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_61_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27367_ _01272_ clknet_leaf_95_i_clk rbzero.wall_tracer.trackDistX\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15381_ rbzero.spi_registers.buf_leak\[4\] _09103_ _09108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24579_ _05251_ _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__22665__A2 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17120_ rbzero.pov.ready_buffer\[2\] _10489_ _10496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19530__A2 _12301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26318_ _00228_ clknet_leaf_236_i_clk rbzero.spi_registers.buf_mapdx\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14332_ rbzero.debug_overlay.vplaneX\[-3\] _08142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_163_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27298_ _01203_ clknet_leaf_208_i_clk rbzero.row_render.size\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__25603__A2 _05998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14355__A1 _08159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17051_ rbzero.pov.ready_buffer\[31\] _10425_ _10442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14355__B2 _08160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14263_ rbzero.debug_overlay.facingX\[0\] _08073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26249_ _00159_ clknet_leaf_4_i_clk rbzero.spi_registers.texadd2\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__23614__A1 _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16002_ _09542_ _09562_ _09571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13214_ _07014_ _07028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_94_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14194_ _07976_ _08003_ _08004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23090__A2 _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_210_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13145_ rbzero.spi_registers.texadd1\[7\] _06915_ _06959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_210_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23917__A2 _08814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17953_ _11096_ _11097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13076_ _06858_ _06892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__21928__A1 _10478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16904_ _10168_ _10323_ _10324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17884_ rbzero.debug_overlay.facingX\[-2\] _11001_ _11028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_228_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_218_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_217_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24021__B _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19623_ rbzero.wall_tracer.stepDistX\[-11\] _12395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_189_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16835_ _10164_ _10264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19554_ _12320_ _12322_ _10184_ _12325_ _12326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_13978_ _07253_ _07779_ _07782_ _07787_ _07788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_87_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16766_ rbzero.debug_overlay.playerX\[-5\] _10195_ _10203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_232_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14291__B1 _08047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14830__A2 _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13633__A3 _07330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18505_ _11564_ _11565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15717_ rbzero.spi_registers.texadd2\[19\] _09350_ _09357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19485_ rbzero.wall_tracer.stepDistY\[-5\] _12256_ _11384_ _12257_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16697_ rbzero.wall_tracer.rayAddendY\[9\] _10140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_186_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18436_ rbzero.tex_g1\[35\] rbzero.tex_g1\[34\] _11523_ _11526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24247__I _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15648_ _09305_ _09306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14594__A1 _07842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15579_ _09251_ _09252_ _09253_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18367_ rbzero.tex_g1\[5\] rbzero.tex_g1\[4\] _11486_ _11487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17318_ rbzero.pov.spi_buffer\[34\] _10638_ _10635_ _10644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18298_ _07190_ _11433_ _11437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13389__I gpout0.vpos\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17249_ _10590_ _10583_ _10592_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20260_ _12979_ _13031_ _13032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18088__A2 _11227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25358__A1 _05996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20191_ _12334_ _12963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14649__A2 _07599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21919__A1 _10113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23950_ _04749_ _04743_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22901_ _12036_ _03755_ _03759_ _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_23881_ rbzero.wall_tracer.stepDistX\[-3\] _04694_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25620_ _06359_ _06360_ _06404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_212_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22832_ _02504_ _01918_ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21147__A2 _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25551_ _06333_ _06288_ _06334_ _06335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_140_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22763_ _03612_ _03622_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__19679__C _12352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24502_ _05257_ _05286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_177_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21714_ _02760_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_25482_ _06171_ _06135_ _06170_ _06266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_220_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22694_ _03556_ _03559_ _03561_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_228_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27221_ _01126_ clknet_leaf_113_i_clk rbzero.wall_tracer.stepDistY\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24433_ _05171_ _05216_ _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_240_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18155__I _11298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21645_ _09942_ rbzero.wall_tracer.rayAddendY\[-7\] _09907_ _02719_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__22647__A2 _12864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23996__I _08810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27152_ _01057_ clknet_leaf_182_i_clk reg_rgb\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_214_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24364_ _05041_ _05107_ _05108_ _05109_ _05148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_173_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21576_ _02660_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16326__A2 _09669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26103_ _00013_ clknet_leaf_244_i_clk rbzero.spi_registers.spi_counter\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14337__A1 _07205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23315_ _04057_ _04168_ _04169_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_20527_ _01619_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_27083_ _00993_ clknet_leaf_151_i_clk rbzero.tex_b1\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_127_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24295_ _04976_ net89 _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_162_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14888__A2 _07829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26034_ _06805_ _06807_ _05087_ _06808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_23246_ _04098_ _04101_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_133_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20458_ rbzero.traced_texVinit\[1\] _01551_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23177_ _04030_ _04032_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20389_ _12967_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_140_i_clk clknet_5_14__leaf_i_clk clknet_leaf_140_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_197_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22128_ _03113_ _03115_ _03116_ _03118_ _02887_ _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_219_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13312__A2 _07035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14950_ _08752_ _08753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_22059_ _03062_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26936_ _00846_ clknet_leaf_185_i_clk rbzero.tex_r1\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_227_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13901_ gpout0.vpos\[2\] _07712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__18251__A2 _11390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14881_ rbzero.tex_b1\[37\] _08631_ _08687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26867_ _00777_ clknet_leaf_166_i_clk rbzero.tex_r0\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
Xclkbuf_leaf_155_i_clk clknet_5_11__leaf_i_clk clknet_leaf_155_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_242_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16620_ _10067_ _10039_ _10053_ _10068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13832_ rbzero.tex_r0\[30\] _07641_ _07642_ _07643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25818_ _06593_ _06594_ _06599_ _06602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14273__B1 _08047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26798_ _00708_ clknet_leaf_131_i_clk rbzero.tex_g1\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_242_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21138__A2 _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14812__A2 _08614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16551_ _10001_ _10002_ _10003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25749_ _06491_ _06492_ _06533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_134_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13763_ _07507_ _07574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16014__A1 _08957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15502_ rbzero.spi_registers.buf_texadd0\[12\] _09194_ _09197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16482_ _09938_ _09939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19270_ _12071_ _12093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13694_ _07500_ _07502_ _07503_ _07504_ _07333_ _07505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_57_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15433_ _09140_ _09145_ _09146_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_18221_ _11120_ _11349_ _11306_ _11307_ _11365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_27419_ _01324_ clknet_leaf_84_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18152_ rbzero.wall_tracer.visualWallDist\[10\] _11296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15364_ _09094_ _09095_ _09089_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14315_ rbzero.debug_overlay.vplaneX\[-2\] _08125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17103_ _10481_ _10482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_230_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18083_ _11225_ _11226_ _11227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15295_ _08884_ _09045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__24016__B _08811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17034_ _10427_ _10428_ _10429_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14879__A2 _08250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14246_ rbzero.debug_overlay.playerY\[1\] _08053_ _08055_ _07681_ _08056_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17409__I _10546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14177_ _07211_ _07986_ _07987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_74_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_108_i_clk clknet_5_30__leaf_i_clk clknet_leaf_108_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_74_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_245_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13128_ rbzero.spi_registers.texadd0\[10\] _06911_ _06942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_239_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18985_ _11865_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_225_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__18227__C1 _07743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17936_ rbzero.wall_tracer.rayAddendX\[-1\] _11080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13059_ _06868_ _06876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__22574__A1 _11278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_177_i_clk_I clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22574__B2 rbzero.traced_texa\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17867_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] _11011_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__19290__I1 rbzero.tex_b1\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13672__I _07482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19606_ rbzero.wall_tracer.stepDistY\[-3\] _12310_ _12294_ _12378_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_178_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16818_ _10236_ _10244_ _10248_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14264__B1 _08023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22326__A1 _11284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17798_ _10958_ _10711_ _10961_ _10962_ _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_108_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14264__C2 _08073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19537_ _12308_ _12309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16749_ rbzero.debug_overlay.playerX\[-7\] _10188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_88_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19468_ _12213_ _12239_ _12240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_192_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18419_ rbzero.tex_g1\[28\] rbzero.tex_g1\[27\] _11512_ _11516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19399_ _07235_ _12170_ _12171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21430_ _02499_ _02515_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_146_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25579__A1 _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14008__I _07518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21361_ _02317_ _02439_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23100_ _03933_ _03956_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_140_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20312_ _12987_ _12259_ _12988_ _12481_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_24080_ _04746_ _04802_ _04863_ _04811_ _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_21292_ _12691_ _01805_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23031_ _02746_ _03887_ _03888_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_247_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20243_ _13013_ _13014_ _13015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__17808__A2 rbzero.pov.ready_buffer\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20174_ _12943_ _12944_ _12946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_229_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24554__A2 _05333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_72_i_clk clknet_5_29__leaf_i_clk clknet_leaf_72_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_196_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24982_ _05567_ _05575_ _05765_ _05766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_110_Left_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23933_ _04734_ _04735_ _04736_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26721_ _00631_ clknet_leaf_33_i_clk rbzero.pov.ready_buffer\[51\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16244__A1 _08915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26652_ _00562_ clknet_leaf_145_i_clk rbzero.tex_b0\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23864_ _02988_ _04690_ _04691_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_224_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25603_ _05951_ _05998_ _06387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_233_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22815_ _03667_ _03673_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26583_ _00493_ clknet_leaf_28_i_clk rbzero.pov.spi_buffer\[52\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23795_ _03612_ _04630_ _04631_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_196_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_175_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25534_ _06264_ _06315_ _06316_ _06317_ _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__19733__A2 _12485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22746_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] _03607_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_39_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16547__A2 rbzero.debug_overlay.vplaneY\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21540__A2 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25465_ _06029_ _06062_ _06249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13531__B _07341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22677_ _02789_ _03545_ _03546_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_10_i_clk clknet_5_4__leaf_i_clk clknet_leaf_10_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27204_ _01109_ clknet_leaf_108_i_clk rbzero.wall_tracer.stepDistY\[-11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_212_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24416_ _05186_ _05180_ _05163_ _05200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21628_ _10455_ rbzero.wall_tracer.rayAddendX\[-7\] _02705_ _02706_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_25396_ _06141_ _06179_ _06180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_191_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27135_ _01045_ clknet_leaf_31_i_clk rbzero.wall_tracer.rayAddendX\[-9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24347_ _04913_ _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21559_ _02536_ _02555_ _02643_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_106_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14100_ rbzero.tex_r1\[43\] _07625_ _07910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_62_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27066_ _00976_ clknet_leaf_151_i_clk rbzero.tex_b1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_15080_ _08869_ _08871_ _08872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_25_i_clk clknet_5_20__leaf_i_clk clknet_leaf_25_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_24278_ _04967_ _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_200_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_91_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26017_ _06792_ _06793_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14031_ _07468_ _07841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23229_ _03851_ _02079_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13533__A2 _07343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_227_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_227_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15972__I _09547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18770_ _11716_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_219_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15982_ rbzero.spi_registers.buf_mapdx\[2\] _09548_ _09556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22556__A1 _11292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17721_ _10904_ _10634_ _10908_ _10911_ _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14933_ _07767_ _08622_ _08623_ _07258_ _08739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_26919_ _00829_ clknet_leaf_130_i_clk rbzero.tex_r1\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_145_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_240_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17652_ _10844_ _10866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_215_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14864_ rbzero.tex_b1\[6\] _07617_ _08670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_202_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_225_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16603_ _10014_ _10033_ _10051_ _10009_ _10052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_13815_ _07625_ _07626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__19024__I1 rbzero.tex_g0\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14795_ _08595_ _08598_ _08601_ _08602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17583_ _10821_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_230_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19322_ rbzero.tex_b1\[39\] rbzero.tex_b1\[38\] _12120_ _12123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16534_ _09983_ _09986_ _09987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13746_ rbzero.tex_r0\[42\] _07545_ _07546_ _07557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_27_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17586__I1 rbzero.tex_b0\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14549__A1 _08201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__26610__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19253_ rbzero.tex_b1\[9\] rbzero.tex_b1\[8\] _12083_ _12084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16465_ _09901_ _09913_ _09922_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13677_ _07335_ _07488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15210__A2 _08975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18204_ _11338_ _11111_ _11120_ _11107_ _11348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_183_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15416_ _09133_ _09134_ _09112_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16396_ _09864_ _09866_ _09867_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19184_ _11307_ _12016_ _12027_ _12028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18135_ rbzero.wall_tracer.visualWallDist\[8\] _11279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15347_ rbzero.map_overlay.i_mapdy\[5\] _09075_ _09083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_207_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18160__A1 _11301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_247_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18066_ _11209_ _11210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15278_ _09030_ _09031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__24461__S _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21047__A1 _12210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13667__I _07348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_17017_ _08160_ _10401_ _10417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13524__A2 _07334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14229_ _08038_ _08034_ _08039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__16043__I _09564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24260__I _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_237_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18968_ _11850_ _11856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17919_ _11042_ _11061_ _11062_ _11063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_206_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18899_ _11769_ _11812_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_240_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20930_ _02018_ _02019_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_221_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20861_ _01949_ _01950_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19015__I1 rbzero.tex_g0\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22600_ _03080_ _03482_ _03485_ _03199_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_178_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23580_ _04307_ _04432_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20792_ _01869_ _01882_ _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_187_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22531_ _03441_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_146_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13351__B net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16218__I _09711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25250_ _05580_ _06034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_147_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22462_ _11462_ _07187_ _03400_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__24435__I _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_170_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24201_ _04918_ _04983_ _04984_ _04963_ _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_134_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21413_ _02497_ _02498_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_25181_ _05946_ _05961_ _05964_ _05965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_161_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22393_ _01550_ _03329_ _03338_ _03339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_135_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24132_ _04842_ _04883_ _04916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_60_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21344_ _02419_ _02430_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24063_ _04796_ rbzero.wall_tracer.rcp_fsm.operand\[9\] _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_21275_ _12692_ _02212_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_130_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25266__I _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23014_ _03870_ _03871_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_38_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20226_ _12486_ _12586_ _12998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14910__B _08603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16465__A1 _09901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20157_ rbzero.wall_tracer.visualWallDist\[1\] _12200_ _12929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13279__A1 _07053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22538__A1 rbzero.wall_tracer.visualWallDist\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24965_ _05678_ _05681_ _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20088_ _12858_ _12806_ _12830_ _12857_ _12860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_231_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_222_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26704_ _00614_ clknet_leaf_61_i_clk rbzero.pov.ready_buffer\[34\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_222_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23916_ rbzero.wall_tracer.rcp_fsm.i_data\[-11\] _04722_ _04723_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14201__I _08010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24896_ _05678_ _05679_ _05680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23847_ _04674_ _04675_ _04676_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26635_ _00545_ clknet_leaf_161_i_clk rbzero.tex_b0\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14779__B2 _08502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15440__A2 _09151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13600_ rbzero.row_render.size\[8\] _07389_ _07411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_212_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14580_ rbzero.tex_g1\[17\] _07818_ _07646_ _08388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23778_ _04530_ _04615_ _04616_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_138_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26566_ _00476_ clknet_leaf_63_i_clk rbzero.pov.spi_buffer\[35\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_200_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13531_ rbzero.floor_leak\[1\] _07337_ _07341_ rbzero.floor_leak\[0\] _07342_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_39_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25517_ _06299_ _06300_ _06301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22729_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] _03584_
+ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13261__B _07074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26497_ _00407_ clknet_leaf_56_i_clk rbzero.debug_overlay.facingY\[-3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25255__A3 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16250_ rbzero.spi_registers.buf_texadd2\[4\] _09757_ _09758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_125_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25448_ _06229_ _06231_ _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13462_ rbzero.texV\[6\] _07273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__24463__A1 _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15201_ rbzero.spi_registers.spi_buffer\[13\] _08960_ _08972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19439__I _12210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_209_Right_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13754__A2 _07543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16181_ _08968_ _09698_ _09706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25379_ _06115_ _06116_ _06163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13393_ gpout0.vpos\[4\] _07204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15132_ _08912_ _08907_ _08914_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_229_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27118_ _01028_ clknet_leaf_225_i_clk reg_hsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24215__A1 _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21029__A1 _12777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19940_ _12707_ _12710_ _12711_ _12712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_15063_ _08837_ _08838_ _08850_ _08855_ _08856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_27049_ _00959_ clknet_leaf_203_i_clk rbzero.wall_tracer.mapY\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__14703__B2 _08294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14014_ rbzero.tex_r1\[26\] _07821_ _07823_ _07824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19871_ rbzero.wall_tracer.stepDistY\[0\] _12642_ _12167_ _12643_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_242_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_242_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15259__A2 _08879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18822_ _11746_ _11748_ _11749_ _11750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__24518__A2 _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_207_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18753_ _11706_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15965_ _09542_ _09527_ _09543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_234_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19902__I _12427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17704_ _10896_ _10617_ _10899_ _10900_ _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_136_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14916_ rbzero.tex_b1\[58\] _08226_ _08722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_18684_ _11667_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15896_ _09429_ _09491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17635_ _10849_ _10549_ _10851_ _10854_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14847_ _08315_ _08652_ _08653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_199_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15431__A2 _08879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17566_ _10801_ _10812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_187_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14778_ rbzero.tex_b0\[12\] _08499_ _08584_ _08585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22701__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19305_ rbzero.tex_b1\[32\] rbzero.tex_b1\[31\] _12109_ _12113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16517_ _07240_ _08869_ _09971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_191_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13729_ rbzero.tex_r0\[32\] _07535_ _07539_ _07540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17497_ rbzero.tex_b0\[11\] rbzero.tex_b0\[10\] _10770_ _10773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_82_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19236_ _12074_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16448_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] _09906_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19167_ _12002_ _11951_ _12011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__13745__A2 _07543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16379_ _08932_ _09855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_182_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18118_ rbzero.debug_overlay.playerX\[4\] _11259_ _11260_ _07681_ _11261_ _11262_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_53_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19098_ _11920_ _11940_ _11941_ _11942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18049_ rbzero.wall_tracer.trackDistY\[-5\] _11193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22768__A1 _11163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21060_ _01922_ _01927_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_113_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19633__A1 rbzero.debug_overlay.playerY\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22503__I _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16447__A1 rbzero.debug_overlay.vplaneY\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20011_ _12705_ _12782_ _12783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16501__I rbzero.wall_tracer.rayAddendY\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24750_ _05527_ _05528_ _05529_ _05533_ _05534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_21962_ rbzero.wall_tracer.rcp_fsm.o_data\[-7\] rbzero.wall_tracer.size\[1\] _02983_
+ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_222_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23701_ _04543_ _04547_ _04548_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_20913_ _12661_ _01743_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24681_ _04919_ _05464_ _05465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21893_ _02927_ _02928_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26420_ _00330_ clknet_leaf_252_i_clk rbzero.spi_registers.buf_texadd3\[16\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23632_ _04479_ _04480_ _04483_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20844_ _01816_ _01821_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26351_ _00261_ clknet_leaf_2_i_clk rbzero.spi_registers.buf_texadd0\[19\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23563_ _04321_ _01972_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20775_ _12209_ _01743_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25302_ _05971_ _06086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22514_ rbzero.wall_tracer.texu\[1\] _03429_ _03430_ rbzero.row_render.texu\[1\]
+ _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_130_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26282_ _00192_ clknet_leaf_230_i_clk rbzero.spi_registers.buf_sky\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23494_ _03898_ _04347_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15787__I _09117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25233_ _06008_ _06016_ _06017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22445_ _03374_ _03377_ _03387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25164_ _05639_ _05948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_162_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22376_ _11394_ _12173_ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_60_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24115_ _04896_ _04898_ _04899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21327_ _02410_ _02413_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25095_ _05331_ _05725_ _05879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22759__A1 _11165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24046_ _04829_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_198_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19624__A1 _12395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21258_ _02068_ _01437_ _01604_ _02066_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_53_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_224_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20209_ _12903_ _12921_ _12981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21189_ _12383_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_244_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_148_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17951__B _11094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_51_i_clk_I clknet_5_23__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25997_ _06701_ _06705_ _06707_ _06775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__23184__A1 _12428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15750_ rbzero.spi_registers.texadd3\[4\] _09373_ _09381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24948_ _05730_ _05731_ _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_14701_ rbzero.tex_b0\[50\] _08506_ _08507_ _08508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_202_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15681_ rbzero.spi_registers.texadd2\[10\] _09326_ _09330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24879_ _05661_ _05662_ _05663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_213_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17420_ rbzero.pov.spi_buffer\[59\] _10720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_200_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26618_ _00528_ clknet_leaf_163_i_clk rbzero.tex_b0\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14632_ _08436_ _08437_ _08438_ _08439_ _07638_ _08440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_157_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14563_ _08371_ _07697_ _07242_ _08372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17351_ rbzero.pov.spi_buffer\[42\] _10662_ _10659_ _10669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26549_ _00459_ clknet_leaf_25_i_clk rbzero.pov.spi_buffer\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16302_ _08994_ _09793_ _09797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15177__A1 _08950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13514_ _07323_ _07324_ _07325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_235_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17282_ rbzero.pov.spi_buffer\[24\] _10617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14494_ _08297_ _08299_ _08302_ _08255_ _08262_ _08303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_43_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19021_ rbzero.tex_g0\[44\] rbzero.tex_g0\[43\] _11882_ _11886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13727__A2 _07537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16233_ _08821_ _08833_ _09745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13445_ _07253_ _07255_ _07207_ _07256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__14924__B2 _08360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16164_ _09692_ _09693_ _09689_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13376_ _07056_ _06904_ _07187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_50_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15115_ _08894_ _08900_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16095_ _08980_ _09635_ _09641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_192_Right_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19923_ _12689_ _12691_ _12693_ _12694_ _12695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_15046_ rbzero.spi_registers.spi_cmd\[3\] _08839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_121_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19615__A1 _12260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__21422__A1 _12788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19854_ _12486_ _12626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_236_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18805_ _11736_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19785_ _12500_ _12557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16997_ _08072_ _10401_ _10402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15652__A2 _09306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18736_ rbzero.tex_r1\[36\] rbzero.tex_r1\[35\] _11693_ _11697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15948_ _08822_ _08845_ _09530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18667_ rbzero.tex_r1\[6\] rbzero.tex_r1\[5\] _11656_ _11658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15879_ _08908_ _09478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17618_ _10841_ _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22993__I _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24675__A1 _05328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18598_ _11607_ _11618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_164_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13966__A2 _07750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17549_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _10802_ _10803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18354__A1 _07041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15168__A1 _08944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20560_ _01640_ _01652_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_15_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24427__A1 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16904__A2 _10323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13179__B1 _06992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19219_ _12054_ _12049_ _12050_ _12060_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_117_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14915__A1 rbzero.tex_b1\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20491_ _01515_ _01538_ _01583_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_15_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22989__B2 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22230_ _03200_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22161_ _11986_ _03134_ _03145_ _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21112_ _02198_ _02199_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14143__A2 _07583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22092_ _11393_ _03085_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_140_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_246_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25920_ _05089_ _06702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_165_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21043_ _01915_ _01929_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__16231__I _09742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25544__I _06271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25851_ _06571_ _06635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_199_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5_0_i_clk clknet_0_i_clk clknet_3_5_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_226_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24802_ _05533_ _05585_ _05586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_25782_ _06561_ _06565_ _06566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22994_ _01437_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_179_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21945_ _02982_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24733_ _05509_ _05511_ _05516_ _05517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_241_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18158__I _11252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27452_ _01357_ clknet_leaf_72_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24664_ _05446_ _05447_ _05448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_139_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21876_ _02908_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_194_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23615_ _04465_ _04466_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26403_ _00313_ clknet_leaf_248_i_clk rbzero.spi_registers.buf_texadd2\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24130__A3 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20827_ _01916_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_27383_ _01288_ clknet_leaf_103_i_clk rbzero.wall_tracer.trackDistY\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24595_ _05305_ _05264_ _05353_ _05379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_148_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26334_ _00244_ clknet_leaf_242_i_clk rbzero.spi_registers.buf_texadd0\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23546_ _04283_ _04299_ _04398_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_20758_ _01832_ _01847_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24269__I1 _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26265_ _00175_ clknet_leaf_15_i_clk rbzero.spi_registers.texadd3\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23477_ _04329_ _04330_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16406__I _09814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20689_ _01773_ _01774_ _01772_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25216_ _05999_ _06000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13230_ gpout0.hpos\[1\] _07044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22428_ _03370_ _03371_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14382__A2 _07230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26196_ _00106_ clknet_leaf_12_i_clk rbzero.spi_registers.texadd0\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__23641__A2 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16659__A1 _09953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25147_ _05929_ _05930_ _05931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13161_ rbzero.texu_hot\[5\] _06939_ _06975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22359_ _11330_ _11359_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15331__A1 rbzero.map_overlay.i_mapdy\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25394__A2 _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25078_ _05828_ _05860_ _05861_ _05862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_13092_ _06905_ _06906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_130_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24029_ _04733_ rbzero.wall_tracer.rcp_fsm.operand\[-9\] rbzero.wall_tracer.rcp_fsm.operand\[-10\]
+ rbzero.wall_tracer.rcp_fsm.operand\[-11\] _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_16920_ rbzero.debug_overlay.playerY\[-1\] _10335_ _10338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23683__B _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16851_ _10277_ _10278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__19452__I _12223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24354__B1 _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15802_ _09117_ _09420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_176_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19570_ _08172_ _11097_ _12341_ _12158_ _12342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_16782_ rbzero.debug_overlay.playerX\[-3\] _10216_ _10217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_13994_ _07534_ _07804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_88_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22904__A1 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18521_ _11574_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15733_ rbzero.spi_registers.buf_texadd2\[23\] _09364_ _09369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13714__B _07524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18452_ rbzero.tex_g1\[42\] rbzero.tex_g1\[41\] _11533_ _11535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_237_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15664_ rbzero.spi_registers.buf_texadd2\[5\] _09317_ _09318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_200_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17403_ _10704_ _10700_ _10707_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14615_ _07848_ _08421_ _08422_ _08423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13948__A2 _07757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18383_ _11495_ _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_185_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17139__A2 _10507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15595_ rbzero.spi_registers.buf_texadd1\[12\] _09259_ _09266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14070__A1 _07842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17334_ rbzero.pov.spi_buffer\[38\] _10650_ _10646_ _10656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__24409__A1 _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20143__A1 rbzero.wall_tracer.stepDistY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14546_ _07349_ _08355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18887__A2 rbzero.texV\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23880__A2 _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21891__A1 _11069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17265_ _10601_ _10594_ _10604_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14477_ _08278_ _08281_ _08283_ _08284_ _08285_ _08286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__15220__I _08987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19004_ _11876_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16216_ _09674_ _09732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13428_ rbzero.trace_state\[1\] rbzero.trace_state\[0\] _07239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__14373__A2 _08007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17196_ rbzero.pov.spi_buffer\[3\] _10547_ _10552_ _10553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16147_ rbzero.spi_registers.buf_texadd1\[2\] _09672_ _09681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13359_ net24 _07171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_178_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23149__I _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16078_ _09627_ _09628_ _09626_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_110_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13675__I _07418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19906_ _12315_ _12318_ _12328_ _12352_ _12678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_15029_ _08821_ _08822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_227_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22988__I _12212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13884__A1 _07694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19837_ _12543_ _12602_ _12609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_224_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23148__A1 _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19768_ _12508_ _12538_ _12540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput2 i_debug_trace_overlay net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_190_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23699__A2 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18719_ _11671_ _11687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_19699_ _12470_ _12471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_108_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22371__A2 _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21730_ _10258_ _02784_ _02786_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_125_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24648__A1 _05406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21661_ _02727_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23400_ _04143_ _04232_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__22123__A2 _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20612_ _13024_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24380_ _05099_ _05157_ _05162_ _05163_ _05164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_145_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21592_ _02646_ _02675_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16889__A1 rbzero.pov.ready_buffer\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23331_ _04176_ _04178_ _04185_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20543_ _01634_ _01635_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_149_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21882__A1 _10477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26050_ _06758_ rbzero.wall_tracer.rcp_fsm.o_data\[1\] _06759_ _06822_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23262_ _03900_ _04116_ _04117_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14364__A2 _08064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20474_ _01562_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_41_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25001_ _05571_ _05573_ _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22213_ _03177_ _03187_ _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23193_ _02621_ _03929_ _04048_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_42_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14902__C _07839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22144_ _11990_ _03121_ _03125_ _03131_ _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15313__A1 _09056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_224_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22075_ _03072_ _03070_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26952_ _00862_ clknet_leaf_183_i_clk rbzero.tex_r1\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_195_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25903_ _06643_ _06686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21026_ _02114_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_145_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26883_ _00793_ clknet_leaf_164_i_clk rbzero.tex_r0\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_145_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25834_ _06547_ _06616_ _06617_ _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__13627__A1 _07433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25765_ _06518_ _06543_ _06549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22977_ _03833_ _03834_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24716_ _05389_ _05391_ _05405_ _05500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_219_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20373__A1 _12403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21928_ _10478_ _10474_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_25696_ _06479_ _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_178_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_219_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27435_ _01340_ clknet_leaf_78_i_clk rbzero.wall_tracer.rcp_done vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24103__A3 _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24647_ _05430_ _05406_ _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__18616__I _11564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21859_ _02715_ _02899_ _02903_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18318__A1 _07712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14052__B2 _07861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14400_ _07498_ _08209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27366_ _01271_ clknet_leaf_100_i_clk rbzero.wall_tracer.trackDistX\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15380_ rbzero.floor_leak\[4\] _09101_ _09107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24578_ _05361_ _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26317_ _00227_ clknet_leaf_214_i_clk rbzero.spi_registers.buf_mapdx\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14331_ _08138_ _08006_ _08036_ _08140_ _08141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__16136__I _09671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23529_ _04059_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27297_ _01202_ clknet_leaf_208_i_clk rbzero.row_render.size\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17050_ _08159_ _10423_ _10441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14262_ rbzero.debug_overlay.facingX\[-3\] _08072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14355__A2 _08016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26248_ _00158_ clknet_leaf_18_i_clk rbzero.spi_registers.texadd2\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13213_ _06927_ _07027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16001_ rbzero.spi_registers.buf_mapdy\[1\] _09560_ _09570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15975__I _09550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20428__A2 _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14193_ _08002_ _08003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_94_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26179_ _00089_ clknet_leaf_223_i_clk rbzero.spi_registers.vshift\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_94_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13144_ rbzero.spi_registers.texadd0\[7\] _06958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__14812__C _08198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_210_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_210_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17952_ _11095_ _11096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13075_ _06890_ _06869_ _06891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__21928__A2 _10474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16903_ rbzero.debug_overlay.playerY\[-3\] _10322_ _10323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_17883_ _11003_ _11024_ _11026_ _11027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_19622_ _12309_ _12373_ _12389_ _12394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_16834_ _10171_ _10262_ _10263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13618__A1 gpout0.vinf vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_221_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19553_ _12324_ _12325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_232_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16765_ _10178_ _10202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_221_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14291__A1 _08099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13977_ _07783_ _07784_ _07785_ _07786_ _07787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_88_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15215__I rbzero.spi_registers.spi_buffer\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18504_ _10757_ _11564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_17_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15716_ _09355_ _09356_ _09348_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19484_ _12255_ _12256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16696_ _09998_ _10138_ _10139_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18435_ _11525_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15647_ _09257_ _09305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_185_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14043__A1 _07841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23302__A1 _12428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18366_ _11480_ _11486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_127_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15578_ _09241_ _09253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17317_ rbzero.pov.spi_buffer\[33\] _10643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14529_ _08335_ _08336_ _08337_ _08338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_173_i_clk_I clknet_5_9__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25055__A1 _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18297_ _07190_ _11433_ _11435_ _11436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_83_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17248_ rbzero.pov.spi_buffer\[16\] _10591_ _10588_ _10592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19809__A1 _12171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17179_ rbzero.pov.ss_buffer\[1\] _10515_ _10539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_101_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20190_ _12841_ _12961_ _12962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13306__B1 _07109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22900_ _03756_ _03757_ _03758_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_224_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23880_ _12287_ _04686_ _04701_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__24869__A1 _05328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_98_i_clk_I clknet_5_27__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22831_ _02634_ _02635_ _03689_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14282__A1 _08076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15125__I _08908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25550_ _06036_ _06088_ _06282_ _06284_ _06334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_22762_ _03619_ _03620_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_177_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23342__I _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24501_ _05241_ _05266_ _05285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21713_ _02768_ _02771_ _02772_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25481_ _06174_ _06177_ _06265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_78_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22693_ _03560_ _01661_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17771__A2 rbzero.pov.ready_buffer\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27220_ _01125_ clknet_leaf_109_i_clk rbzero.wall_tracer.stepDistY\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24432_ _05102_ _05113_ _05057_ _05216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_21644_ _02708_ _02717_ _02718_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14585__A2 _07872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24374__S _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23844__A2 _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_214_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24363_ _04898_ _05035_ _05052_ _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_173_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20658__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27151_ _01056_ clknet_leaf_225_i_clk reg_rgb\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21575_ _02544_ _02657_ _02659_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23314_ _04061_ _04069_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26102_ _00012_ clknet_leaf_244_i_clk rbzero.spi_registers.spi_counter\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20526_ rbzero.wall_tracer.stepDistX\[5\] _01524_ _01618_ _01619_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_138_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15534__A1 rbzero.spi_registers.buf_texadd0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27082_ _00992_ clknet_leaf_150_i_clk rbzero.tex_b1\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14337__A2 _08120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24294_ _04946_ _04942_ _05046_ _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_26033_ _06662_ _06739_ _06806_ _06807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_23245_ _04099_ _04100_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__18171__I _11112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20457_ _10019_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_41_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14632__C _07638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25349__A2 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23176_ _03928_ _04031_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20388_ _12971_ _12779_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_242_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22127_ _11993_ _03095_ _03117_ _11079_ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_246_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17039__A1 _08153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22058_ rbzero.wall_tracer.rcp_fsm.o_data\[1\] rbzero.wall_tracer.stepDistY\[1\]
+ _03051_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_26935_ _00845_ clknet_leaf_185_i_clk rbzero.tex_r1\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_21009_ _02097_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13900_ gpout0.vpos\[1\] _07704_ _07706_ _07707_ _07710_ _07711_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_199_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20594__A1 _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26866_ _00776_ clknet_leaf_165_i_clk rbzero.tex_r0\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14880_ rbzero.tex_b1\[39\] _08494_ _08321_ _08686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_230_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25817_ _06592_ _06600_ _06601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_214_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13831_ _07343_ _07642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_3_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26797_ _00707_ clknet_leaf_130_i_clk rbzero.tex_g1\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__19730__I _12501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23532__A1 _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16550_ _08117_ rbzero.debug_overlay.vplaneY\[-7\] _10002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_97_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25748_ _06491_ _06492_ _06532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__20876__I _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13762_ _07477_ _07572_ _07573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_193_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15501_ rbzero.spi_registers.texadd0\[12\] _09192_ _09196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_214_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16481_ _09919_ _09938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25679_ _06428_ _06462_ _06463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_210_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13693_ rbzero.tex_r0\[52\] _07487_ _07493_ _07504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18220_ _11344_ _11349_ _11300_ _11347_ _11363_ _11364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_194_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27418_ _01323_ clknet_leaf_85_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15432_ rbzero.spi_registers.buf_floor\[5\] _08885_ _09146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14576__A2 _07811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_18151_ _11280_ _11285_ _11289_ _11294_ _11295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_65_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27349_ _01254_ clknet_leaf_91_i_clk rbzero.wall_tracer.trackDistX\[-9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15363_ rbzero.spi_registers.buf_mapdyw\[1\] _09092_ _09095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17102_ rbzero.debug_overlay.vplaneX\[10\] _10481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14314_ _08123_ _08078_ _08124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18082_ _11191_ _11226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_135_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15294_ rbzero.map_overlay.i_othery\[2\] _09043_ _09044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17033_ rbzero.pov.ready_buffer\[26\] _10425_ _10429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14245_ _07998_ _08054_ _08055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_1_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14176_ _07423_ _07209_ _07986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_238_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14114__I _07526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13127_ rbzero.spi_registers.texadd3\[10\] _06921_ _06924_ rbzero.spi_registers.texadd2\[10\]
+ _06916_ rbzero.spi_registers.texadd1\[10\] _06941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_245_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18984_ rbzero.tex_g0\[28\] rbzero.tex_g0\[27\] _11861_ _11865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24012__A2 _08814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17935_ _08084_ _11047_ _11011_ _11079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_13058_ _06874_ _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14500__A2 _07898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23771__A1 _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22574__A2 _09974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17866_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] _11010_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_19605_ rbzero.wall_tracer.size\[5\] _12181_ _12376_ _12252_ _12377_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_16817_ rbzero.pov.ready_buffer\[69\] _10228_ _10229_ _10247_ _10248_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_108_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14264__A1 _08071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17797_ _10959_ rbzero.pov.ready_buffer\[56\] _10962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_220_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19536_ _12286_ _12307_ _12308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_191_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16748_ _10176_ _10180_ _10186_ _10187_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_221_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24258__I _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_159_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19467_ _12224_ _12238_ _12239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_16679_ _10112_ _10114_ _10120_ _10123_ _10124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__18256__I _11399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18418_ _11515_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19398_ _07774_ _07238_ _12170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_1_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18349_ _11475_ _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_200_i_clk clknet_5_12__leaf_i_clk clknet_leaf_200_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_155_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_20_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21360_ _02309_ _02442_ _02445_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__25579__A2 _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20311_ _12997_ _13004_ _01405_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21291_ _02146_ _02377_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_6_i_clk clknet_5_4__leaf_i_clk clknet_leaf_6_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_215_i_clk clknet_5_6__leaf_i_clk clknet_leaf_215_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_23030_ _03767_ _03759_ _03886_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_20242_ _12263_ _12917_ _13014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20173_ _12943_ _12944_ _12945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24981_ _05764_ _05574_ _05765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23762__A1 _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26720_ _00630_ clknet_leaf_29_i_clk rbzero.pov.ready_buffer\[50\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_192_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23932_ _10491_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input21_I i_reg_outs_enb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26651_ _00561_ clknet_leaf_145_i_clk rbzero.tex_b0\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23863_ _12214_ _04687_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25602_ _05234_ _06047_ _06385_ _06386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__17992__A2 _08374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22814_ _03668_ _03672_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_0_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26582_ _00492_ clknet_leaf_28_i_clk rbzero.pov.spi_buffer\[51\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23794_ _04628_ _04629_ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_196_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25533_ _06141_ _06179_ _06317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_175_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13812__B _07478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19733__A3 _12504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22745_ _03547_ _03604_ _03606_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14627__C _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25464_ _06235_ _06245_ _06246_ _06247_ _06248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_22676_ _11201_ _03522_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27203_ _01108_ clknet_leaf_75_i_clk rbzero.wall_tracer.size_full\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_192_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24415_ _05057_ _05177_ _05199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21627_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] _02701_
+ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25395_ _06170_ _06172_ _06178_ _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__19497__A2 _11991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27134_ _01044_ clknet_leaf_183_i_clk gpout1.clk_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24346_ _04907_ _05130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_21558_ _02539_ _02554_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22416__I _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20509_ _01596_ _01601_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_133_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22628__I0 rbzero.wall_tracer.texu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24277_ _04922_ _04860_ _05060_ _05061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27065_ _00975_ clknet_leaf_149_i_clk rbzero.tex_b1\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_21489_ _02453_ _02456_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_120_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14030_ _07830_ _07833_ _07837_ _07838_ _07839_ _07840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_91_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26016_ _06758_ rbzero.wall_tracer.rcp_fsm.o_data\[-4\] _06759_ _06793_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_23228_ _12212_ _02482_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14730__A2 _08298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19725__I _12496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23159_ _03899_ _04002_ _04014_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_227_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_227_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_246_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15981_ _09554_ _09555_ _09553_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_121_i_clk_I clknet_5_18__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13773__I _07583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24787__B _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17720_ _10906_ rbzero.pov.ready_buffer\[30\] _10911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14932_ _07431_ _08734_ _08737_ _08738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26918_ _00828_ clknet_leaf_126_i_clk rbzero.tex_r1\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_209_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_240_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17651_ _10857_ _10865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_215_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26849_ _00759_ clknet_leaf_192_i_clk rbzero.tex_r0\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14863_ _08665_ _08666_ _08668_ _08522_ _08532_ _08669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_230_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14246__A1 rbzero.debug_overlay.playerY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14246__B2 _07681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16602_ _08094_ _10031_ _10051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13814_ _07582_ _07625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17582_ rbzero.tex_b0\[48\] rbzero.tex_b0\[47\] _10817_ _10821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14794_ _07462_ _08599_ _08600_ _08601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_97_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19321_ _12122_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16533_ _09902_ _08100_ _09985_ _09986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13745_ rbzero.tex_r0\[43\] _07543_ _07556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25258__A1 _06037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19252_ _12072_ _12083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16464_ _09915_ _09918_ _09921_ rbzero.wall_tracer.rayAddendY\[-5\] _09922_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13676_ _07486_ _07487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_241_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18203_ _11332_ _11347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_100_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15415_ rbzero.spi_registers.buf_floor\[0\] _09131_ _09134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_100_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19183_ _12017_ _12026_ _12027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16395_ _09855_ _09867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__24481__A2 _05264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18134_ rbzero.wall_tracer.visualWallDist\[9\] _11278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_5_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_46_i_clk_I clknet_5_19__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15346_ _07754_ _09065_ _09082_ _09068_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_14_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_247_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18065_ rbzero.wall_tracer.trackDistY\[-10\] _11209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22619__I0 rbzero.wall_tracer.texu\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15277_ _09029_ _09030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16171__A1 _08948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17016_ _10415_ _10416_ _10414_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21047__A2 _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14228_ _08037_ _08009_ _08038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14159_ rbzero.color_floor\[1\] _07966_ _07670_ _07968_ _07969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_10_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18967_ _11855_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_237_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17918_ _08079_ _11001_ _11062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18898_ rbzero.traced_texa\[7\] _07267_ _11811_ _11812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_234_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17849_ _10994_ _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_240_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25497__A1 _06034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20860_ _12361_ _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_221_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15831__C _09441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14728__B _07867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19519_ _12249_ _11073_ _12291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20791_ _01870_ _01881_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22530_ rbzero.wall_tracer.visualWallDist\[-9\] _03436_ _03438_ rbzero.traced_texa\[-9\]
+ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14447__C _08222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22461_ _07147_ _07150_ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14019__I _07804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19479__A2 _11990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21412_ _02359_ _02365_ _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24200_ _04920_ _04851_ _04888_ _04960_ _04984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_173_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25180_ _05962_ _05963_ _05964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22392_ _03330_ _03333_ _03337_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24131_ _04833_ _04836_ _04838_ _04915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_135_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_21343_ _02421_ _02429_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_154_i_clk clknet_5_11__leaf_i_clk clknet_leaf_154_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_163_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24062_ _04844_ _04834_ _04845_ _04812_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_142_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24451__I _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21274_ _12698_ _02097_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14712__A2 _08518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23013_ _02251_ _03736_ _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_229_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20225_ _12992_ _12996_ _12997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_38_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_169_i_clk clknet_5_10__leaf_i_clk clknet_leaf_169_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20156_ _12660_ _12223_ _12928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_5_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14689__I _07822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13807__B _07462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23735__A1 _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20087_ _12806_ _12828_ _12830_ _12857_ _12858_ _12859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_24964_ _05686_ _05717_ _05746_ _05747_ _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__18206__A3 _11306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26703_ _00613_ clknet_leaf_61_i_clk rbzero.pov.ready_buffer\[33\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_222_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23915_ _04721_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_222_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24895_ _05623_ _05625_ _05679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__19280__I _12093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26634_ _00544_ clknet_leaf_162_i_clk rbzero.tex_b0\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_169_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23846_ _11142_ _03076_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15976__A1 _08965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26565_ _00475_ clknet_leaf_63_i_clk rbzero.pov.spi_buffer\[34\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20989_ _01729_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23777_ _04613_ _04614_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_200_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18914__A1 _11779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_107_i_clk clknet_5_31__leaf_i_clk clknet_leaf_107_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25516_ _05921_ _06039_ _06300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13530_ _07340_ _07341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22728_ rbzero.wall_tracer.trackDistX\[-1\] _01993_ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24626__I _05205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26496_ _00406_ clknet_leaf_55_i_clk rbzero.debug_overlay.facingY\[-4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25447_ _06228_ _06230_ _06231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13461_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] rbzero.texV\[7\]
+ _07272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_125_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22659_ _03526_ _03528_ _03530_ _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24463__A2 _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_173_Right_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15200_ _08967_ _08970_ _08971_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_152_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16180_ rbzero.spi_registers.buf_texadd1\[11\] _09696_ _09705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22474__A1 _10256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25378_ _06115_ _06116_ _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13392_ _07199_ _07203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15131_ _08913_ _08906_ _08909_ _08914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_27117_ _01027_ clknet_leaf_226_i_clk reg_gpout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24329_ _05044_ _05104_ _05112_ _05113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_229_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15062_ rbzero.spi_registers.spi_counter\[1\] _08854_ _08855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_27048_ _00958_ clknet_leaf_204_i_clk rbzero.wall_tracer.mapY\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14013_ rbzero.tex_r1\[27\] _07822_ _07823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_19870_ _12172_ _12639_ _12640_ _12641_ _12642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_242_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18821_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] _11749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_234_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_4__f_i_clk clknet_3_1_0_i_clk clknet_5_4__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_207_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18752_ rbzero.tex_r1\[43\] rbzero.tex_r1\[42\] _11703_ _11706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15964_ rbzero.spi_registers.spi_buffer\[5\] _09542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_234_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17703_ _10897_ rbzero.pov.ready_buffer\[24\] _10900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14915_ rbzero.tex_b1\[56\] _08698_ _08214_ _08721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18683_ rbzero.tex_r1\[13\] rbzero.tex_r1\[12\] _11666_ _11667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_215_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15895_ _08937_ _09476_ _09490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_216_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17634_ _10852_ rbzero.pov.ready_buffer\[1\] _10854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14846_ _08295_ _08648_ _08651_ _08652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_216_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20960__A1 _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25920__I _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17565_ _10811_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14777_ rbzero.tex_b0\[13\] _07930_ _08584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18905__A1 rbzero.traced_texa\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22765__B _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19304_ _12112_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16516_ _09966_ _09969_ _09970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13728_ _07443_ _07539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_168_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17496_ _10772_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19235_ rbzero.tex_b1\[1\] rbzero.tex_b1\[0\] _12073_ _12074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16447_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] _09905_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16392__A1 rbzero.spi_registers.buf_texadd3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13659_ _07450_ rbzero.row_render.texu\[1\] _07468_ _07469_ _07470_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xclkbuf_leaf_71_i_clk clknet_5_29__leaf_i_clk clknet_leaf_71_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19166_ _11950_ _11948_ _12010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22465__A1 _10255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16378_ rbzero.spi_registers.spi_buffer\[12\] _09853_ _09854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_205_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13678__I _07488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18117_ rbzero.debug_overlay.playerX\[0\] rbzero.map_rom.f4 _11261_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15329_ rbzero.spi_registers.buf_mapdy\[0\] _09060_ _09070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19097_ rbzero.debug_overlay.facingY\[-2\] _11919_ _11941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_170_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18048_ rbzero.wall_tracer.trackDistX\[-5\] _11192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__16695__A2 _10020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_86_i_clk clknet_5_25__leaf_i_clk clknet_leaf_86_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22768__A2 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14170__A3 _07979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20010_ _12694_ _12782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14458__A1 _08211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19999_ _12761_ _12766_ _12770_ _12771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21961_ _02994_ _02984_ _02995_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_206_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23700_ rbzero.wall_tracer.trackDistY\[-9\] _03037_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20912_ _02000_ _02001_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24680_ _05377_ _05464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21892_ _02811_ _02933_ _02934_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15958__A1 _09522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19149__A1 _08157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_24_i_clk clknet_5_20__leaf_i_clk clknet_leaf_24_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__24142__A1 _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20843_ _01931_ _01932_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_23631_ _04481_ _04482_ _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_230_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26350_ _00260_ clknet_leaf_2_i_clk rbzero.spi_registers.buf_texadd0\[18\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20774_ _01863_ _01864_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__20703__A1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23562_ _04413_ _04414_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_162_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16673__B _08096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25301_ _06084_ _06085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_130_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22513_ _03411_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23493_ _04252_ _04346_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26281_ _00191_ clknet_leaf_227_i_clk rbzero.spi_registers.buf_sky\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_39_i_clk clknet_5_16__leaf_i_clk clknet_leaf_39_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1_0_i_clk clknet_0_i_clk clknet_3_1_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_25232_ _06010_ _06015_ _06016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22444_ _02033_ _03373_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25163_ _05932_ _05935_ _05947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22375_ _03321_ _03250_ _12040_ _03193_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__26563__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24114_ _04897_ _04742_ _04898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__22208__A1 _11281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21326_ _02411_ _02412_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25094_ _05838_ _05853_ _05878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14697__A1 rbzero.tex_b0\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14921__B _08726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22759__A2 rbzero.wall_tracer.stepDistX\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24045_ _04813_ _04814_ _04815_ _04828_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_21257_ _02340_ _02343_ _01701_ _01726_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_53_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_224_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20208_ _12903_ _12921_ _12980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_183_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21188_ _02118_ _02274_ _02275_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15308__I _08986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20139_ rbzero.wall_tracer.size\[9\] _12640_ _12911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_148_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21754__B _09988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25996_ _06694_ _02997_ _06770_ _06774_ _06719_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_95_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23184__A2 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24381__A1 _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24947_ _05705_ _05706_ _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_225_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14700_ rbzero.tex_b0\[51\] _07938_ _08507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_242_Right_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_206_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15680_ _09327_ _09329_ _09325_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_206_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24878_ _05337_ _05329_ _05252_ _05607_ _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_202_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26617_ _00527_ clknet_leaf_169_i_clk rbzero.tex_b0\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14631_ rbzero.tex_g1\[37\] _07901_ _07630_ _08439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_23829_ _03296_ _03074_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_212_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14621__A1 _07803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17350_ rbzero.pov.spi_buffer\[41\] _10668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_138_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14562_ _07258_ _08371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_26548_ _00458_ clknet_leaf_25_i_clk rbzero.pov.spi_buffer\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_219_i_clk_I clknet_5_6__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16301_ rbzero.spi_registers.buf_texadd2\[17\] _09791_ _09796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13513_ _07266_ _07271_ _07312_ _07324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_17281_ _10614_ _10606_ _10616_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14493_ rbzero.tex_g0\[46\] _08298_ _08301_ _08302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_82_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26479_ _00389_ clknet_leaf_207_i_clk rbzero.debug_overlay.playerY\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_235_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19020_ _11885_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_180_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16232_ rbzero.spi_registers.buf_texadd2\[0\] _09743_ _09744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13444_ _07139_ _07254_ _07148_ _07255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_67_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14924__A2 _08222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16126__A1 rbzero.spi_registers.buf_texadd0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16163_ _08939_ _09687_ _09693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13375_ _07185_ _07186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15114_ rbzero.spi_registers.spi_counter\[5\] _08899_ _08900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_106_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17874__A1 rbzero.debug_overlay.facingX\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16094_ rbzero.spi_registers.buf_texadd0\[14\] _09633_ _09640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14831__B _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19922_ _12284_ _12694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15045_ _08836_ _08831_ _08835_ _08838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__13360__A1 _07171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18674__I0 rbzero.tex_r1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19853_ _12620_ _12624_ _12625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__21422__A2 _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15218__I _07166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18804_ _11449_ _11734_ _11735_ _11736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_247_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19784_ _12473_ _12554_ _12555_ _12556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_16996_ _10392_ _10401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__24372__A1 _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15947_ _08911_ _09528_ _09529_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18735_ _11696_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_222_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18666_ _11657_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_204_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15878_ _09476_ _09477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_84_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17617_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _10838_ _10841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14829_ _08630_ _08632_ _08634_ _08502_ _08285_ _08635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_18597_ _11617_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14612__B2 _08211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17548_ _10801_ _10802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_114_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19551__A1 _08076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15168__A2 _08940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17479_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _10760_ _10763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13179__A1 rbzero.spi_registers.texadd3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19218_ _12055_ _12059_ _12060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22438__A1 rbzero.wall_tracer.texu\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20490_ _01500_ _01514_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14915__A2 _08698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19149_ _08157_ _09991_ _11929_ _11993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_15_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21110__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22160_ _11287_ _03135_ _03130_ _11070_ _03114_ _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_41_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__26133__D _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21111_ _12498_ _02078_ _01723_ _12570_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_22091_ _03081_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__19606__A2 _12310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21042_ _02128_ _02129_ _02130_ _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_165_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25850_ _05212_ _06634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14032__I _07586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_168_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24801_ _05388_ _05534_ _05585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_242_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25781_ _06562_ _06564_ _06565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_198_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22993_ _02257_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_158_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24732_ _05512_ _05515_ _05516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21944_ _09925_ _02981_ _02091_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__13804__C _07589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21972__I0 rbzero.wall_tracer.rcp_fsm.o_data\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24115__A1 _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27451_ _01356_ clknet_leaf_72_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24663_ _05269_ _05270_ _05239_ _05447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14603__A1 rbzero.tex_g1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21875_ _10482_ _11069_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_210_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26402_ _00312_ clknet_leaf_248_i_clk rbzero.spi_registers.buf_texadd2\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_210_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23614_ _02260_ _04308_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27382_ _01287_ clknet_leaf_103_i_clk rbzero.wall_tracer.trackDistY\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__22677__A1 _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20826_ rbzero.wall_tracer.visualWallDist\[8\] _12228_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_148_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24130__A4 _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24594_ _05229_ _05377_ _05378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_166_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19542__A1 _08029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_26333_ _00243_ clknet_leaf_232_i_clk rbzero.spi_registers.buf_texadd0\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23545_ _04397_ _04298_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20757_ _01832_ _01847_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_119_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14367__B1 _08060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22429__A1 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26264_ _00174_ clknet_leaf_13_i_clk rbzero.spi_registers.texadd3\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23476_ _04222_ _02079_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20688_ _01773_ _01774_ _01772_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_134_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14906__A2 _08698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25215_ _05998_ _05999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14207__I _08016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22427_ rbzero.wall_tracer.texu\[2\] _03361_ _02715_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__21101__A1 _12465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14382__A3 _08191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26195_ _00105_ clknet_leaf_12_i_clk rbzero.spi_registers.texadd0\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25146_ _05913_ _05914_ _05928_ _05930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_13160_ _06946_ _06973_ _06974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_206_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21652__A2 _07772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22358_ _11376_ _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21309_ _02370_ _02395_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13091_ _06904_ _06905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25077_ _05830_ _05831_ _05859_ _05861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22289_ _10048_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24197__A4 _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24441__I2 _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13342__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_22__f_i_clk clknet_3_5_0_i_clk clknet_5_22__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_24028_ _04811_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__22601__A1 _07236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_218_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16850_ rbzero.pov.ready_buffer\[73\] _10274_ _10269_ _10276_ _10277_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__17084__A2 _10445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24354__A1 _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23157__A2 _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15801_ rbzero.spi_registers.texadd3\[17\] _09418_ _09419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_69_Left_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__24354__B2 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16781_ rbzero.debug_overlay.playerX\[-4\] _10203_ _10216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25979_ _10255_ _06759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21168__A1 _12210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13993_ _07329_ _07803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13781__I _07591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14842__A1 _08308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18520_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _11571_ _11574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15732_ rbzero.spi_registers.texadd2\[23\] _09362_ _09368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_66_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18451_ _11534_ _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_185_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15663_ _09305_ _09317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_237_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17402_ rbzero.pov.spi_buffer\[55\] _10697_ _10706_ _10707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14614_ rbzero.tex_g1\[0\] _07843_ _08422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18382_ rbzero.tex_g1\[12\] rbzero.tex_g1\[11\] _11491_ _11495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_201_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15594_ rbzero.spi_registers.texadd1\[12\] _09255_ _09265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_233_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19533__A1 _12300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14826__B _08280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17333_ rbzero.pov.spi_buffer\[37\] _10655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_200_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14545_ _08304_ _08345_ _08353_ _08354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__20143__A2 _12906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Left_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17264_ rbzero.pov.spi_buffer\[20\] _10603_ _10599_ _10604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21891__A2 _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14476_ _07551_ _08285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19003_ rbzero.tex_g0\[36\] rbzero.tex_g0\[35\] _11872_ _11876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16215_ rbzero.spi_registers.buf_texadd1\[20\] _09730_ _09731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13427_ _07237_ rbzero.trace_state\[2\] _07238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_141_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17195_ _08908_ _10552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16146_ _09679_ _09680_ _09678_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13358_ net41 _07159_ _07170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21643__A2 _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16332__I _09819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16077_ _08962_ _09624_ _09628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13289_ _07063_ _07089_ _07099_ _07102_ _07103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_110_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14280__C _08089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19905_ _12675_ _12676_ _12677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23396__A2 _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15028_ rbzero.spi_registers.spi_done _08821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__19643__I _10310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Left_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_19836_ _12242_ _12606_ _12607_ _12608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_209_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19767_ _12508_ _12538_ _12539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_224_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21159__A1 _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16979_ rbzero.pov.ready_buffer\[35\] _10383_ _10388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput3 i_debug_vec_overlay net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_160_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18718_ _11686_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19698_ _12267_ _12350_ _12469_ _12470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_79_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19772__A1 _12468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18649_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _11644_ _11647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_125_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21660_ _02724_ _08741_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14061__A2 _07832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_96_Left_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20611_ _12492_ _12496_ _01607_ _13025_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_21591_ _02646_ _02675_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20542_ _12688_ _12957_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23330_ _04181_ _04184_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_61_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21882__A2 _10466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23261_ _03902_ _03996_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20473_ _01479_ _01564_ _01565_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_94_i_clk_I clknet_5_19__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25000_ _05783_ _05308_ _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__24820__A2 _05429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22212_ _11279_ _03096_ _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23192_ _03667_ _03930_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22143_ rbzero.wall_tracer.visualWallDist\[-5\] _03100_ _03130_ _11074_ _03131_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20988__A4 _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_246_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__23387__A2 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22074_ rbzero.wall_tracer.stepDistY\[7\] _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26951_ _00861_ clknet_leaf_183_i_clk rbzero.tex_r1\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_77_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25902_ _06663_ _06684_ _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21025_ _02112_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_195_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__17066__A2 _10434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26882_ _00792_ clknet_leaf_164_i_clk rbzero.tex_r0\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_145_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25833_ _06611_ _06617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_25764_ _06547_ _06548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_230_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22976_ _03779_ _03832_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24715_ _05452_ _05486_ _05498_ _05499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_48_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21927_ _10484_ _02963_ _02966_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_25695_ _05980_ _05984_ _05978_ _06479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16577__A1 _08112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_178_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_219_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_178_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27434_ _01339_ clknet_leaf_82_i_clk rbzero.wall_tracer.rcp_fsm.operand\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24646_ _05428_ _05429_ _05430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21858_ _11072_ _09921_ _02902_ _10071_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__18318__A2 _11449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19366__I1 rbzero.tex_b1\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27365_ _01270_ clknet_leaf_101_i_clk rbzero.wall_tracer.trackDistX\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16329__A1 rbzero.spi_registers.buf_texadd3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20809_ _01791_ _01792_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_24577_ net90 _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_38_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21789_ _11080_ _09977_ _02838_ _09918_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_61_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_232_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26316_ _00226_ clknet_leaf_214_i_clk rbzero.spi_registers.buf_mapdx\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14330_ _08139_ _08140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_232_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23528_ _04377_ _04380_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21873__A2 _10087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27296_ _01201_ clknet_leaf_208_i_clk rbzero.row_render.size\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16861__B _10174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14261_ rbzero.debug_overlay.facingX\[-1\] _08071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26247_ _00157_ clknet_leaf_18_i_clk rbzero.spi_registers.texadd2\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23459_ _03849_ _03965_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16000_ _09568_ _09569_ _09565_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13212_ _07020_ _07026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22154__I _10151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26178_ _00088_ clknet_leaf_222_i_clk rbzero.color_floor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14192_ _07212_ _07224_ _07991_ _08002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_94_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13776__I _07586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25129_ _05894_ _05899_ _05913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13143_ _06956_ _06957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_143_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_210_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_210_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17951_ _11039_ _11086_ _11094_ _11095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13074_ _06889_ _06890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_218_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16902_ rbzero.debug_overlay.playerY\[-4\] _10316_ _10322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__18254__A1 _11134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17882_ _08072_ _11025_ _11026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24327__A1 _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19621_ _12309_ _12391_ _12392_ _12393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__13725__B _07337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16833_ _10258_ _10250_ _10262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13618__A2 _07428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19552_ _12323_ _11035_ _11036_ _12324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__14400__I _07498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16764_ _10182_ _10201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13976_ _07777_ _07780_ _07786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_233_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_220_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__19754__A1 _12382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23713__I _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14291__A2 _08036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23550__A2 _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18503_ _11563_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15715_ rbzero.spi_registers.buf_texadd2\[18\] _09353_ _09356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_17_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18807__I _11737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16695_ _10128_ _10020_ _10139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19483_ _12254_ _12255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_17_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17711__I _10843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15646_ rbzero.spi_registers.texadd2\[1\] _09303_ _09304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18434_ rbzero.tex_g1\[34\] rbzero.tex_g1\[33\] _11523_ _11525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19506__A1 rbzero.wall_tracer.visualWallDist\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18309__A2 _08753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23302__A2 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18365_ _11485_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_173_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16327__I _09814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15577_ rbzero.spi_registers.buf_texadd1\[8\] _09245_ _09252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17316_ _10640_ _10641_ _10642_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_116_i_clk_I clknet_5_19__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14528_ rbzero.tex_g0\[63\] _07894_ _08337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18296_ _11434_ _07707_ _08873_ _11435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__25055__A2 _05308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19638__I _12409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17247_ _10555_ _10591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18542__I _11564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14459_ rbzero.tex_g0\[11\] _07626_ _08268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_148_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17178_ rbzero.pov.spi_buffer\[0\] _10538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_40_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16129_ rbzero.spi_registers.buf_texadd0\[23\] _09655_ _09666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_162_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17048__A2 _10434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_127_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19819_ _12160_ _12279_ _12591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14806__A1 _07888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22830_ _02501_ _01919_ _02636_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_223_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14282__A2 _08078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22761_ _03619_ _03620_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_189_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17621__I rbzero.pov.spi_done vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24500_ _05283_ _05255_ _05284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21712_ _02769_ _11424_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25480_ _06101_ _06180_ _06260_ _06263_ _06264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_22692_ _11133_ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14034__A2 _07843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19348__I1 rbzero.tex_b1\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24431_ _05077_ _05093_ _05214_ _05215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_192_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21643_ rbzero.wall_tracer.rayAddendY\[-8\] _02689_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23779__B _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27150_ _01055_ clknet_leaf_183_i_clk reg_rgb\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20982__I _12464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24362_ _05144_ _05145_ _05080_ _05146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_214_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_173_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21574_ _02658_ _02553_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_214_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26101_ _00011_ clknet_leaf_243_i_clk rbzero.spi_registers.spi_counter\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23313_ _04061_ _04069_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20525_ _12399_ _01617_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_160_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27081_ _00991_ clknet_leaf_154_i_clk rbzero.tex_b1\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24293_ _04947_ _04838_ _05046_ _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_138_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16731__A1 _08182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26032_ _06781_ _06806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14913__C _08595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20456_ _01455_ _01457_ _01549_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_23244_ _01380_ _03852_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23175_ _03931_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_20387_ _01389_ _01480_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_203_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15298__A1 rbzero.map_overlay.i_othery\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22126_ _03083_ _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22702__I _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13848__A2 _07599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18236__A1 _08379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17039__A2 _10432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26934_ _00844_ clknet_leaf_174_i_clk rbzero.tex_r1\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_22057_ _03010_ _03060_ _03061_ _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20043__A1 _12750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21008_ rbzero.wall_tracer.stepDistX\[9\] _11389_ _02096_ _02097_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_26865_ _00775_ clknet_leaf_176_i_clk rbzero.tex_r0\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_25816_ _06595_ _06599_ _06600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13830_ _07341_ _07641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_203_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24629__I _05304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26796_ _00706_ clknet_leaf_130_i_clk rbzero.tex_g1\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_242_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14273__A2 _08045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25747_ _06480_ _06529_ _06530_ _06531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13761_ _07478_ _07530_ _07554_ _07571_ _07572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_69_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22959_ _02120_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19200__A3 _12043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15500_ _09193_ _09195_ _09191_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16480_ _09927_ _09932_ _09936_ _09937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25678_ _06442_ _06445_ _06461_ _06462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_13692_ rbzero.tex_r0\[53\] _07499_ _07503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27417_ _01322_ clknet_leaf_85_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_15431_ rbzero.color_floor\[5\] _08879_ _09145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23296__A1 _12676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24629_ _05304_ _05413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_214_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18150_ _11290_ _11291_ _11292_ _11293_ _11294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__20892__I _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27348_ _01253_ clknet_leaf_97_i_clk rbzero.wall_tracer.trackDistX\[-10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15362_ rbzero.mapdyw\[1\] _09090_ _09094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_96_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14981__C2 _07046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17101_ _10479_ _10480_ _10462_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14313_ _08122_ _08123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18081_ rbzero.wall_tracer.trackDistX\[-4\] _11225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_151_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15293_ _08878_ _09043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_27279_ _01184_ clknet_leaf_205_i_clk rbzero.wall_tracer.texu\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_22_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17032_ _08161_ _10423_ _10428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23909__S _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14244_ _08037_ _08004_ _08054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14175_ _07144_ _07189_ _07984_ _07985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_221_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15289__A1 rbzero.map_overlay.i_othery\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24313__B _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13126_ rbzero.texu_hot\[5\] _06939_ _06940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_245_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18983_ _11864_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__18227__A1 _09056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17934_ _08081_ _11077_ _11051_ _11078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__18227__B2 _07736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13057_ _06873_ _06874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_178_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17865_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] _11009_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16789__A1 _07699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_42_i_clk_I clknet_5_22__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15226__I _08916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19921__I _12692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19604_ _12289_ _11988_ _12290_ _12375_ _12376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_16816_ _10238_ _10245_ _10246_ _10247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17796_ _10946_ _10961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14264__A2 _08007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19535_ _12305_ _12306_ _12307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_89_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_187_Right_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_159_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13959_ net3 _07212_ _07215_ _07221_ _07770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_16747_ _09067_ _10187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_105_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19466_ _12237_ _12238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16678_ _10121_ _10122_ _10123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_202_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_235_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18417_ rbzero.tex_g1\[27\] rbzero.tex_g1\[26\] _11512_ _11515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15629_ _09254_ _09291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19397_ _12168_ _12169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_174_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18348_ _11474_ net22 _11475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15896__I _09429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18279_ _11404_ _11420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20310_ _12992_ _12996_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13527__A1 _07299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21290_ _01579_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20241_ _12592_ _13012_ _13013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21847__B _09899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20172_ _12773_ _12673_ _12944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22522__I _09972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18218__A1 _11338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16520__I _09973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18218__B2 _11331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24980_ _05569_ _05764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_243_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_196_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23931_ rbzero.wall_tracer.rcp_fsm.i_data\[-8\] _04728_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13365__B net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15136__I _08917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26650_ _00560_ clknet_leaf_145_i_clk rbzero.tex_b0\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23862_ _04689_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19718__A1 _12337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14255__A2 _08033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25601_ _05237_ _06385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input14_I i_gpout2_sel[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22813_ _03670_ _02603_ _03671_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_169_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23514__A2 _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26581_ _00491_ clknet_leaf_28_i_clk rbzero.pov.spi_buffer\[50\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23793_ _04628_ _04629_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_212_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_154_Right_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25532_ _06101_ _06180_ _06316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_175_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22744_ _11169_ _03605_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24385__S _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_175_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14007__A2 _07816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_177_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25463_ _06236_ _06239_ _06247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22675_ _02731_ _03543_ _03544_ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16952__A1 _07685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27202_ _01107_ clknet_leaf_75_i_clk rbzero.wall_tracer.size_full\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24414_ net67 _04995_ _05198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_192_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21626_ _09900_ _02701_ _02702_ _02703_ _02704_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_25394_ _06174_ _06177_ _06178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_191_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27133_ _01043_ clknet_leaf_224_i_clk gpout1.clk_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24345_ _05116_ _05128_ _05129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_21557_ _02585_ _02641_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_173_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20508_ _01599_ _01600_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_27064_ _00974_ clknet_leaf_150_i_clk rbzero.tex_b1\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24276_ _04967_ _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21488_ _02323_ _02564_ _02572_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26015_ _06785_ _06789_ _06791_ _06756_ _06792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_23227_ _03845_ _03709_ _03968_ _04082_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_160_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20439_ rbzero.wall_tracer.stepDistX\[4\] _01524_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23158_ _03997_ _04001_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_247_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_227_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_227_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22109_ _12216_ _03093_ _03094_ _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_101_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15980_ _08968_ _09551_ _09555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_219_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23089_ _03814_ _01920_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_247_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14931_ rbzero.color_floor\[5\] _07669_ _08198_ _08736_ _08737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_26917_ _00827_ clknet_leaf_126_i_clk rbzero.tex_r1\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_240_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_240_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14862_ rbzero.tex_b1\[2\] _08528_ _08667_ _08668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17650_ _10858_ _10563_ _10861_ _10864_ _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_26848_ _00758_ clknet_leaf_191_i_clk rbzero.tex_r0\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_230_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16601_ _08094_ _10038_ _10050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13813_ _07608_ _07624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_202_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17581_ _10820_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_138_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14793_ rbzero.tex_b0\[1\] _08209_ _08600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26779_ _00689_ clknet_leaf_122_i_clk rbzero.tex_g1\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__18357__I _11480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16532_ _08109_ rbzero.debug_overlay.vplaneY\[-9\] _09984_ _09985_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_35_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19320_ rbzero.tex_b1\[38\] rbzero.tex_b1\[37\] _12120_ _12122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13744_ _07468_ _07555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25258__A2 _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16463_ _09920_ _09921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19251_ _12082_ _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_167_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13675_ _07418_ _07486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_155_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15414_ rbzero.color_floor\[0\] _09129_ _09133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18202_ _11331_ _11343_ _11344_ _11345_ _11346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_100_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19182_ _12018_ _12024_ _12025_ _12026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_100_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16394_ rbzero.spi_registers.spi_buffer\[16\] _09865_ _09866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18133_ _11267_ _11268_ _11273_ _11276_ _11277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_15345_ rbzero.spi_registers.buf_mapdy\[4\] _09080_ _09082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25918__I _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18064_ _11204_ rbzero.wall_tracer.trackDistY\[-8\] _11206_ _11207_ _11208_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_0_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15276_ _09028_ _09029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_145_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17015_ rbzero.pov.ready_buffer\[43\] _10412_ _10416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19916__I _12472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14227_ _08024_ _08037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23438__I _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14158_ _07967_ _07668_ _07968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13109_ _06908_ _06914_ _06923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_238_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14089_ rbzero.tex_r1\[38\] _07898_ _07819_ _07899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18966_ rbzero.tex_g0\[20\] rbzero.tex_g0\[19\] _11851_ _11855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_238_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17917_ _11043_ _11059_ _11060_ _11061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18897_ rbzero.traced_texa\[6\] _07273_ _11810_ _11811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_206_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19651__I _12422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_201_Left_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_234_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17848_ _09892_ net28 _10994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__15434__A1 rbzero.spi_registers.vshift\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__18267__I _11409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17779_ _10944_ rbzero.pov.ready_buffer\[50\] _10950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_221_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19176__A2 _12007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19518_ _12179_ _12290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20790_ _01873_ _01880_ _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22180__A1 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19449_ _12162_ _12220_ _12221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16943__C _10357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22460_ _07150_ _08887_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_134_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14744__B _08355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21411_ _02360_ _02364_ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_211_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22391_ _01453_ _03332_ _03336_ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24130_ _04894_ _04902_ _04911_ _04913_ _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_TAPCELL_ROW_135_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21342_ _02423_ _02428_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25421__A2 _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24061_ rbzero.wall_tracer.rcp_fsm.operand\[8\] _04787_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14035__I _07483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21273_ _02197_ _02200_ _02198_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20246__A1 rbzero.wall_tracer.size\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23012_ _03725_ _03734_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20224_ _12993_ _12994_ _12995_ _12996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_38_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22252__I _11248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13874__I rbzero.debug_overlay.playerY\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__17346__I _10546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_223_Right_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20155_ _12663_ _12664_ _12927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_168_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20086_ _12761_ _12766_ _12759_ _12858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_24963_ _05691_ _05713_ _05714_ _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_51_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18206__A4 rbzero.map_rom.i_row\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23914_ _08812_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26702_ _00612_ clknet_leaf_62_i_clk rbzero.pov.ready_buffer\[32\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_222_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24894_ _05652_ _05676_ _05677_ _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_58_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_222_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26633_ _00543_ clknet_leaf_161_i_clk rbzero.tex_b0\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_240_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23845_ _04670_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_200_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26564_ _00474_ clknet_leaf_63_i_clk rbzero.pov.spi_buffer\[33\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23776_ _04613_ _04614_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_170_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20988_ _01947_ _01952_ _01954_ _01945_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_200_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25515_ _05321_ _06045_ _06299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22727_ _11134_ _02306_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_24_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26495_ _00405_ clknet_leaf_55_i_clk rbzero.debug_overlay.facingY\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16925__A1 _08018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25446_ _06227_ _06221_ _06225_ _06230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_13460_ _07267_ _07268_ _07270_ _07271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__23032__B _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22658_ _02730_ _03529_ _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_137_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21609_ _11456_ _02691_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25377_ _06148_ _06160_ _06161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_13391_ _07201_ _07202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22474__A2 _11449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22589_ _06908_ _03475_ _03477_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15130_ rbzero.spi_registers.spi_buffer\[1\] _08913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_27116_ net84 clknet_leaf_225_i_clk reg_gpout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_211_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24328_ _05105_ _05106_ _05110_ _05111_ _05112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_133_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_188_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_229_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25412__A2 _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15061_ _08851_ _08852_ _08845_ _08853_ _08854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_65_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27047_ _00957_ clknet_leaf_203_i_clk rbzero.wall_tracer.mapY\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24259_ _04871_ _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_239_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_248_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14012_ _07575_ _07822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21985__A1 rbzero.wall_tracer.size\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_242_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18820_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] _11748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_215_i_clk_I clknet_5_6__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17653__A2 rbzero.pov.ready_buffer\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_207_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18751_ _11705_ _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15963_ rbzero.spi_registers.buf_vshift\[5\] _09530_ _09541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21737__A1 _11107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19471__I rbzero.wall_tracer.stepDistX\[-5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17702_ _10884_ _10899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_216_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14914_ rbzero.tex_b1\[57\] _08526_ _08720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15894_ rbzero.spi_registers.buf_leak\[4\] _09482_ _09489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18682_ _11650_ _11666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_231_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17633_ _10849_ _10538_ _10851_ _10853_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_187_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14845_ _07814_ _08649_ _08650_ _08651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_230_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20960__A2 _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_5_i_clk clknet_5_4__leaf_i_clk clknet_leaf_5_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_203_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14776_ rbzero.tex_b0\[15\] _08554_ _08497_ _08583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17564_ rbzero.tex_b0\[40\] rbzero.tex_b0\[39\] _10807_ _10811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_214_i_clk clknet_5_6__leaf_i_clk clknet_leaf_214_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_216_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19303_ rbzero.tex_b1\[31\] rbzero.tex_b1\[30\] _12109_ _12112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16515_ _08102_ _09956_ _09968_ _09969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13727_ rbzero.tex_r0\[33\] _07537_ _07538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_196_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17495_ rbzero.tex_b0\[10\] rbzero.tex_b0\[9\] _10770_ _10772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16916__A1 _07713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19234_ _12072_ _12073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_128_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13658_ rbzero.row_render.texu\[4\] _07452_ _07469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16446_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] _09904_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18118__B1 _11260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_229_i_clk clknet_5_2__leaf_i_clk clknet_leaf_229_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_152_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16377_ _09819_ _09853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19165_ _12008_ _12009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22465__A2 _11444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13589_ _07367_ _07370_ _07365_ _07400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15328_ rbzero.map_overlay.i_mapdy\[0\] _09058_ _09069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18116_ rbzero.map_rom.a6 _11260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_117_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19096_ _11921_ _11938_ _11939_ _11940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_117_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__22217__A2 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18047_ rbzero.wall_tracer.trackDistY\[-4\] _11191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_10_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15259_ rbzero.map_overlay.i_otherx\[0\] _08879_ _09016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_10_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21976__A1 rbzero.wall_tracer.size\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20779__A2 _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19998_ _12764_ _12765_ _12770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23717__A2 _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18949_ _11829_ _11845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__21728__A1 _11344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21960_ rbzero.wall_tracer.size\[0\] _02992_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20911_ _12300_ _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21891_ _11069_ _02696_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16080__A1 _08965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23630_ _04381_ _04390_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20842_ _01829_ _01851_ _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__27250__D _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14630__A2 _07857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23561_ _04285_ _04288_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20773_ _12659_ _01641_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_147_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25300_ _05869_ _05909_ _06084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22512_ _03409_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26280_ _00190_ clknet_leaf_244_i_clk rbzero.spi_registers.texadd3\[23\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23492_ _04342_ _04345_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25231_ _06014_ _06015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22443_ _03384_ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__19857__B1 _12527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_164_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25162_ _05871_ _05908_ _05942_ _05946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_162_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22374_ _03320_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19556__I _12327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24113_ _04737_ _04869_ _04811_ _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_5_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21325_ _01483_ _12647_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14146__B2 _07955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25093_ _05836_ _05875_ _05876_ _05877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_107_Left_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14921__C _08357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24044_ rbzero.wall_tracer.rcp_fsm.operand\[4\] rbzero.wall_tracer.rcp_fsm.operand\[3\]
+ rbzero.wall_tracer.rcp_fsm.operand\[2\] rbzero.wall_tracer.rcp_fsm.operand\[1\]
+ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_21256_ _02341_ _02342_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__21967__A1 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25158__A1 _05912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_224_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20207_ _12877_ _12924_ _12978_ _12979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_183_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_224_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21187_ _02119_ _02121_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_159_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23708__A2 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20138_ _12907_ _11981_ _12909_ _12910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_25995_ _06773_ _06774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_148_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21719__A1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24946_ _05724_ _05728_ _05613_ _05729_ _05730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_20069_ _12750_ _12841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_clkbuf_leaf_89_i_clk_I clknet_5_24__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24877_ _05613_ _05660_ _05614_ _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_202_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_116_Left_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_202_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14630_ rbzero.tex_g1\[36\] _07857_ _08438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23828_ _03296_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_26616_ _00526_ clknet_leaf_168_i_clk rbzero.tex_b0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_185_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22144__A1 _11990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_198_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14561_ _07971_ _08369_ _08370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26547_ _00457_ clknet_leaf_24_i_clk rbzero.pov.spi_buffer\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23759_ rbzero.wall_tracer.trackDistY\[-2\] _03056_ _04592_ _04600_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18899__A1 _11769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16300_ _09792_ _09794_ _09795_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13512_ _07322_ _07323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__19560__A2 _12271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17280_ rbzero.pov.spi_buffer\[24\] _10615_ _10612_ _10616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14492_ rbzero.tex_g0\[47\] _08300_ _08301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_26478_ _00388_ clknet_leaf_211_i_clk rbzero.debug_overlay.playerY\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_235_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16231_ _09742_ _09743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25429_ _06204_ _06211_ _06212_ _06213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13443_ _07079_ _07254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16155__I _09675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16162_ rbzero.spi_registers.buf_texadd1\[6\] _09685_ _09692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13374_ net21 _07185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_125_Left_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__19466__I _12237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14137__A1 rbzero.tex_r1\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15113_ _08865_ _08898_ _08899_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_134_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16093_ _09638_ _09639_ _09637_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_239_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14688__A2 _08494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19921_ _12692_ _12693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15044_ _08831_ _08835_ _08836_ _08837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21958__A1 _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_248_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19852_ _12621_ _12622_ _12623_ _12624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__19871__I0 rbzero.wall_tracer.stepDistY\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18674__I1 rbzero.tex_r1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_247_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18803_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] _11735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19783_ _12402_ _12553_ _12477_ _12482_ _12555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__19415__B _12182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16995_ _10345_ _10399_ _10400_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_223_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13112__A2 _06922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24372__A2 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18734_ rbzero.tex_r1\[35\] rbzero.tex_r1\[34\] _11693_ _11696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15946_ rbzero.spi_registers.buf_vshift\[0\] _09527_ _09478_ _09529_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_134_Left_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18665_ rbzero.tex_r1\[5\] rbzero.tex_r1\[4\] _11656_ _11657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15877_ _08829_ _09444_ _09476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_153_i_clk clknet_5_11__leaf_i_clk clknet_leaf_153_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__16062__A1 _09542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17616_ _10840_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14828_ rbzero.tex_b1\[29\] _08279_ _08633_ _08634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18596_ rbzero.tex_r0\[40\] rbzero.tex_r0\[39\] _11613_ _11617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_148_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17547_ _10758_ _10801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23883__A1 rbzero.wall_tracer.rcp_fsm.o_data\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22686__A2 _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14759_ _08560_ _08561_ _08563_ _08564_ _08565_ _08566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_59_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_168_i_clk clknet_5_10__leaf_i_clk clknet_leaf_168_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17478_ _10762_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_15_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13179__A2 _06922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14376__A1 _07694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19217_ _12057_ _12052_ _12058_ _12059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16429_ _09457_ _09886_ _09890_ _08888_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__14376__B2 _07687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_143_Left_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19148_ _08156_ _10008_ _11931_ _11992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_132_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24282__I _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19079_ _08161_ rbzero.wall_tracer.rayAddendY\[3\] _11923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15876__A1 _09462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21110_ _01947_ _01951_ _01944_ _01834_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_160_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22090_ _03080_ _03083_ _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__15409__I _09074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21041_ _02010_ _02023_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_106_i_clk clknet_5_30__leaf_i_clk clknet_leaf_106_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__18665__I1 rbzero.tex_r1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20621__A1 _12706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24800_ _05578_ _05582_ _05583_ _05584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_226_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25780_ _06051_ _05970_ _06563_ _06385_ _06564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_119_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_213_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22992_ _03844_ _03849_ _02524_ _02336_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA_clkbuf_leaf_90_i_clk_I clknet_5_24__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14851__A2 _07906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24731_ _05513_ _05514_ _05515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_21943_ rbzero.wall_tracer.rcp_done _11392_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_119_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21972__I1 rbzero.wall_tracer.size\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27450_ _01355_ clknet_leaf_74_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_143_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24662_ _05420_ _05314_ _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_173_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21874_ _10072_ _02909_ _02916_ _02887_ _02917_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_221_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26401_ _00311_ clknet_leaf_248_i_clk rbzero.spi_registers.buf_texadd2\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23613_ _04399_ _04427_ _04464_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_27381_ _01286_ clknet_leaf_104_i_clk rbzero.wall_tracer.trackDistY\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20825_ _01831_ _01850_ _01848_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__23874__A1 rbzero.wall_tracer.stepDistX\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24593_ net47 _05245_ _05377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26332_ _00242_ clknet_leaf_242_i_clk rbzero.spi_registers.buf_texadd0\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23544_ _04284_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20756_ _01837_ _01846_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_46_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14367__A1 _08175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26263_ _00173_ clknet_leaf_13_i_clk rbzero.spi_registers.texadd3\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23475_ _04220_ _04223_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22429__A2 _07705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20687_ _09939_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_163_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25214_ _05823_ _05997_ _05815_ _05998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_135_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22426_ _03351_ _03368_ _03369_ _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26194_ _00104_ clknet_leaf_214_i_clk rbzero.spi_registers.texadd0\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14119__A1 rbzero.tex_r1\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25145_ _05913_ _05914_ _05928_ _05929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22357_ _02779_ _03248_ _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21308_ _02373_ _02394_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25076_ _05830_ _05831_ _05859_ _05860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_13090_ gpout0.hpos\[0\] _06904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22288_ _11288_ _03250_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13878__B1 _07676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24441__I3 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24027_ _04810_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13342__A2 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21239_ _02182_ _02242_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__18281__A2 _11420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15800_ _09037_ _09418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_70_i_clk clknet_5_29__leaf_i_clk clknet_leaf_70_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__24354__A2 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23980__B _09113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13992_ _07326_ _07802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16780_ _10202_ _10215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25978_ _06901_ _06758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21168__A2 _13012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14379__B _07195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15731_ _09366_ _09367_ _09361_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24929_ _05693_ _05708_ _05709_ _05711_ _05712_ _05713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_TAPCELL_ROW_66_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18450_ rbzero.tex_g1\[41\] rbzero.tex_g1\[40\] _11533_ _11534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_213_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15662_ rbzero.spi_registers.texadd2\[5\] _09315_ _09316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_196_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_237_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_85_i_clk clknet_5_25__leaf_i_clk clknet_leaf_85_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17401_ _10705_ _10706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14613_ rbzero.tex_g1\[1\] _07878_ _08421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15593_ _09263_ _09264_ _09253_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18381_ _11494_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__23865__A1 _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14544_ _08346_ _08349_ _08352_ _08353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17332_ _10652_ _10653_ _10654_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_154_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24409__A3 _05139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14358__A1 _08089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14475_ _07642_ _08284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17263_ _10602_ _10603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_181_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25198__I _05321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19002_ _11875_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13426_ rbzero.trace_state\[3\] _07237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16214_ _09670_ _09730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17194_ rbzero.pov.spi_buffer\[2\] _10551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__24290__A1 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16145_ _08913_ _09676_ _09680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17709__I _10847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13357_ _07156_ _07162_ _07163_ _07168_ _07169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_87_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16076_ rbzero.spi_registers.buf_texadd0\[9\] _09622_ _09627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_23_i_clk clknet_5_20__leaf_i_clk clknet_leaf_23_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13288_ _07101_ _07102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_121_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_19904_ _12430_ _12676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19924__I _12596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15027_ _08820_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_110_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_248_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__24051__B _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19835_ _12537_ _12605_ _12607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_112_i_clk_I clknet_5_31__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_38_i_clk clknet_5_7__leaf_i_clk clknet_leaf_38_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_19766_ _12510_ _12532_ _12538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_30_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16978_ _08081_ _10381_ _10387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput4 i_gpout0_sel[0] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14833__A2 _08568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18717_ rbzero.tex_r1\[28\] rbzero.tex_r1\[27\] _11682_ _11686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_160_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15929_ _09515_ _09508_ _09516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19697_ rbzero.wall_tracer.stepDistX\[-8\] _11384_ _12469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19772__A2 _12485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18648_ _11646_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_125_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22108__A1 _09956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22108__B2 _12595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14597__A1 _07480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18579_ _11564_ _11607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_176_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20610_ _12731_ _01701_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21590_ _02656_ _02661_ _02674_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_151_Left_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_188_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20541_ _01632_ _01633_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_144_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23260_ _03902_ _03996_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_37_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22525__I _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20472_ _01481_ _01563_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_171_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22211_ _03176_ _03186_ _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_41_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23191_ _03943_ _03953_ _03951_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_30_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22142_ _03083_ _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__20045__I _12789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22073_ _03019_ _03060_ _03071_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26950_ _00860_ clknet_leaf_181_i_clk rbzero.tex_r1\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__21398__A2 _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25901_ _06683_ _06615_ _06684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21024_ _12427_ _12433_ _01917_ _02112_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_26881_ _00791_ clknet_leaf_164_i_clk rbzero.tex_r0\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14978__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13882__I rbzero.debug_overlay.playerY\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15077__A2 _08751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25832_ _06571_ _06590_ _06616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14824__A2 _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25763_ _06514_ _06545_ _06546_ _06547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_22975_ _03779_ _03832_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__16026__A1 _09522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__26089__A2 _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24714_ _05384_ _05453_ _05485_ _05498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21926_ _02947_ _02964_ _02965_ _02941_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_25694_ _05235_ _06195_ _06478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_241_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_219_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_219_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27433_ _01338_ clknet_leaf_83_i_clk rbzero.wall_tracer.rcp_fsm.operand\[9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_195_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24645_ net72 _05360_ _05429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__14588__B2 _08211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21857_ _02900_ _02901_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_210_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20808_ _01785_ _01889_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24576_ _05349_ _05355_ _05359_ _05360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_27364_ _01269_ clknet_leaf_102_i_clk rbzero.wall_tracer.trackDistX\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_239_Left_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_61_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21788_ _10463_ _02837_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_194_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21322__A2 _12207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23527_ _04378_ _04379_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_26315_ _00225_ clknet_leaf_232_i_clk rbzero.spi_registers.buf_vinf vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20739_ _01724_ _01731_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_191_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27295_ _01200_ clknet_leaf_210_i_clk rbzero.row_render.size\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26246_ _00156_ clknet_leaf_18_i_clk rbzero.spi_registers.texadd2\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14260_ _08027_ _08052_ _08056_ _08069_ _08070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_23458_ _03846_ _04259_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13211_ rbzero.spi_registers.texadd0\[22\] _07025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22409_ _01776_ _03353_ _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26177_ _00087_ clknet_leaf_223_i_clk rbzero.color_floor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14760__A1 rbzero.tex_b0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13563__A2 _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14191_ _07999_ _08000_ _08001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_23389_ _04124_ _04006_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14381__C _07222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20833__A1 _12432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25128_ _05873_ _05906_ _05911_ _05912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_13142_ rbzero.texu_hot\[2\] _06955_ _06956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_210_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_210_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13315__A2 _07111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25059_ _05783_ _05641_ _05842_ _05843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17950_ _11037_ _11091_ _11093_ _11094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_57_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13073_ _06861_ _06889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_248_Left_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16901_ rbzero.pov.ready_buffer\[50\] _10274_ _10321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_168_Right_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17881_ rbzero.wall_tracer.rayAddendX\[5\] _11025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18254__A2 _11397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13792__I _07331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19620_ _12373_ _12390_ _12392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20061__A2 _12224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24327__A2 _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16832_ _10258_ _10250_ _10261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14276__B1 _08040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24878__A3 _05252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19551_ _08076_ _11092_ _12323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_221_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16763_ rbzero.debug_overlay.playerX\[-5\] _10200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_13975_ _07200_ _07079_ _07785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16017__A1 _08962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21010__A1 _12836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18502_ net25 rbzero.tex_g1\[63\] _11559_ _11563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_244_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15714_ rbzero.spi_registers.texadd2\[18\] _09350_ _09355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19482_ _07237_ _08373_ _07239_ _12254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_17_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16694_ _09953_ _10130_ _10135_ _10137_ _10138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_107_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18433_ _11524_ _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14579__A1 rbzero.tex_g1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15645_ _09302_ _09303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_200_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18364_ rbzero.tex_g1\[4\] rbzero.tex_g1\[3\] _11481_ _11485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15576_ rbzero.spi_registers.texadd1\[8\] _09243_ _09251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22510__A1 rbzero.wall_tracer.texu\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__22510__B2 _08360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17315_ rbzero.pov.spi_buffer\[33\] _10638_ _10635_ _10642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14527_ rbzero.tex_g0\[62\] _07901_ _08336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18295_ _07979_ _11434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17246_ rbzero.pov.spi_buffer\[15\] _10590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__23066__A2 _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14458_ _08211_ _08265_ _08266_ _08267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_142_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13409_ _07219_ _07220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_148_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14389_ _07430_ _08198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17177_ _10518_ _10534_ _10537_ _10512_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_109_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16128_ _09664_ _09665_ _09661_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19690__A1 _12417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19654__I _12397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13306__A2 _07108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14503__A1 _08245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16059_ _09614_ _09615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_162_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_127_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25515__A1 _05321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19818_ _12381_ _12590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_127_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19749_ _12520_ _12521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22760_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] _03613_
+ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_116_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_140_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13490__A1 _07299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21711_ _08171_ _02731_ _02770_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22691_ _11195_ _12266_ _03558_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_177_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24430_ _05045_ _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14466__C _07802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21642_ _08099_ rbzero.wall_tracer.rayAddendY\[-8\] _09904_ _02717_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_176_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24361_ _04720_ _05131_ _05037_ _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21573_ _02542_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14038__I _07343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_214_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18181__A1 rbzero.map_overlay.i_othery\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26100_ _00010_ clknet_leaf_227_i_clk gpout0.vinf vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_90_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23312_ _04149_ _04166_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20524_ rbzero.wall_tracer.stepDistY\[5\] _01530_ _01526_ _01616_ _01617_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_7_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27080_ _00990_ clknet_leaf_155_i_clk rbzero.tex_b1\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_105_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24292_ _05075_ _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_145_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26031_ _05028_ _06803_ _06804_ _05022_ _06805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_160_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23243_ _02404_ _02546_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20455_ _01544_ _01548_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23174_ _03919_ _03927_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19681__A1 _12425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20386_ _12933_ _12963_ _01391_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_203_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22125_ rbzero.wall_tracer.visualWallDist\[-8\] _03105_ _03115_ _03116_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_246_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22568__A1 _11282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22568__B2 rbzero.traced_texa\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22056_ rbzero.wall_tracer.stepDistY\[0\] _03054_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19433__A1 _07708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26933_ _00843_ clknet_leaf_174_i_clk rbzero.tex_r1\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_234_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13826__B _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16247__A1 _08922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21007_ _11389_ _02095_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_215_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26864_ _00774_ clknet_leaf_166_i_clk rbzero.tex_r0\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_25815_ _06582_ _06598_ _06599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_173_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_230_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26795_ _00705_ clknet_leaf_131_i_clk rbzero.tex_g1\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_98_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13760_ _07555_ _07569_ _07570_ _07571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25746_ _06479_ _06529_ _06493_ _06530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_186_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22958_ _03814_ _03815_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13481__A1 rbzero.traced_texVinit\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21909_ _02950_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13691_ rbzero.tex_r0\[54\] _07487_ _07501_ _07502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25677_ _06446_ _06460_ _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_211_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22889_ _03746_ _03747_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15222__A2 _08975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27416_ _01321_ clknet_leaf_85_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15430_ _09143_ _09144_ _09112_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24628_ _05411_ _05348_ _05412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__23296__A2 _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15361_ _09091_ _09093_ _09089_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24559_ _05291_ _05294_ _05342_ _05343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_27347_ _01252_ clknet_leaf_97_i_clk rbzero.wall_tracer.trackDistX\[-11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14981__A1 _06892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14981__B2 _07153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18172__A1 rbzero.map_overlay.i_othery\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17100_ rbzero.pov.ready_buffer\[20\] _10460_ _10480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14312_ _08121_ _08122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_18080_ _11194_ _11223_ _11224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15292_ _09040_ _09041_ _09042_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27278_ _01183_ clknet_leaf_119_i_clk rbzero.wall_tracer.texu\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_22_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_237_Right_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_22_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17031_ _06899_ _10427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14243_ _07997_ _08043_ _08053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_180_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26229_ _00139_ clknet_leaf_1_i_clk rbzero.spi_registers.texadd1\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14174_ _06862_ _07189_ _07984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19474__I _12179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13125_ _06912_ _06937_ _06938_ _06939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__25745__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18982_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _11861_ _11864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_245_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17933_ _11014_ _11077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18227__A2 _11343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13056_ _06872_ _06873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_237_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13736__B _07546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17864_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] _11008_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_17_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19603_ _12176_ _11071_ _12375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16815_ _10243_ _10239_ _10246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_219_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17795_ _10958_ _10708_ _10954_ _10960_ _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_75_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19534_ _12265_ _12285_ _12306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16746_ rbzero.pov.ready_buffer\[60\] _10183_ _10179_ _10185_ _10186_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_191_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13958_ _07258_ _07674_ _07717_ _07768_ _07242_ _07769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_TAPCELL_ROW_89_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19465_ _12236_ _12237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16677_ _10115_ _10116_ _10119_ _10122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_33_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13889_ _07699_ _07700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_201_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18416_ _11514_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__25160__B _05943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15628_ _09287_ _09288_ _09290_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19396_ _12167_ _12168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_174_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13224__A1 _07026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_228_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21298__A1 _12689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18347_ _08806_ _11474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15559_ rbzero.spi_registers.texadd1\[4\] _09230_ _09238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18278_ rbzero.wall_tracer.mapX\[9\] _11419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17910__A1 _08085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13697__I _07481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_204_Right_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17229_ rbzero.pov.spi_buffer\[11\] _10568_ _10577_ _10578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20240_ _12644_ _13012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_24_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_i_clk_I i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20171_ _12867_ _12940_ _12942_ _12943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_244_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__18218__A2 _11360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_23930_ _04733_ _04725_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_243_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23861_ _04684_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18728__I _11649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25600_ _06362_ _06363_ _06384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22812_ _02601_ _02602_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__19718__A2 _12339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23792_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.stepDistY\[2\] _04623_
+ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_168_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13463__A1 rbzero.traced_texVinit\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26580_ _00490_ clknet_leaf_28_i_clk rbzero.pov.spi_buffer\[49\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_196_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25531_ _06265_ _06314_ _06315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_22743_ _02766_ _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_175_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_175_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22694__B _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15152__I _08931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25462_ _06214_ _06215_ _06217_ _06246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_181_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22674_ _02737_ _01453_ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_164_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13215__A1 rbzero.spi_registers.texadd3\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27201_ _01106_ clknet_leaf_75_i_clk rbzero.wall_tracer.size_full\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24413_ _05056_ _05197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21625_ rbzero.wall_tracer.rayAddendX\[-8\] _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_25393_ _06119_ _06175_ _06176_ _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_47_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24344_ _05086_ _05119_ _05125_ _05127_ _05128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_192_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27132_ _01042_ clknet_leaf_225_i_clk gpout0.clk_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_21556_ _02617_ _02640_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17901__A1 rbzero.debug_overlay.facingX\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20507_ _12626_ _13025_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27063_ _00973_ clknet_leaf_151_i_clk rbzero.tex_b1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__25975__A1 _06737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24275_ _05036_ _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21487_ _02450_ _02563_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26014_ _06745_ _06734_ _06790_ _05242_ _06791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_23226_ _03967_ _03970_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20438_ rbzero.wall_tracer.stepDistY\[4\] _01525_ _01526_ _01531_ _01532_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_28_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21461__A1 _12383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23157_ _04008_ _04009_ _04012_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_28_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20369_ _01398_ _01443_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_246_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_227_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22108_ _09956_ _03085_ _03100_ _12595_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_8_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_227_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23088_ _03824_ _03944_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_2_0_i_clk_I clknet_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22039_ _03048_ _03039_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14930_ _08735_ _07669_ _08736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26916_ _00826_ clknet_leaf_126_i_clk rbzero.tex_r1\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_209_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_i_clk_I clknet_5_4__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_159_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26847_ _00757_ clknet_leaf_192_i_clk rbzero.tex_r0\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14861_ rbzero.tex_b1\[3\] _08529_ _08667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_240_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16600_ _10048_ _10049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13812_ _07609_ _07622_ _07478_ _07623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_242_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17580_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _10817_ _10820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14792_ rbzero.tex_b0\[0\] _08247_ _08599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26778_ _00688_ clknet_leaf_122_i_clk rbzero.tex_g1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__22713__A1 _11190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16531_ _09978_ _09984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_86_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25729_ _06509_ _06511_ _06513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_230_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13743_ _07480_ _07553_ _07554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17196__A2 _10547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19250_ rbzero.tex_b1\[8\] rbzero.tex_b1\[7\] _12078_ _12082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_195_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16462_ _09919_ _09920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_5_9__f_i_clk_I clknet_3_2_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24466__A1 _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13674_ rbzero.tex_r0\[51\] _07484_ _07485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_211_i_clk_I clknet_5_16__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18201_ _11315_ _11259_ _11345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_15413_ _09130_ _09132_ _09112_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14954__A1 _07164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19181_ _11354_ _12008_ _12025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_100_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16393_ _09818_ _09865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_100_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18145__A1 _11286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18132_ rbzero.wall_tracer.mapX\[7\] rbzero.wall_tracer.mapX\[6\] _11274_ _11275_
+ _11276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_183_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15344_ _07757_ _09065_ _09081_ _09068_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__18306__C _10992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18063_ rbzero.wall_tracer.trackDistY\[-9\] _11207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14406__I _08214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15275_ _08876_ _09028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_184_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17014_ _08076_ _10410_ _10415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14226_ _08035_ _08036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__19645__A1 _08062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22623__I _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14850__B _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14157_ rbzero.color_sky\[1\] _07967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_238_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15131__A1 _08913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13108_ _06921_ _06922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_238_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14088_ _07632_ _07898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18965_ _11854_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__19932__I _12553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15237__I _08951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17916_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] _11060_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_237_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18896_ _11807_ _11809_ _11810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23454__I _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17847_ _10993_ _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_206_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17778_ _10943_ _10690_ _10947_ _10949_ _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_88_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19517_ _12175_ _12289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_53_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16729_ _10167_ _10170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_221_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19448_ rbzero.wall_tracer.stepDistY\[-10\] _12169_ _12219_ _12220_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__15198__A1 _08968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19379_ net26 rbzero.tex_b1\[63\] _12151_ _12155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__18283__I _11399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18136__A1 _11278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_211_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21410_ _02382_ _02392_ _02390_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_174_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_211_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_170_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22390_ _12577_ _08182_ _03334_ _03335_ _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__19884__A1 _10231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23680__A2 _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21341_ _02424_ _02427_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_135_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21691__A1 _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__27248__D _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24060_ _04830_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21272_ _02357_ _02217_ _02358_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__19636__A1 rbzero.debug_overlay.playerX\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15856__B _08909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23011_ _03727_ _03868_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17627__I _10847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25709__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20223_ _12421_ _12296_ _12995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21443__A1 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25844__I _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20154_ _12668_ _12728_ _12926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_168_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16870__A1 rbzero.pov.ready_buffer\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20085_ _12831_ _12827_ _12856_ _12857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_24962_ _05736_ _05743_ _05744_ _05745_ _05746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__23364__I _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_160_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26701_ _00611_ clknet_leaf_62_i_clk rbzero.pov.ready_buffer\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23913_ _04719_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_222_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24893_ _05675_ _05672_ _05674_ _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__17362__I _10665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15425__A2 _08879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16622__B2 _10036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26632_ _00542_ clknet_leaf_161_i_clk rbzero.tex_b0\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_170_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23844_ _11142_ _03076_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13436__A1 _07244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23499__A2 _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23775_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] _04610_
+ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26563_ _00473_ clknet_leaf_63_i_clk rbzero.pov.spi_buffer\[32\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20987_ _12732_ _02075_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_200_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25514_ _05235_ _06102_ _06298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15189__A1 _08962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_22726_ _03547_ _03588_ _03589_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26494_ _00404_ clknet_leaf_55_i_clk rbzero.debug_overlay.facingY\[-6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19289__I _12093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22657_ _12943_ _12944_ _12866_ _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_25445_ _06181_ _06103_ _06229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18193__I _11112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21608_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13390_ _07199_ _07200_ _07201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_5_16__f_i_clk clknet_3_4_0_i_clk clknet_5_16__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25376_ _06151_ _06158_ _06159_ _06160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_22588_ rbzero.wall_tracer.wall\[0\] _03476_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_211_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27115_ _01025_ clknet_leaf_141_i_clk rbzero.tex_b1\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_65_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24327_ _05065_ _05067_ _05069_ _05041_ _05111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_21539_ _02277_ _02377_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14226__I _08035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_85_i_clk_I clknet_5_25__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_229_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15060_ _08830_ _08835_ _08840_ _08844_ _08853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_24258_ _04877_ _05042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_161_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27046_ _00956_ clknet_leaf_160_i_clk rbzero.tex_g0\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_239_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14011_ _07341_ _07821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_189_Left_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23209_ _01642_ _03814_ _04058_ _04064_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_24189_ _04968_ _04969_ _04971_ _04972_ _04973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_248_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_242_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22599__B _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16861__A1 _08049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_207_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18750_ rbzero.tex_r1\[42\] rbzero.tex_r1\[41\] _11703_ _11705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_207_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15962_ _09539_ _09540_ _09536_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_234_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17701_ _10896_ _10614_ _10892_ _10898_ _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_175_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14913_ _08715_ _08716_ _08718_ _08558_ _08595_ _08719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_18681_ _11665_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_234_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15893_ _09487_ _09488_ _09473_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20945__B1 _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_216_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17632_ _10852_ rbzero.pov.ready_buffer\[0\] _10853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_203_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14844_ rbzero.tex_b1\[20\] _07595_ _08650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_198_Left_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_102_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17563_ _10810_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14775_ rbzero.tex_b0\[14\] _08494_ _08582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19302_ _12111_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16514_ _09967_ _09968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13726_ _07531_ _07537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17494_ _10771_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19233_ _12071_ _12072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16445_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] _09903_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13657_ _07328_ _07468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18118__A1 rbzero.debug_overlay.playerX\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18118__B2 _07681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19164_ _12007_ _12008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16376_ rbzero.spi_registers.buf_texadd3\[12\] _09851_ _09852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_152_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13588_ _07062_ _07397_ _07399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_18115_ rbzero.map_rom.i_col\[4\] _11259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_15327_ _07740_ _09065_ _09066_ _09068_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__21673__A1 _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19095_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] _11939_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14136__I _07488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18046_ rbzero.wall_tracer.trackDistX\[-4\] _11190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__14155__A2 _07960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15258_ _08811_ _09015_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23414__A2 _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14580__B _07646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21425__A1 _12689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14209_ _07713_ _08007_ _08011_ _07698_ _08017_ _08018_ _08019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_15189_ _08962_ _08952_ _08963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19997_ _12537_ _12605_ _12242_ _12769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__15655__A2 _09306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16852__A1 _08175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18948_ _11844_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21728__A2 _11420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18879_ _11795_ _11796_ _11797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_241_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20910_ _12930_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_222_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21890_ _10022_ _02924_ _02930_ _02932_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_20841_ _01814_ _01828_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24142__A3 _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13969__A2 _07720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23560_ _04286_ _04287_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16954__C _10293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20772_ _12929_ _12261_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22511_ _03428_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23491_ _04134_ _04343_ _04344_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14918__B2 _08564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18109__A1 rbzero.debug_overlay.playerY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_107_i_clk_I clknet_5_31__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25230_ _06013_ _06014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_22442_ _02167_ _03383_ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_147_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14394__A2 _08202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19857__A1 _12260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16970__B _10214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25161_ _05942_ _05944_ _05945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_161_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22373_ _12577_ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24112_ _04876_ _04746_ _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_143_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21324_ _12971_ _02261_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25092_ _05874_ _05858_ _05876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_248_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14490__B _07826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24043_ _04826_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21255_ _12442_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_102_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20206_ _12879_ _12923_ _12978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_224_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21186_ _02119_ _02121_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_224_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15646__A2 _09303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20137_ _12178_ _12908_ _12172_ _12909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25994_ _05208_ _06772_ _06680_ _06659_ _06773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_148_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22916__A1 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20068_ _12833_ _12839_ _12840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24945_ _05702_ _05704_ _05729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__18188__I _11331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24876_ _05439_ _05461_ _05640_ _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26615_ _00525_ clknet_leaf_168_i_clk rbzero.tex_b0\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23827_ _11150_ _04536_ _04659_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18916__I _11825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_198_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14560_ _08200_ _08368_ _08369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26546_ _00456_ clknet_leaf_24_i_clk rbzero.pov.spi_buffer\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_220_Left_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23758_ rbzero.wall_tracer.trackDistY\[-2\] _03056_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17020__A1 _08157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14665__B _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13511_ _07321_ _07322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22709_ _03556_ _03573_ _03574_ _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25094__A1 _05838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14491_ _07509_ _08300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26477_ _00387_ clknet_leaf_211_i_clk rbzero.debug_overlay.playerY\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23689_ _11240_ _03032_ _04537_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_138_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_235_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16230_ _09741_ _09742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25428_ _06207_ _06208_ _06212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_181_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13442_ _06869_ _07142_ _07252_ _07253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_153_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23644__A2 _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19747__I _12518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21655__A1 _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13373_ _07184_ net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16161_ _09690_ _09691_ _09689_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25359_ _06079_ _06080_ _06081_ _06003_ _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_134_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15112_ _08836_ _08897_ _08899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14137__A2 _07938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16092_ _08977_ _09635_ _09639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__17267__I _10571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19920_ _12525_ _12692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15043_ rbzero.spi_registers.spi_counter\[4\] _08836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27029_ _00939_ clknet_leaf_134_i_clk rbzero.tex_g0\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XANTENNA__24602__B _05275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19851_ _12420_ _12274_ _12623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_248_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18802_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] _11734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__20630__A2 _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19782_ _12553_ _12477_ _12482_ _12401_ _12554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16994_ rbzero.pov.ready_buffer\[38\] _10397_ _10400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_207_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18036__B1 _11173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18733_ _11695_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15945_ _09527_ _09528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_222_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22383__A2 _08042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18664_ _11650_ _11656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_222_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15876_ _09462_ _09474_ _09475_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17615_ rbzero.tex_b0\[62\] rbzero.tex_b0\[61\] _10838_ _10840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14827_ rbzero.tex_b1\[28\] _07932_ _08633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_18595_ _11616_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14073__A1 _07848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18339__A1 _07176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17546_ _10800_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14758_ _07603_ _08565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__17011__A1 rbzero.pov.ready_buffer\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14575__B _07808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13709_ _07335_ _07520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17477_ rbzero.tex_b0\[2\] rbzero.tex_b0\[1\] _10760_ _10762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_172_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14689_ _07822_ _08496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_15_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19216_ rbzero.wall_tracer.mapY\[7\] _12056_ _12058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16428_ _08824_ _09887_ _09890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24563__I _05264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19147_ _08155_ _10031_ _11967_ _11991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_172_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16359_ _09838_ _09839_ _09833_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__21646__B2 _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19078_ rbzero.debug_overlay.facingY\[-4\] _10062_ _11922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18029_ _11172_ _11173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21040_ _02010_ _02023_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_165_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16949__C _10293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22991_ _01388_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_33_i_clk_I clknet_5_22__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24730_ net94 _05271_ _05283_ _05514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_21942_ rbzero.wall_tracer.rcp_fsm.o_data\[-11\] _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__20385__A1 _12235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24661_ _05362_ _05254_ _05445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21873_ _02904_ _10087_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17640__I _10857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26400_ _00310_ clknet_leaf_248_i_clk rbzero.spi_registers.buf_texadd2\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23612_ _04396_ _04428_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20824_ _01810_ _01912_ _01913_ _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_27380_ _01285_ clknet_leaf_104_i_clk rbzero.wall_tracer.trackDistY\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__22258__I _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24592_ _05334_ _05295_ _05376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21162__I _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26331_ _00241_ clknet_leaf_234_i_clk rbzero.spi_registers.buf_mapdyw\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20755_ _12835_ _01845_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_23543_ _04320_ _04334_ _04395_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23474_ _03862_ _04327_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26262_ _00172_ clknet_leaf_13_i_clk rbzero.spi_registers.texadd3\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20686_ _01777_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25213_ _05808_ net48 _05997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__21637__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22425_ _03346_ _03368_ _03347_ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26193_ _00103_ clknet_leaf_214_i_clk rbzero.spi_registers.texadd0\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25144_ _05918_ _05927_ _05928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_149_Right_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22356_ _03304_ _03305_ _03252_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14119__A2 _07629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21307_ _02376_ _02393_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25075_ _05836_ _05856_ _05858_ _05859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xclkbuf_leaf_4_i_clk clknet_5_4__leaf_i_clk clknet_leaf_4_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22287_ _03249_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_213_i_clk clknet_5_6__leaf_i_clk clknet_leaf_213_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_206_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24026_ rbzero.wall_tracer.rcp_fsm.operand\[10\] _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__24422__B _05205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17069__A1 _10455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21238_ _02323_ _02324_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21169_ _02000_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__25000__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25977_ _06751_ _06754_ _06755_ _06756_ _06757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_13991_ _07437_ _07801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_228_i_clk clknet_5_2__leaf_i_clk clknet_leaf_228_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_204_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15335__I _08877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15730_ rbzero.spi_registers.buf_texadd2\[22\] _09364_ _09367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24928_ _05671_ _05673_ _05707_ _05712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__20376__A1 _12398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15661_ _09302_ _09315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_241_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_24859_ _05642_ _05643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_83_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_237_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_237_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17400_ _06897_ _10705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_240_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14612_ _08416_ _08417_ _08419_ _08211_ _07604_ _08420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xclkbuf_5_31__f_i_clk clknet_3_7_0_i_clk clknet_5_31__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_212_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18380_ rbzero.tex_g1\[11\] rbzero.tex_g1\[10\] _11491_ _11494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15592_ rbzero.spi_registers.buf_texadd1\[11\] _09259_ _09264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17331_ rbzero.pov.spi_buffer\[37\] _10650_ _10646_ _10654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14543_ _08335_ _08350_ _08351_ _08352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26529_ _00439_ clknet_leaf_38_i_clk rbzero.pov.spi_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17262_ _10542_ _10602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_12_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14474_ rbzero.tex_g0\[37\] _08279_ _08282_ _08283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_165_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19001_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _11872_ _11875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__19477__I rbzero.wall_tracer.side vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16213_ _09728_ _09729_ _09723_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__21628__A1 _10455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13425_ _07235_ _07236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_107_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17193_ _10549_ _10545_ _10550_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16144_ rbzero.spi_registers.buf_texadd1\[1\] _09672_ _09679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_114_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13739__B _07549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13356_ _07164_ _07161_ _07159_ _07167_ gpout2.clk_div\[1\] _07154_ _07168_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_52_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16075_ _09623_ _09625_ _09626_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__24042__A2 _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13869__A1 rbzero.debug_overlay.playerX\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13287_ _07100_ _07101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22053__A1 _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19903_ _12674_ _12675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15026_ _08818_ rbzero.spi_registers.ss_buffer\[0\] _08820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_227_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16807__A1 rbzero.debug_overlay.playerX\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21800__A1 _09982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19834_ _12537_ _12605_ _12606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19765_ _12393_ _12535_ _12536_ _12537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_208_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16977_ _10382_ _10384_ _10386_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 i_gpout0_sel[1] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15928_ rbzero.spi_registers.spi_buffer\[1\] _09515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18716_ _11685_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19696_ _12369_ _12465_ _12466_ _12467_ _12468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_160_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18647_ rbzero.tex_r0\[62\] rbzero.tex_r0\[61\] _11644_ _11646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15859_ _09444_ _09458_ _09463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14046__A1 rbzero.tex_r1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22108__A2 _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17783__A2 rbzero.pov.ready_buffer\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18578_ _11606_ _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17529_ _10780_ _10791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20540_ _12968_ _01377_ _01631_ _12431_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23608__A2 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20471_ _01481_ _01563_ _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21619__B2 _10036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16804__I _09139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22210_ _03182_ _03183_ _03185_ _03180_ rbzero.wall_tracer.rcp_fsm.i_data\[7\] _03186_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_172_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14752__C _08334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23190_ _03931_ _04045_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_41_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22141_ _03119_ _03129_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22419__I0 _08061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_22072_ _03069_ _03070_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14521__A2 _07834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25900_ _06650_ _06683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_239_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21023_ _02111_ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22595__A2 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26880_ _00790_ clknet_leaf_161_i_clk rbzero.tex_r0\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__19460__A2 _12227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17471__A1 _07052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25831_ _05995_ _06614_ _06615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_227_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25762_ _06515_ _06544_ _06546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20358__A1 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22974_ _03805_ _03831_ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_24713_ _05491_ _05496_ _05497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_223_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_21925_ _02920_ _02952_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25693_ _06439_ _06440_ _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14037__A1 _07842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27432_ _01337_ clknet_leaf_78_i_clk rbzero.wall_tracer.rcp_fsm.operand\[8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_195_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24644_ _05417_ _05426_ _05427_ _05428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_21856_ _10484_ _02879_ _02891_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_218_Right_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_27363_ _01268_ clknet_leaf_102_i_clk rbzero.wall_tracer.trackDistX\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20807_ _01788_ _01896_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24575_ _05357_ _05358_ _05359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21787_ _10448_ _02836_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_61_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26314_ _00224_ clknet_leaf_232_i_clk rbzero.spi_registers.buf_vshift\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23526_ _04219_ _04054_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15537__A1 rbzero.spi_registers.buf_texadd0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_232_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20738_ _01814_ _01828_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_147_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_27294_ _01199_ clknet_leaf_210_i_clk rbzero.row_render.size\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_232_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26245_ _00155_ clknet_leaf_20_i_clk rbzero.spi_registers.texadd2\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_247_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23457_ _04202_ _04205_ _04310_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_20669_ _01634_ _01635_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13210_ _07019_ _07023_ _07024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_208_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__22283__A1 _11175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22408_ _03320_ _10200_ _03352_ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26176_ _00086_ clknet_leaf_228_i_clk rbzero.color_floor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14190_ _06888_ _07974_ _08000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23388_ _03491_ _04129_ _04242_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_152_i_clk clknet_5_11__leaf_i_clk clknet_leaf_152_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25127_ _05877_ _05905_ _05911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13141_ _06910_ _06952_ _06954_ _06955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22339_ rbzero.wall_tracer.trackDistY\[7\] _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__25221__A1 _05869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_210_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13072_ _06884_ _06887_ _06888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_76_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25058_ net79 _05385_ _05840_ _05842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_20_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23783__A1 rbzero.wall_tracer.trackDistY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16900_ _10309_ _10320_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_218_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24009_ _04794_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_218_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17880_ _11005_ _11022_ _11023_ _11024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_245_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16831_ _10209_ _10260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14276__A1 _08084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22338__A2 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14276__B2 _08085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19550_ _12321_ _12322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_73_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16762_ _10193_ _10180_ _10199_ _10187_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_13974_ _07720_ _07139_ _07784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18501_ _11562_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15713_ _09351_ _09354_ _09348_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19481_ rbzero.wall_tracer.size\[3\] _12247_ _12251_ _12252_ _12253_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_220_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16693_ _10015_ _10136_ _10137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_17_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17765__A2 rbzero.pov.ready_buffer\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18432_ rbzero.tex_g1\[33\] rbzero.tex_g1\[32\] _11523_ _11524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_107_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15644_ _09204_ _09302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13741__C _07551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14579__A2 _07816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23838__A2 _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18363_ _11484_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_186_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15575_ _09249_ _09250_ _09242_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13313__I _06981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_105_i_clk clknet_5_30__leaf_i_clk clknet_leaf_105_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17314_ _10618_ _10641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14526_ _07549_ _08335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18294_ _07180_ _11433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13539__B1 _07329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17245_ _10587_ _10583_ _10589_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14457_ rbzero.tex_g0\[9\] _07584_ _08266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16624__I _09972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25460__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13408_ gpout0.vpos\[6\] _07219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__20146__I _12917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17176_ _10520_ _10536_ _10518_ _10515_ _10537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14388_ rbzero.color_floor\[2\] _08197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16127_ _09011_ _09657_ _09665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13339_ net41 _07146_ _07152_ net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_84_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24062__B _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22026__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16058_ _09428_ _09614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15009_ _08808_ _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_206_i_clk_I clknet_5_18__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19817_ _12381_ _12262_ _12282_ _12521_ _12589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_127_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25515__A2 _06045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19748_ _12519_ _12520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_155_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19679_ _12355_ _12357_ _12360_ _12352_ _12451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_140_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21710_ _02769_ _02733_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22690_ _11238_ _12499_ _03557_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__20760__A1 _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23829__A2 _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21641_ _02714_ _02716_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_220_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24360_ _04905_ _04910_ _05052_ _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_21572_ _02552_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26008__I _06737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20512__A1 _12685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14990__A2 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_214_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_173_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20523_ _01614_ _01615_ _12906_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23311_ _03931_ _04165_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24291_ _05011_ _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_28_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26030_ _06771_ _06780_ _06804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20454_ _01372_ _01545_ _01547_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_23242_ _12961_ _03714_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14742__A2 _08526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23173_ _03933_ _03956_ _04028_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20385_ _12235_ _01478_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19681__A2 _12447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22124_ _03114_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_84_i_clk clknet_5_28__leaf_i_clk clknet_leaf_84_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_11_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22055_ _03030_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_203_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26932_ _00842_ clknet_leaf_174_i_clk rbzero.tex_r1\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_21006_ rbzero.wall_tracer.stepDistY\[9\] _01838_ _01839_ _02094_ _02095_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_227_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26863_ _00773_ clknet_leaf_176_i_clk rbzero.tex_r0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14258__A1 _07720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25814_ _05993_ _06596_ _06597_ _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xclkbuf_leaf_99_i_clk clknet_5_27__leaf_i_clk clknet_leaf_99_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26794_ _00704_ clknet_leaf_194_i_clk rbzero.tex_g1\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__19197__A1 _09895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25745_ _06031_ _05970_ _06452_ _06385_ _06529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__16709__I _09988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22957_ _02502_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13481__A2 rbzero.spi_registers.vshift\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15613__I _09254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17747__A2 rbzero.pov.ready_buffer\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14657__C _07464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21908_ _11064_ _02949_ _10125_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20751__A1 _12173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25676_ _06448_ _06458_ _06459_ _06460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_193_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13690_ _07488_ _07501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_85_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22888_ _03640_ _03745_ _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_22_i_clk clknet_5_5__leaf_i_clk clknet_leaf_22_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_27415_ _01320_ clknet_leaf_85_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_210_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24627_ _05410_ _05411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_214_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21839_ _02883_ _02884_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_195_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27346_ _01251_ clknet_leaf_94_i_clk rbzero.wall_tracer.w\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15360_ rbzero.spi_registers.buf_mapdyw\[0\] _09092_ _09093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24558_ _05326_ _05341_ _05342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18172__A2 _11256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_2_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14311_ rbzero.debug_overlay.vplaneX\[10\] _08121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_230_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23509_ _04301_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16444__I _08110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_155_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15291_ _08987_ _09042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_37_i_clk clknet_5_5__leaf_i_clk clknet_leaf_37_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_27277_ _01182_ clknet_leaf_205_i_clk rbzero.wall_tracer.texu\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_124_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24489_ _05272_ _05273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17030_ _10407_ _10424_ _10426_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_22_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22256__A1 rbzero.wall_tracer.visualWallDist\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26228_ _00138_ clknet_leaf_0_i_clk rbzero.spi_registers.texadd1\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14242_ _08029_ _08036_ _08040_ _08041_ _08051_ _08052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__14733__A2 _08233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_170_Left_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26159_ _00069_ clknet_leaf_185_i_clk rbzero.mapdyw\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14173_ _06862_ _07981_ _07982_ _07983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_22_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold45_I i_gpout0_sel[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13124_ rbzero.spi_registers.texadd0\[11\] _06911_ _06938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18981_ _11863_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_245_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17275__I _10611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17932_ _08085_ _11075_ _11016_ _11076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_13055_ _06871_ _06872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19424__A2 _12006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17863_ _11006_ _11007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_109_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19602_ rbzero.wall_tracer.stepDistX\[-3\] _12374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_16814_ _10243_ _10239_ _10245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_233_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17794_ _10959_ rbzero.pov.ready_buffer\[55\] _10960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19533_ _12300_ _12304_ _12305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16745_ _10168_ _10184_ _10185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13957_ _07735_ _07766_ _07767_ _07768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_89_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19464_ _12235_ _12236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_122_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16676_ _09897_ _10121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13888_ rbzero.debug_overlay.playerX\[-3\] _07699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_201_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15627_ _09289_ _09290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18415_ rbzero.tex_g1\[26\] rbzero.tex_g1\[25\] _11512_ _11514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_19395_ _12166_ _12167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_189_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24484__A2 _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24057__B _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18346_ _07179_ _11471_ _11472_ _11473_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_15558_ _09236_ _09237_ _09229_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14509_ rbzero.tex_g0\[53\] _08317_ _08318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_155_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18277_ _11402_ _11417_ _11418_ _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15489_ rbzero.spi_registers.buf_texadd0\[9\] _09178_ _09187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_226_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17228_ _10564_ _10577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14724__A2 _08528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19112__A1 _08151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17159_ _10513_ _10523_ rbzero.pov.spi_counter\[1\] _10525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_130_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20170_ _12240_ _12672_ _12941_ _12942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14488__A1 rbzero.tex_g0\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17185__I _10543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19415__A2 rbzero.wall_tracer.rayAddendY\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_236_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_236_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23860_ _02980_ _04686_ _04688_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_22811_ _12817_ _03669_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_0_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23791_ _04627_ rbzero.wall_tracer.stepDistY\[3\] _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16529__I _09934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13463__A2 rbzero.spi_registers.vshift\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25530_ _06268_ _06313_ _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22742_ _03548_ _03602_ _03603_ _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_189_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_175_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_175_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25461_ _06236_ _06239_ _06242_ _06244_ _06245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_192_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22673_ _11201_ _03539_ _03542_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_48_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27200_ _01105_ clknet_leaf_74_i_clk rbzero.wall_tracer.size_full\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_192_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24412_ _05190_ _05195_ _05196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_21624_ _10086_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22486__A1 rbzero.wall_tracer.size\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25392_ _06122_ _06128_ _06176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_176_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21170__I _12522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13888__I rbzero.debug_overlay.playerX\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27131_ _01041_ clknet_leaf_224_i_clk gpout0.clk_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24343_ _05126_ _05053_ _05127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21555_ _02620_ _02639_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__26566__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20506_ _01597_ _01598_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_145_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27062_ _00972_ clknet_leaf_148_i_clk rbzero.tex_b1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24274_ _05057_ _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15912__A1 _08957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21486_ _02446_ _02566_ _02570_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_200_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20249__B1 _13017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26013_ _06721_ _06724_ _06749_ _06790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20437_ _01527_ _01529_ _01530_ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_205_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23225_ _12949_ _04080_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_200_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20514__I _12917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23156_ _04010_ _04011_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21461__A2 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20368_ _01458_ _01461_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_56_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_227_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22107_ _03090_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23087_ _03823_ _03826_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_8_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14512__I _07493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20299_ _01384_ _01387_ _01393_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_246_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13151__A1 _06962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22038_ rbzero.wall_tracer.stepDistY\[-5\] _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26915_ _00825_ clknet_leaf_135_i_clk rbzero.tex_r1\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__22410__A1 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26846_ _00756_ clknet_leaf_193_i_clk rbzero.tex_r0\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14860_ rbzero.tex_b1\[1\] _08241_ _07861_ _08666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_240_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_240_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_6_0_i_clk_I clknet_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_81_i_clk_I clknet_5_28__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13811_ _07615_ _07621_ _07622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_230_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16439__I _09896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14791_ _07601_ _08596_ _08597_ _08598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_26777_ _00687_ clknet_leaf_122_i_clk rbzero.tex_g1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_98_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23989_ _04779_ _08814_ _04780_ _11473_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_230_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16530_ _08111_ _08098_ _09983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25728_ _06509_ _06511_ _06512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13742_ _07542_ _07552_ _07553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_27_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16461_ _09895_ _09898_ _09919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_27_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25659_ _06399_ _06411_ _06443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_183_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13673_ _07483_ _07484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__18654__I _11649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18200_ _11109_ _11344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_182_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15412_ rbzero.spi_registers.buf_sky\[5\] _09131_ _09132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19180_ _11340_ _12008_ _12023_ _12024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16392_ rbzero.spi_registers.buf_texadd3\[16\] _09863_ _09864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_100_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18145__A2 _11287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13798__I _07608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18131_ rbzero.debug_overlay.playerY\[4\] _11250_ _11275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_15343_ rbzero.spi_registers.buf_mapdy\[3\] _09080_ _09081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_27329_ _01234_ clknet_leaf_201_i_clk rbzero.row_render.wall\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16156__A1 _08926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18062_ _11205_ _11206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_124_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14706__A2 _08506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15274_ rbzero.map_overlay.i_otherx\[4\] _09027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__26523__D _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17013_ _10411_ _10413_ _10414_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14225_ _08015_ _08034_ _08035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_34_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14156_ _07425_ _07966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_186_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23729__A1 _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15518__I _09208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13107_ _06920_ _06921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_81_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14087_ rbzero.tex_r1\[39\] _07834_ _07897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18964_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _11851_ _11854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24340__B _05123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17915_ _11044_ _11057_ _11058_ _11059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18895_ rbzero.traced_texa\[6\] _07273_ _11809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_218_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17846_ _10845_ _10992_ _10520_ _10539_ _10993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_234_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21255__I _12442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24154__A1 _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23671__S _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16349__I _09806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14989_ _08789_ _08790_ _08791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17777_ _10944_ rbzero.pov.ready_buffer\[49\] _10949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18908__A1 rbzero.traced_texa\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23901__A1 _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19516_ _12244_ _12288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_191_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16728_ _10168_ _10169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__20715__A1 _12426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19447_ _12168_ _12215_ _12218_ _12219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_187_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16659_ _09953_ _10096_ _10102_ _10104_ _10105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25654__A1 _05889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19378_ _12154_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18136__A2 _11279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_211_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18329_ _10988_ _07202_ _11459_ _11460_ _11461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_211_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19884__A2 _12160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25397__I _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21340_ _02425_ _02426_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__26433__D _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21271_ _02215_ _02216_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_8_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16812__I _07677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20222_ _12560_ _12273_ _12994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23010_ _02404_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21443__A2 _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25709__A2 _06051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20153_ _12877_ _12924_ _12925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_168_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24393__A1 _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20084_ _12823_ _12824_ _12855_ _12856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24961_ _05734_ _05735_ _05721_ _05745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__16870__A2 _10252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_103_i_clk_I clknet_5_30__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26700_ _00610_ clknet_leaf_63_i_clk rbzero.pov.ready_buffer\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23912_ _04718_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24892_ _05672_ _05674_ _05675_ _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_222_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16622__A2 _09977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26631_ _00541_ clknet_leaf_161_i_clk rbzero.tex_b0\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_169_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23843_ _11143_ _04536_ _04673_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_212_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26562_ _00472_ clknet_leaf_63_i_clk rbzero.pov.spi_buffer\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_240_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23774_ _11167_ rbzero.wall_tracer.stepDistY\[1\] _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20986_ _01966_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_196_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25513_ _06277_ _06292_ _06296_ _06297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_22725_ rbzero.wall_tracer.trackDistX\[-2\] _03522_ _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26493_ _00403_ clknet_leaf_55_i_clk rbzero.debug_overlay.facingY\[-7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_24_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16386__A1 rbzero.spi_registers.spi_buffer\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25444_ _06221_ _06225_ _06227_ _06228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_165_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22656_ _02733_ _03527_ _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16138__A1 _08843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21607_ gpout0.clk_div\[0\] _11826_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25375_ _06108_ _06114_ _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14507__I _07501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22587_ _03474_ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__24425__B _05111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27114_ _01024_ clknet_leaf_141_i_clk rbzero.tex_b1\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_106_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24326_ _05043_ _05107_ _05108_ _05109_ _05110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA_clkbuf_leaf_28_i_clk_I clknet_5_20__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21538_ _02484_ _02621_ _02622_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_105_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_248_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17818__I _09035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_229_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27045_ _00955_ clknet_leaf_160_i_clk rbzero.tex_g0\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24257_ _04895_ _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21469_ _02539_ _02554_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_133_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14010_ rbzero.tex_r1\[25\] _07818_ _07819_ _07820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23208_ _02633_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24188_ _04840_ _04921_ _04972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22660__S _11400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15338__I _08883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23139_ _03908_ _03995_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_242_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_248_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_235_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18850__A3 _11772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24384__A1 _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15961_ _09525_ _09527_ _09540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_207_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14872__A1 _07889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17700_ _10897_ rbzero.pov.ready_buffer\[23\] _10898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14912_ rbzero.tex_b1\[61\] _07592_ _08717_ _08718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_234_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15892_ _08928_ _09477_ _09488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18680_ rbzero.tex_r1\[12\] rbzero.tex_r1\[11\] _11661_ _11665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_216_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20945__A1 rbzero.traced_texVinit\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21993__I0 rbzero.wall_tracer.rcp_fsm.o_data\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20945__B2 _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14843_ rbzero.tex_b1\[21\] _07633_ _08649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17631_ _10844_ _10852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26829_ _00739_ clknet_leaf_177_i_clk rbzero.tex_g1\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_216_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17562_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _10807_ _10810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14774_ _07624_ _08559_ _08566_ _08572_ _08580_ _08581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_98_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16513_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.wall_tracer.rayAddendY\[-2\] _09959_
+ _09967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_19301_ rbzero.tex_b1\[30\] rbzero.tex_b1\[29\] _12109_ _12111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13725_ rbzero.tex_r0\[34\] _07535_ _07337_ _07536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_168_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17493_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _10770_ _10771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__18384__I _11480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24439__A2 _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16444_ _08110_ _09902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19232_ _11478_ _12071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13656_ _07458_ _07466_ _07467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_67_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23111__A2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19163_ _12006_ _12007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16129__A1 rbzero.spi_registers.buf_texadd0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14417__I _07511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16375_ _09815_ _09851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__21122__A1 rbzero.wall_tracer.stepDistY\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13587_ _07364_ _07385_ _07398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18114_ rbzero.debug_overlay.playerY\[2\] _11255_ _11256_ _10358_ _11257_ _11258_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_15326_ _09067_ _09068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19094_ _11922_ _11936_ _11937_ _11938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18045_ _11160_ _11162_ _11188_ _11189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15257_ rbzero.pov.sclk_buffer\[1\] _09015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_152_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14208_ rbzero.debug_overlay.playerY\[0\] _08018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15188_ rbzero.spi_registers.spi_buffer\[9\] _08962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_130_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14139_ rbzero.tex_r1\[60\] _07940_ _07948_ _07949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_130_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25166__B _05949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19996_ _12759_ _12767_ _12768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_226_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24375__A1 _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18947_ rbzero.tex_g0\[12\] rbzero.tex_g0\[11\] _11840_ _11844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_225_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14863__B2 _08522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18878_ rbzero.traced_texa\[2\] rbzero.texV\[2\] _11794_ _11796_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_33_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17829_ _09035_ _10982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14615__A1 _07848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_222_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20840_ _01915_ _01929_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24296__I _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18294__I _07180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20771_ _01749_ _01750_ _01861_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_119_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15711__I _09352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22510_ rbzero.wall_tracer.texu\[0\] _03423_ _03424_ _08360_ _03428_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23490_ _04023_ _04235_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_162_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18109__A2 _11252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22441_ _03341_ _07704_ _03382_ _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19857__A2 _12496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13231__I _07044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25160_ _05871_ _05908_ _05943_ _05944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_190_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22544__I _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22372_ _03318_ _03319_ _03079_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24111_ _04749_ _04864_ _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__17638__I rbzero.pov.spi_done vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21323_ _02409_ _02250_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25091_ _05874_ _05858_ _05875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24042_ _04809_ _04825_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21254_ _12439_ _12440_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22613__A1 _12163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20064__I _12835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20205_ _12962_ _12976_ _12977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_21185_ _02270_ _02272_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_224_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24366__A1 _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20136_ _10996_ _11032_ _12908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25993_ _06771_ _06772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_148_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14854__A1 rbzero.tex_b1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_20067_ _12667_ _12837_ _12838_ _12839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_24944_ _05330_ _05728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__19793__A1 _12556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24875_ _05658_ _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26614_ _00524_ clknet_leaf_163_i_clk rbzero.tex_b0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23826_ _04242_ _04658_ _04528_ _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19545__A1 rbzero.wall_tracer.visualWallDist\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18348__A2 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14082__A2 _07855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_198_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26545_ _00455_ clknet_leaf_24_i_clk rbzero.pov.spi_buffer\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23757_ _11178_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_178_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_20969_ _01943_ _01960_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13510_ _07260_ _07319_ _07320_ _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_22708_ _03560_ _01892_ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_14490_ rbzero.tex_g0\[44\] _08298_ _07826_ _08299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__14909__A2 _08568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26476_ _00386_ clknet_leaf_208_i_clk rbzero.debug_overlay.playerY\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_23688_ rbzero.wall_tracer.trackDistY\[-11\] _03032_ _04537_ _04538_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_165_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_235_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25427_ _06207_ _06208_ _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13441_ _07080_ _07251_ _06868_ _07252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_22639_ rbzero.wall_tracer.w\[1\] _03508_ _03493_ _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14237__I _08046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16160_ _09542_ _09687_ _09691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25358_ _05996_ _05973_ _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__21655__A2 _08377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13372_ _07169_ _07183_ net15 _07184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__26043__A1 _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15111_ _08836_ _08897_ _08898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24309_ _04932_ _05091_ _05092_ _05093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_134_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16091_ rbzero.spi_registers.buf_texadd0\[13\] _09633_ _09638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25289_ _05530_ _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_146_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15042_ _08825_ _08832_ _08834_ _08835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_27028_ _00938_ clknet_leaf_136_i_clk rbzero.tex_g0\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XPHY_EDGE_ROW_2_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_39_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_19850_ _12470_ _12560_ _12622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_112_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24357__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18801_ _11733_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19781_ _12476_ _12553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16993_ _08088_ _10393_ _10399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14845__A1 _07814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17283__I _10543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22907__A2 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18732_ rbzero.tex_r1\[34\] rbzero.tex_r1\[33\] _11693_ _11695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15944_ _09437_ _08845_ _09527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_235_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24109__A1 _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15875_ _08942_ _09460_ _09475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18663_ _11655_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17614_ _10839_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14826_ rbzero.tex_b1\[30\] _08631_ _08280_ _08632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19431__C _12202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18594_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _11613_ _11616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_188_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_48_Left_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13760__B _07570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14757_ _07636_ _08564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17545_ rbzero.tex_b0\[32\] rbzero.tex_b0\[31\] _10796_ _10800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13820__A2 _07629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13708_ rbzero.tex_r0\[63\] _07518_ _07519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17476_ _10761_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14688_ rbzero.tex_b0\[54\] _08494_ _08495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19215_ rbzero.wall_tracer.mapY\[7\] _12056_ _12057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_172_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16427_ _08828_ _09886_ _09889_ _08888_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_13639_ rbzero.row_render.texu\[2\] _07450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16770__A1 rbzero.pov.ready_buffer\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19146_ _11925_ _11969_ _11990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_15_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16358_ _08944_ _09831_ _09839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21646__A2 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21110__A4 _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15309_ _09054_ _09055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16362__I _09819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19077_ _08153_ rbzero.wall_tracer.rayAddendY\[5\] _11921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16522__A1 _09974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16289_ rbzero.spi_registers.buf_texadd2\[14\] _09780_ _09787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18028_ rbzero.wall_tracer.trackDistX\[-2\] _11172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_238_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_227_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21708__I _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25545__B1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19979_ _12750_ _12676_ _12723_ _12681_ _12751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_158_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22990_ _03846_ _03709_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20909__A1 _12211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21941_ _02979_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__20385__A2 _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13226__I _07039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24660_ _05284_ _05442_ _05443_ _05444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_143_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21872_ _02912_ _02915_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_143_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14064__A2 _07872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23611_ _04461_ _04460_ _04462_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__17142__B _10508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20823_ _01812_ _01852_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20137__A2 _12908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24591_ _05304_ _05374_ _05375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_148_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15441__I _08883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26330_ _00240_ clknet_leaf_234_i_clk rbzero.spi_registers.buf_mapdyw\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23542_ _04318_ _04336_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20754_ rbzero.wall_tracer.stepDistX\[7\] _12206_ _01844_ _01845_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_64_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26261_ _00171_ clknet_leaf_10_i_clk rbzero.spi_registers.texadd3\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_174_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23473_ _01969_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14057__I _07501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16761__A1 rbzero.pov.ready_buffer\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20685_ rbzero.traced_texVinit\[3\] _01553_ _01776_ _01662_ _01777_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25212_ _05372_ _05996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_162_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22424_ _03364_ _03367_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22834__A1 _12684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26192_ _00102_ clknet_leaf_239_i_clk rbzero.spi_registers.texadd0\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25143_ _05926_ _05927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22355_ _11296_ _03249_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13327__A1 _06879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21306_ _02382_ _02392_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_20_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25074_ _05792_ _05797_ _05857_ _05858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_22286_ _11138_ _03248_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13878__A2 _07685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24025_ _04772_ _04808_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__17069__A2 _10432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21237_ _02318_ _02319_ _02322_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_130_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21168_ _12210_ _13012_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__25000__A2 _05308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20119_ _12421_ _12258_ _12891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25976_ _06742_ _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21099_ _02074_ _02082_ _02186_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_13990_ _07776_ _07799_ _07767_ _07800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_205_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24927_ _05710_ _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__25839__A1 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15660_ _09312_ _09313_ _09314_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24858_ _05640_ _05641_ _05642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_213_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14055__A2 _07822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_237_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14611_ rbzero.tex_g1\[5\] _07832_ _08418_ _08419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_237_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23809_ _04639_ _04642_ _04643_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15591_ rbzero.spi_registers.texadd1\[11\] _09255_ _09263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24789_ _05572_ _05573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17330_ _10618_ _10653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_185_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14542_ rbzero.tex_g0\[58\] _08342_ _08351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26528_ _00438_ clknet_leaf_38_i_clk rbzero.pov.spi_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__26084__C _11825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17261_ rbzero.pov.spi_buffer\[19\] _10601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_138_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14473_ rbzero.tex_g0\[36\] _07909_ _08282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_26459_ _00369_ clknet_leaf_207_i_clk rbzero.debug_overlay.playerX\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_193_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14358__A3 _08167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16752__A1 _10168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16212_ _09000_ _09721_ _09729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19000_ _11874_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13424_ _07234_ _07235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_64_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22184__I _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22825__A1 _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17192_ rbzero.pov.spi_buffer\[2\] _10547_ _10174_ _10550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16143_ _09673_ _09677_ _09678_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_114_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13355_ _07166_ _07167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_107_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16074_ _09614_ _09626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13286_ _06878_ _07100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19707__B _12442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19902_ _12427_ _12674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__24332__C _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15025_ _08819_ _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_209_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19833_ _12543_ _12602_ _12604_ _12605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__20432__I _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14818__A1 _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19764_ _12456_ _12534_ _12536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_236_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16976_ _10385_ _10386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23743__I _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18715_ rbzero.tex_r1\[27\] rbzero.tex_r1\[26\] _11682_ _11685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput6 net95 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15927_ rbzero.spi_registers.buf_othery\[1\] _09510_ _09514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19695_ _12437_ _12443_ _12467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_160_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_56_Left_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18646_ _11645_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15858_ _09139_ _09462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__19509__A1 _08181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14046__A2 _07855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14809_ rbzero.row_render.side _07446_ _08616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__20119__A2 _12258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18577_ rbzero.tex_r0\[32\] rbzero.tex_r0\[31\] _11602_ _11606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15261__I _08987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15789_ _09408_ _09410_ _09406_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17528_ _10790_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__25058__A2 _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_202_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17459_ rbzero.pov.spi_buffer\[70\] _10743_ _10740_ _10749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21619__A2 _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22094__I _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20470_ _01487_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_171_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_Left_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__17188__I _10546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19129_ _11959_ _11971_ _11972_ _11973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_125_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22140_ rbzero.wall_tracer.rcp_fsm.i_data\[-6\] _03126_ _03128_ _03129_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22071_ _03038_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_199_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21438__I _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21022_ rbzero.wall_tracer.visualWallDist\[9\] _12228_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__23792__A2 rbzero.wall_tracer.stepDistY\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14809__A1 rbzero.row_render.side vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15436__I _09111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25830_ _06548_ _06607_ _06613_ _06614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_145_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15482__A1 _06962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Left_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_199_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25761_ _06515_ _06544_ _06545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22973_ _03808_ _03830_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__18747__I _11692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17651__I _10857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24712_ _05492_ _05493_ _05494_ _05495_ _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_21924_ _02921_ _02952_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25692_ _06442_ _06474_ _06475_ _06476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_241_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21173__I _12587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27431_ _01336_ clknet_leaf_73_i_clk rbzero.wall_tracer.rcp_fsm.operand\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_182_Right_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24643_ _05424_ _05425_ _05427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_219_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_178_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21307__A1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16267__I _09747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21855_ _10481_ _11072_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_195_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27362_ _01267_ clknet_leaf_102_i_clk rbzero.wall_tracer.trackDistX\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20806_ _01888_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_24574_ _05349_ _05355_ _05358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__21858__A2 _09921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21786_ _08127_ _08129_ _08139_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_148_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26313_ _00223_ clknet_leaf_235_i_clk rbzero.spi_registers.buf_vshift\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23525_ _03979_ _04052_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20737_ _01822_ _01827_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_136_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27293_ _01198_ clknet_leaf_211_i_clk rbzero.row_render.size\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16734__A1 _08182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_232_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20530__A2 _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_232_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Left_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26244_ _00154_ clknet_leaf_21_i_clk rbzero.spi_registers.texadd2\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_98_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23456_ _04199_ _03965_ _04203_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_18_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20668_ _01758_ _01759_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_208_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17098__I _10477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22407_ _03320_ _08062_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26175_ _00085_ clknet_leaf_233_i_clk rbzero.color_floor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__22283__A2 _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23387_ _03898_ _04241_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20599_ _12424_ _12587_ _01593_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__20294__A1 _12660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25126_ _05909_ _05869_ _05910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_13140_ rbzero.spi_registers.texadd0\[8\] _06953_ _06954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22338_ _03274_ _03289_ _03291_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20833__A3 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_210_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25057_ _05840_ _05639_ _05841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13071_ _06885_ _06886_ _06887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_76_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19287__I0 rbzero.tex_b1\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22269_ _03225_ _03233_ _03234_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_76_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20046__A1 _12816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24008_ rbzero.wall_tracer.rcp_fsm.operand\[10\] _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__20252__I _13023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23783__A2 rbzero.wall_tracer.stepDistY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_92_Left_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16830_ _10258_ _10212_ _10259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14276__A2 _08035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_151_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13973_ _07203_ _06875_ _06865_ _07226_ _07783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_16761_ rbzero.pov.ready_buffer\[62\] _10183_ _10179_ _10198_ _10199_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_25959_ _06667_ _06675_ _06740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18500_ rbzero.tex_g1\[63\] rbzero.tex_g1\[62\] _11559_ _11562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15712_ rbzero.spi_registers.buf_texadd2\[17\] _09353_ _09354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19480_ _12165_ _12252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16692_ _10132_ _10112_ _10134_ _10136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_198_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18431_ _11522_ _11523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_107_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15643_ _09299_ _09300_ _09301_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15574_ rbzero.spi_registers.buf_texadd1\[7\] _09245_ _09250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18362_ rbzero.tex_g1\[3\] rbzero.tex_g1\[2\] _11481_ _11484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_185_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_201_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18175__B1 rbzero.map_rom.i_row\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17313_ rbzero.pov.spi_buffer\[32\] _10640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14525_ _07541_ _08334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_127_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18293_ _07790_ _11432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14853__C _08346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14456_ rbzero.tex_g0\[8\] _07816_ _08265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17244_ rbzero.pov.spi_buffer\[15\] _10580_ _10588_ _10589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13407_ _07216_ _07217_ _07218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_153_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17175_ _10532_ rbzero.pov.spi_counter\[4\] _10535_ _10536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__17525__I0 rbzero.tex_b0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14387_ _07186_ _08194_ _08196_ net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_40_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_76_i_clk_I clknet_5_30__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16126_ rbzero.spi_registers.buf_texadd0\[22\] _09655_ _09664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13338_ _07064_ _07147_ _07149_ _07151_ _06887_ _07152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_40_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16057_ _09525_ _09612_ _09613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13269_ _06930_ _06984_ _06986_ _07083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15700__A2 _09338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20037__A1 _12780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15008_ _08807_ rbzero.wall_tracer.rcp_fsm.state\[3\] _08808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_209_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23774__A2 rbzero.wall_tracer.stepDistY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20588__A2 _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21785__A1 _10036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19816_ _12302_ _12587_ _12588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23473__I _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19747_ _12518_ _12519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16959_ _10370_ _10371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_212_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19678_ _12338_ _12340_ _12343_ _12334_ _12450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_211_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18629_ rbzero.tex_r0\[54\] rbzero.tex_r0\[53\] _11634_ _11636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_177_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_29__f_i_clk_I clknet_3_7_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_i_clk clknet_5_1__leaf_i_clk clknet_leaf_3_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21640_ _09904_ _09971_ _02715_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_212_i_clk clknet_5_7__leaf_i_clk clknet_leaf_212_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18166__B1 _11306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21721__I _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21571_ _02647_ _02655_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__16716__A1 _10151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20512__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14990__A3 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23310_ _04154_ _04164_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20522_ rbzero.wall_tracer.size_full\[5\] _01527_ _12182_ _01615_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_214_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_173_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24290_ _05058_ _05073_ _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_133_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25451__A2 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23241_ _03940_ _03941_ _04096_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_138_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_227_i_clk clknet_5_2__leaf_i_clk clknet_leaf_227_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20453_ _01374_ _01546_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20276__A1 _12949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13950__A1 gpout0.vpos\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23172_ _03915_ _03932_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20384_ _12260_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__17141__A1 rbzero.pov.ready_buffer\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22123_ _03084_ _03086_ _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_101_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23765__A2 rbzero.wall_tracer.stepDistY\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22054_ _03008_ _03045_ _03059_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26931_ _00841_ clknet_leaf_173_i_clk rbzero.tex_r1\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_100_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21005_ _02090_ _02093_ _01838_ _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_195_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26862_ _00772_ clknet_leaf_179_i_clk rbzero.tex_r0\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14258__A2 _07202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25813_ _05949_ _05990_ _05981_ _06597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26793_ _00703_ clknet_leaf_195_i_clk rbzero.tex_g1\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_242_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25744_ _06439_ _06440_ _06483_ _06528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__24190__A2 _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22956_ _02277_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20200__A1 _12432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21907_ _02939_ _02940_ _02946_ _02948_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_25675_ _06073_ _05969_ _06459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22887_ _03640_ _03745_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_222_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27414_ _01319_ clknet_leaf_85_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24626_ _05205_ _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_167_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_214_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21838_ _02857_ _02871_ _02869_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21631__I _09899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27345_ _01250_ clknet_leaf_94_i_clk rbzero.wall_tracer.w\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24557_ _05339_ _05340_ _05341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__16707__A1 _10072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21769_ _02811_ _02819_ _02820_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16707__B2 _10049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14310_ _08097_ _08101_ _08115_ _08119_ _08120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_23508_ _04262_ _04340_ _04360_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_15290_ rbzero.spi_registers.buf_othery\[1\] _09021_ _09041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27276_ _01181_ clknet_leaf_205_i_clk rbzero.wall_tracer.texu\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24488_ _05269_ _05271_ _05272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_230_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26227_ _00137_ clknet_leaf_0_i_clk rbzero.spi_registers.texadd1\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_22_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14194__A1 _07976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14241_ _08050_ _08051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_22_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23439_ _04292_ _04180_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13289__C _07102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26158_ _00068_ clknet_leaf_188_i_clk rbzero.mapdxw\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14172_ _07144_ _07981_ _07982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17132__A1 rbzero.pov.ready_buffer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25109_ _05287_ _05892_ _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13123_ rbzero.spi_registers.texadd3\[11\] _06921_ _06924_ rbzero.spi_registers.texadd2\[11\]
+ _06917_ rbzero.spi_registers.texadd1\[11\] _06937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_21_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_26089_ _06846_ _03024_ _06844_ _06853_ _11825_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_18980_ rbzero.tex_g0\[26\] rbzero.tex_g0\[25\] _11861_ _11863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_108_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14497__A2 _07898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17931_ _11017_ _11075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13054_ gpout0.hpos\[5\] _06871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21767__B2 _09953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17862_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] _11006_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_233_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19601_ _12335_ _12371_ _12372_ _12373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_17_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_7__f_i_clk clknet_3_1_0_i_clk clknet_5_7__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17986__A3 _07775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16813_ _10243_ _10212_ _10244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17793_ _10936_ _10959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__17291__I _10611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24181__A2 _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19532_ _12303_ _12304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16744_ _10176_ _08181_ _10184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_220_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13956_ _07149_ _07194_ _07697_ _07767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_191_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19463_ _12232_ _12234_ _12235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16675_ _10115_ _10116_ _10119_ _10120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16946__A1 _10359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13887_ rbzero.debug_overlay.playerY\[-2\] _07698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_122_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20742__A2 _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13324__I _07137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18414_ _11513_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15626_ _09240_ _09289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_19394_ _12165_ _12166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_185_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14421__A2 _08227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24484__A3 _05228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18345_ _10220_ _11473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_228_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15557_ rbzero.spi_registers.buf_texadd1\[3\] _09232_ _09237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14508_ _07831_ _08317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15488_ rbzero.spi_registers.texadd0\[9\] _09176_ _09186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18276_ rbzero.wall_tracer.mapX\[8\] _11410_ _11418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_155_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput20 i_reg_mosi net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17227_ rbzero.pov.spi_buffer\[10\] _10576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__19648__B1 _12419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14439_ _08247_ _08248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20258__A1 _12984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17158_ rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\] _10523_ _10524_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_80_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17123__A1 rbzero.pov.ready_buffer\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16109_ rbzero.spi_registers.buf_texadd0\[18\] _09644_ _09651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17089_ rbzero.debug_overlay.vplaneX\[-2\] _10471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_229_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14488__A2 _08210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21758__A1 _09998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16229__A3 _09669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24299__I _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22810_ _02485_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_197_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24172__A2 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23790_ rbzero.wall_tracer.trackDistY\[3\] _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22183__A1 _11094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14660__A2 _07938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22741_ _03586_ _02443_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_189_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_151_i_clk clknet_5_11__leaf_i_clk clknet_leaf_151_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_175_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_175_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25460_ _06232_ _06243_ _06244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22672_ _03534_ _03540_ _03541_ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14412__A2 _08210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24411_ net55 _05191_ _05192_ _05194_ _05195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_21623_ _10449_ _02694_ _02700_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25391_ _06122_ _06128_ _06175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_192_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23683__A1 _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27130_ _01040_ clknet_leaf_121_i_clk rbzero.traced_texVinit\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24342_ _05014_ _05051_ _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_145_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21554_ _02623_ _02638_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_166_i_clk clknet_5_8__leaf_i_clk clknet_leaf_166_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_117_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20505_ _12491_ _12917_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27061_ _00971_ clknet_leaf_147_i_clk rbzero.tex_b1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24273_ _05056_ _05057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_105_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15912__A2 _09498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21485_ _02569_ _02565_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26012_ _06772_ _06740_ _06788_ _06789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20249__A1 rbzero.wall_tracer.stepDistY\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23224_ _03652_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_133_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13923__A1 _07214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20436_ _12311_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_200_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13923__B2 _07102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21997__A1 _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23155_ _03892_ _03893_ _03896_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16280__I _09742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20367_ _01384_ _01459_ _01460_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_56_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22106_ _03079_ _03099_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_73_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_227_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23086_ _03939_ _03942_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20298_ _01391_ _01392_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_8_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21749__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22037_ _02997_ _03045_ _03047_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26914_ _00824_ clknet_leaf_134_i_clk rbzero.tex_r1\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
Xclkbuf_leaf_104_i_clk clknet_5_30__leaf_i_clk clknet_leaf_104_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_228_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_199_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26845_ _00755_ clknet_leaf_193_i_clk rbzero.tex_r0\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_240_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_24_i_clk_I clknet_5_20__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13810_ _07616_ _07618_ _07619_ _07620_ _07604_ _07621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_14790_ rbzero.tex_b0\[2\] _07932_ _08597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23988_ rbzero.wall_tracer.rcp_fsm.i_data\[4\] _08813_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26776_ _00686_ clknet_leaf_127_i_clk rbzero.tex_g1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_187_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13741_ _07544_ _07547_ _07548_ _07550_ _07551_ _07552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xclkbuf_leaf_119_i_clk clknet_5_18__leaf_i_clk clknet_leaf_119_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_25727_ _06427_ _06465_ _06510_ _06511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22939_ _03791_ _03793_ _03796_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_35_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16928__A1 _07676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19590__A2 _11081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16460_ _09917_ _09918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_27_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13672_ _07482_ _07483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25658_ _06435_ _06441_ _06442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_27_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14403__A2 _08210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15411_ _09077_ _09131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24609_ _05352_ _05393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_16391_ _09814_ _09863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25589_ _06318_ _06319_ _06371_ _06372_ _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_54_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20488__A1 _12675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18145__A3 _11288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15342_ _09029_ _09080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18130_ rbzero.debug_overlay.playerX\[2\] _11116_ _11249_ rbzero.debug_overlay.playerX\[3\]
+ _11274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_93_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27328_ _01233_ clknet_leaf_115_i_clk rbzero.traced_texa\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_249_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24218__A3 _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18061_ rbzero.wall_tracer.trackDistX\[-9\] _11205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15273_ _09025_ _09026_ _09018_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_27259_ _01164_ clknet_leaf_95_i_clk rbzero.wall_tracer.visualWallDist\[-1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17012_ _10385_ _10414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14224_ _08031_ _08033_ _08034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_112_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25179__A1 _05912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14155_ _07801_ _07960_ _07964_ _07965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__17656__A2 rbzero.pov.ready_buffer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13106_ _06914_ _06920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14086_ _07891_ _07892_ _07893_ _07895_ _07648_ _07896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_18963_ _11853_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_238_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17914_ _08088_ _11004_ _11058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18894_ _11769_ _11808_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20412__A1 _12422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14890__A2 _08518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17845_ _10987_ _10992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_245_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16092__A1 _08977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14578__C _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17776_ _10943_ _10687_ _10947_ _10948_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_135_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14988_ _07164_ _08779_ _08781_ gpout1.clk_div\[1\] net10 _08790_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__22165__B2 _11068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14642__A2 _07920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19515_ rbzero.wall_tracer.stepDistX\[-4\] _12287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_92_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16727_ _10167_ _10168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13939_ _07739_ _07749_ _07750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16793__C _10221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19446_ _12178_ rbzero.wall_tracer.rayAddendY\[-2\] _12182_ _12217_ _12218_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_157_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16658_ _10015_ _10103_ _10104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_233_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_83_i_clk clknet_5_28__leaf_i_clk clknet_leaf_83_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15609_ rbzero.spi_registers.texadd1\[16\] _09268_ _09276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19377_ rbzero.tex_b1\[63\] rbzero.tex_b1\[62\] _12151_ _12154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16589_ rbzero.wall_tracer.rayAddendY\[3\] _10038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18328_ _07205_ _08872_ _11460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_155_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_211_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18259_ _11398_ _11402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_98_i_clk clknet_5_27__leaf_i_clk clknet_leaf_98_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_170_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21270_ _12685_ _02213_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_170_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20221_ _12410_ _12258_ _12993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18844__A1 rbzero.traced_texa\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17647__A2 rbzero.pov.ready_buffer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18695__I1 rbzero.tex_r1\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_21_i_clk clknet_5_5__leaf_i_clk clknet_leaf_21_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_20152_ _12879_ _12923_ _12924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24393__A2 _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24960_ _05734_ _05735_ _05744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20083_ _12847_ _12853_ _12823_ _12854_ _12855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14881__A2 _08631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23911_ rbzero.wall_tracer.rcp_fsm.operand\[-11\] _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24891_ _05621_ _05622_ _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_51_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16083__A1 _08968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_i_clk clknet_5_5__leaf_i_clk clknet_leaf_36_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_222_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23842_ _04533_ _04672_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26630_ _00540_ clknet_leaf_161_i_clk rbzero.tex_b0\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA_clkbuf_leaf_198_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22156__A1 _11988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input12_I i_gpout2_sel[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23773_ _11170_ _04589_ _04612_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26561_ _00471_ clknet_leaf_63_i_clk rbzero.pov.spi_buffer\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_200_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20985_ _02065_ _02073_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_170_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25512_ _06293_ _06294_ _06295_ _06148_ net57 _06296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_22724_ _03548_ _03585_ _03587_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19572__A2 _11079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26492_ _00402_ clknet_leaf_56_i_clk rbzero.debug_overlay.facingY\[-8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25443_ _06226_ _06189_ _06185_ _06227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_149_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22655_ _03524_ _03525_ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_250_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21606_ _02308_ _02688_ _02690_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25374_ _06152_ _06156_ _06157_ _06158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__24492__I _05275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16138__A2 _09669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22586_ _03474_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19586__I _12357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24325_ _04965_ _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14149__A1 _07888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27113_ _01023_ clknet_leaf_141_i_clk rbzero.tex_b1\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_211_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21537_ _02480_ _02492_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22226__B _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27044_ _00954_ clknet_leaf_159_i_clk rbzero.tex_g0\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24256_ _04854_ _05040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__19088__A1 _08156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_229_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21468_ _02542_ _02553_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13848__B _07448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23207_ _04062_ _01920_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20419_ _01509_ _01512_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_24187_ _04947_ _04970_ _04887_ _04890_ _04971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_21399_ _02213_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__20642__A1 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23138_ _03909_ _03994_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_242_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__24384__A2 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23069_ _03920_ _03922_ _03925_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_15960_ rbzero.spi_registers.buf_vshift\[4\] _09531_ _09539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_207_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_25__f_i_clk clknet_3_6_0_i_clk clknet_5_25__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__14679__B _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14911_ rbzero.tex_b1\[60\] _07876_ _08717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15891_ rbzero.spi_registers.buf_leak\[3\] _09482_ _09487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20945__A2 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25333__A1 _05869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17630_ _10850_ _10851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26828_ _00738_ clknet_leaf_177_i_clk rbzero.tex_g1\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14842_ _08308_ _08646_ _08647_ _08648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__17810__A2 rbzero.pov.ready_buffer\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14624__A2 _07855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17561_ _10809_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_86_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14773_ _08315_ _08579_ _08580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26759_ _00669_ clknet_5_3__leaf_i_clk gpout0.vpos\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_19300_ _12110_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16512_ rbzero.debug_overlay.vplaneY\[-1\] _09965_ _09966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13724_ _07534_ _07535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17492_ _10759_ _10770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_151_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19231_ _12067_ _12049_ _12050_ _12070_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_184_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16185__I _09675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16443_ _09900_ _09901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13655_ rbzero.row_render.texu\[0\] _07461_ _07463_ _07465_ _07466_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_19162_ _11954_ _11999_ _12005_ _12006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_13586_ _07366_ _07370_ _07395_ _07396_ _07397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_16374_ _09849_ _09850_ _09844_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__21122__A2 _12194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18113_ rbzero.debug_overlay.playerY\[5\] rbzero.wall_tracer.mapY\[5\] _11257_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15325_ _09034_ _09067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_19093_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] _11937_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_164_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18044_ _11166_ _11186_ _11187_ _11188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19079__A1 _08161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15256_ _09014_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13899__B1 _07709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15529__I _09190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14207_ _08016_ _08017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15187_ _08959_ _08960_ _08961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14138_ rbzero.tex_r1\[61\] _07920_ _07948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_130_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19995_ _12761_ _12766_ _12767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_130_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24375__A2 _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18946_ _11843_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14069_ rbzero.tex_r1\[3\] _07878_ _07879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input4_I i_gpout0_sel[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18877_ rbzero.traced_texa\[3\] rbzero.texV\[3\] _11795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_33_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16065__A1 _08946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17828_ _10979_ _10742_ _10975_ _10981_ _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_240_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17801__A2 rbzero.pov.ready_buffer\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22138__A1 rbzero.wall_tracer.visualWallDist\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22138__B2 _11076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25875__A2 _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23886__A1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22689__A2 rbzero.wall_tracer.stepDistX\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17759_ _10936_ _10937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_234_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20770_ _12660_ _01478_ _01747_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_49_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19429_ rbzero.wall_tracer.visualWallDist\[-1\] _12200_ _12201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22440_ _03341_ _07701_ _03382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22310__A1 _11292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22371_ _02784_ _03248_ rbzero.wall_tracer.wall\[1\] _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24110_ _04827_ _04882_ _04851_ _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_21322_ _12203_ _12207_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25090_ _05856_ _05874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_115_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15439__I _09150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24041_ _04818_ _04820_ _04821_ _04824_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_21253_ _12413_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__14343__I rbzero.debug_overlay.facingY\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20204_ _12964_ _12975_ _12976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_21184_ _02271_ _12959_ _02154_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_224_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_183_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14303__A1 _08110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25563__A1 _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24366__A2 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20135_ _12177_ _12907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14303__B2 _08112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25992_ _05212_ _06771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14854__A2 _08258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20066_ _12816_ _12693_ _12782_ _12675_ _12838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_24943_ _05723_ _05726_ _05727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_225_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24874_ _05653_ _05656_ _05657_ _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_224_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14606__A2 _07821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_174_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26613_ _00523_ clknet_leaf_168_i_clk rbzero.tex_b0\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_206_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23825_ _04653_ _04656_ _04657_ _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__23877__A1 rbzero.wall_tracer.stepDistX\[-5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_68_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15902__I _09494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_198_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23756_ _04588_ _04589_ _04597_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26544_ _00454_ clknet_leaf_24_i_clk rbzero.pov.spi_buffer\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_200_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_198_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20968_ _01930_ _02055_ _02056_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_49_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22707_ _11225_ _12287_ _03572_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_165_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23687_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26475_ _00385_ clknet_leaf_40_i_clk rbzero.debug_overlay.playerY\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_20899_ _01930_ _01988_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13440_ _06875_ _06864_ _07251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_81_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25426_ _06203_ _06209_ _06210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22638_ _03511_ _03513_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_235_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__17829__I _09035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25357_ _06137_ _06139_ _06140_ _06141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_24_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13371_ _07170_ _07174_ _07177_ _07182_ _07183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_36_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22569_ _03464_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16733__I _08908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15110_ _08865_ _08896_ _08897_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24308_ _04930_ _05090_ _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16090_ _09634_ _09636_ _09637_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25288_ _06071_ _06060_ _06072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15041_ _08832_ _08833_ _08834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24239_ _05012_ net89 _05023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_160_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27027_ _00937_ clknet_leaf_134_i_clk rbzero.tex_g0\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XFILLER_0_160_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19481__A1 rbzero.wall_tracer.size\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18800_ _07171_ rbzero.tex_r1\[63\] _11729_ _11733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_19780_ _12547_ _12551_ _12552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16992_ _10345_ _10394_ _10398_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__22368__A1 rbzero.mapdxw\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_196_Right_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18731_ _11694_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15943_ _09524_ _09526_ _09520_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_247_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15084__I _08875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18662_ rbzero.tex_r1\[4\] rbzero.tex_r1\[3\] _11651_ _11655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_216_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15874_ rbzero.spi_registers.buf_floor\[5\] _09464_ _09474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_216_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17613_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _10838_ _10839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_204_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14825_ _07563_ _08631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18593_ _11615_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17544_ _10799_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14756_ rbzero.tex_b0\[30\] _08499_ _08562_ _08563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_103_Left_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__22540__A1 rbzero.wall_tracer.visualWallDist\[-5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13707_ _07508_ _07518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17475_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _10760_ _10761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14687_ _08276_ _08494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_156_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19214_ _12009_ _12056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_172_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16426_ _08826_ _09887_ _09889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13638_ _07444_ _07449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_171_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19145_ _08162_ _10063_ _11971_ _11989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_16357_ rbzero.spi_registers.buf_texadd3\[7\] _09829_ _09838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_146_i_clk_I clknet_5_14__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13569_ _07355_ _07378_ _07380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25956__I _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15308_ _08986_ _09054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24045__A1 _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19076_ rbzero.debug_overlay.facingY\[-2\] _11919_ _11920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_2_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16288_ _09785_ _09786_ _09784_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18027_ _11167_ _11168_ _11169_ _11170_ _11171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15239_ _08987_ _09003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_160_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_112_Left_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_240_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25545__B2 _06328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19978_ _12674_ _12750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14836__A2 _08250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_163_Right_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18929_ rbzero.tex_g0\[4\] rbzero.tex_g0\[3\] _11830_ _11834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_158_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19775__A2 _12527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21940_ _11092_ _02978_ _10125_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_158_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21724__I _11399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23859__A1 _12395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21871_ _02913_ _02914_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_222_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_121_Left_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_143_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15722__I _09336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23610_ _04220_ _04327_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20822_ _01812_ _01852_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24590_ _05371_ _05350_ net77 _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_210_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13272__B2 _06926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23541_ _04367_ _04393_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20753_ _01715_ _01843_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_187_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14338__I rbzero.debug_overlay.facingY\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26260_ _00170_ clknet_leaf_241_i_clk rbzero.spi_registers.texadd3\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23472_ _04324_ _04325_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20684_ _01665_ _01772_ _01775_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__22555__I _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_217_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16761__A2 _10183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25211_ _05235_ _05970_ _05993_ _05994_ _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_17_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22423_ _03365_ _03366_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14772__A1 _08565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26191_ _00101_ clknet_leaf_239_i_clk rbzero.spi_registers.texadd0\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25142_ _05919_ _05925_ _05926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22354_ _11140_ _11247_ _03244_ rbzero.wall_tracer.trackDistY\[10\] _03304_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_116_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24036__A1 _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16513__A2 rbzero.wall_tracer.rayAddendY\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21305_ _02390_ _02391_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14524__A1 _08315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25073_ _05793_ _05796_ _05857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_103_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22285_ _11377_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_131_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22598__A1 _07236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24024_ _04805_ _04807_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_103_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21236_ _02318_ _02319_ _02322_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__21270__A1 _12685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21167_ _02136_ _02253_ _02254_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_141_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14827__A2 _07932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20118_ _12560_ _12500_ _12890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25975_ _06737_ _05028_ _06654_ _06755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_21098_ _02065_ _02073_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_102_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_226_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_20049_ _12819_ _12820_ _12821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24926_ _05689_ _05690_ _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_232_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24010__I _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24857_ _05311_ _05641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16728__I _10168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_237_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14610_ rbzero.tex_g1\[4\] _07563_ _08418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_23808_ _04639_ _04642_ _04594_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_240_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_237_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15590_ _09261_ _09262_ _09253_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24788_ _05410_ _05347_ _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_157_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__21325__A2 _12647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18577__I0 rbzero.tex_r0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23989__C _11473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14541_ rbzero.tex_g0\[59\] _08340_ _08350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26527_ _00437_ clknet_leaf_38_i_clk rbzero.pov.spi_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23739_ rbzero.wall_tracer.trackDistY\[-4\] _03050_ _04577_ _04582_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17260_ _10598_ _10594_ _10600_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_126_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14472_ rbzero.tex_g0\[39\] _08279_ _08280_ _08281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_26458_ _00368_ clknet_leaf_206_i_clk rbzero.debug_overlay.playerX\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16211_ rbzero.spi_registers.buf_texadd1\[19\] _09719_ _09728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25409_ _06184_ _06188_ _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13423_ _07233_ _07234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14763__A1 rbzero.tex_b0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13566__A2 _06884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17191_ rbzero.pov.spi_buffer\[1\] _10549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_183_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22825__A2 _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26389_ _00299_ clknet_leaf_20_i_clk rbzero.spi_registers.buf_texadd2\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__26016__A2 rbzero.wall_tracer.rcp_fsm.o_data\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16142_ _09660_ _09678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13354_ _07165_ _07166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_181_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13318__A2 _07111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14515__A1 _08321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16073_ _08957_ _09624_ _09625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13285_ _07063_ _07093_ _07098_ _07099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_19901_ _12240_ _12672_ _12673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15024_ _08818_ net19 _08819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__18257__A2 _11400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_236_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16268__A1 _08948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19832_ _12603_ _12539_ _12604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__25527__A1 _05996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14711__I _07566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19763_ _12456_ _12534_ _12535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_235_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16975_ _08932_ _10385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_235_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18714_ _11684_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15926_ _08912_ _09498_ _09513_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19694_ _12437_ _12443_ _12466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_127_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 net81 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_160_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_72_i_clk_I clknet_5_29__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18645_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _11644_ _11645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15857_ _08912_ _09460_ _09461_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_204_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_19__f_i_clk_I clknet_3_4_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16440__A1 _07241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19014__I _11871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14808_ _07432_ _07473_ _08361_ _08615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_188_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18576_ _11605_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15788_ rbzero.spi_registers.buf_texadd3\[13\] _09409_ _09410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17527_ rbzero.tex_b0\[24\] rbzero.tex_b0\[23\] _10786_ _10790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14739_ rbzero.tex_b0\[33\] _08233_ _08546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_200_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17458_ rbzero.pov.spi_buffer\[69\] _10748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17940__A1 _11074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13997__I _07518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer2_I _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16409_ rbzero.spi_registers.spi_buffer\[20\] _09876_ _09877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17389_ _10696_ _10697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__26007__A2 _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19128_ _08162_ _10062_ _11972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_232_Right_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19059_ _11907_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22070_ rbzero.wall_tracer.stepDistY\[6\] _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21252__A1 _12465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21021_ _02108_ _02109_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__13190__B1 _06992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21004__A1 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25760_ _06518_ _06543_ _06544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22972_ _03810_ _03829_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24711_ _05444_ _05449_ _05495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21923_ _11033_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25691_ _06445_ _06473_ _06475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_223_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27430_ _01335_ clknet_leaf_69_i_clk rbzero.wall_tracer.rcp_fsm.operand\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24642_ _05424_ _05425_ _05426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_171_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21854_ _02894_ _02896_ _02898_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_219_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21307__A2 _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22504__A1 rbzero.wall_tracer.size\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20805_ _01781_ _01891_ _01894_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_27361_ _01266_ clknet_leaf_103_i_clk rbzero.wall_tracer.trackDistX\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14993__A1 _07171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14068__I _07483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24573_ _05295_ _05356_ _05357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21785_ _10036_ _02834_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26312_ _00222_ clknet_leaf_235_i_clk rbzero.spi_registers.buf_vshift\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20736_ _01823_ _01826_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_23524_ _04223_ _04214_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27292_ _01197_ clknet_leaf_211_i_clk rbzero.row_render.size\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__22285__I _11377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_232_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23455_ _02249_ _04308_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14745__A1 _07888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26243_ _00153_ clknet_leaf_21_i_clk rbzero.spi_registers.texadd2\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_98_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20667_ _01484_ _12957_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13700__I _07418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20818__A1 _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22406_ _03345_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_208_Left_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23386_ _04133_ _04240_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_26174_ _00084_ clknet_leaf_222_i_clk rbzero.color_floor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20598_ _01688_ _01689_ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25125_ _05908_ _05871_ _05909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__20294__A2 _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22337_ _11282_ _03290_ _03278_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16498__B2 _09953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20833__A4 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25056_ _05472_ _05840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15170__A1 _08946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13070_ gpout0.hpos\[4\] _06886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_210_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22268_ rbzero.wall_tracer.visualWallDist\[-6\] _03218_ _03229_ _03234_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24007_ _04792_ _04793_ _04786_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__21243__A1 _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15627__I _09289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21219_ rbzero.traced_texVinit\[7\] _01778_ _02306_ _02034_ _02307_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14531__I _07831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22199_ _10151_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_218_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_245_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22043__I0 rbzero.wall_tracer.rcp_fsm.o_data\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16670__A1 _08096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16760_ _10194_ _10197_ _10198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_25958_ _05212_ _06739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_217_Left_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13972_ _07247_ _07781_ _07782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18798__I0 rbzero.tex_r1\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15711_ _09352_ _09353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24909_ _05672_ _05674_ _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_220_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16691_ _10132_ _10112_ _10134_ _10135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__16458__I _09895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25889_ _05027_ _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_201_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18430_ _11479_ _11522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15642_ _09289_ _09301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_107_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24496__A1 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13787__A2 _07597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18361_ _11483_ _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15573_ rbzero.spi_registers.texadd1\[7\] _09243_ _09249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18673__I _11650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18175__A1 rbzero.map_overlay.i_othery\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18175__B2 _07732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17312_ _10637_ _10630_ _10639_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14524_ _08315_ _08325_ _08332_ _08333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_18292_ _10271_ _11431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24248__B2 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22128__C _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13539__A2 _07349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17243_ _10564_ _10588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14455_ _07479_ _08264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_226_Left_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13406_ _07196_ _07197_ _07217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_142_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17174_ rbzero.pov.spi_counter\[3\] rbzero.pov.spi_counter\[2\] rbzero.pov.spi_counter\[1\]
+ _10513_ _10535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_clkbuf_leaf_19_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19718__B _12342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14386_ _08195_ reg_rgb\[1\] _08196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17525__I1 rbzero.tex_b0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16125_ _09662_ _09663_ _09661_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13337_ _07064_ _07147_ _07150_ _07151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__22144__B _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16056_ _09600_ _09612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__24420__A1 _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13268_ _07064_ _07076_ _07081_ _07082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_121_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13172__B1 _06981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15007_ _08806_ _08807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_209_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14441__I _07532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13199_ _07007_ _07012_ _07013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19815_ _12586_ _12587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_235_Left_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_209_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13057__I _06873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16661__A1 _09998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19746_ _12511_ _12288_ _12516_ _12517_ _12518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_16958_ rbzero.pov.ready_buffer\[58\] _10274_ _10366_ _10369_ _10370_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13475__A1 rbzero.traced_texVinit\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22734__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15909_ _08950_ _09498_ _09501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19677_ _12315_ _12318_ _12328_ _12448_ _12449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_155_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20745__B1 _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16889_ rbzero.pov.ready_buffer\[48\] _10275_ _10311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_205_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18628_ _11635_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23703__B _12036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14975__A1 _07050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18559_ rbzero.tex_r0\[24\] rbzero.tex_r0\[23\] _11592_ _11596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__18166__A1 rbzero.map_overlay.i_mapdy\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21570_ _02649_ _02654_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_244_Left_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__24239__A1 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17199__I _10546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20521_ rbzero.wall_tracer.size_full\[5\] _01527_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14990__A4 _07230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_173_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_190_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23240_ _03725_ _01580_ _03942_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20452_ _01445_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_138_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23171_ _03958_ _03993_ _04026_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_160_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20383_ _01379_ _01476_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13950__A2 rbzero.map_overlay.i_mapdy\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22122_ rbzero.wall_tracer.rcp_fsm.i_data\[-8\] _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_93_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_246_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22053_ _03058_ _03054_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26930_ _00840_ clknet_leaf_173_i_clk rbzero.tex_r1\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_21004_ _02091_ _02092_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22973__A1 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26861_ _00771_ clknet_leaf_192_i_clk rbzero.tex_r0\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__17662__I _10847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25812_ _06581_ _06585_ _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_71_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26792_ _00702_ clknet_leaf_195_i_clk rbzero.tex_g1\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_25743_ _06498_ _06499_ _06496_ _06527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_3_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22955_ _03811_ _03812_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21906_ _10121_ _02947_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24478__A1 _05261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25674_ _06451_ _06457_ _06458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22886_ _03703_ _03744_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_85_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19589__I _12360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27413_ _01318_ clknet_leaf_85_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_66_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24625_ _05296_ _05408_ _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14966__A1 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14966__B2 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21837_ _02872_ _02857_ _02871_ _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27344_ _01249_ clknet_leaf_94_i_clk rbzero.wall_tracer.w\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24556_ _05292_ _05279_ _05290_ _05340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_21768_ _12184_ _02722_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23507_ _04265_ _04339_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15131__B _08909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20719_ _01801_ _01809_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14526__I _07549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14569__I1 _08377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27275_ _01180_ clknet_leaf_205_i_clk rbzero.wall_tracer.texu\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24487_ _05270_ _05271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21699_ _11133_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26226_ _00136_ clknet_leaf_2_i_clk rbzero.spi_registers.texadd1\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_22_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_20_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14240_ _08042_ _08045_ _08047_ _08049_ _08050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__22743__I _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23438_ _03726_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14171_ _07974_ _07981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23369_ _04222_ _04223_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26157_ _00067_ clknet_leaf_221_i_clk rbzero.mapdxw\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13941__A2 rbzero.map_overlay.i_mapdy\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25108_ _05888_ _05891_ _05892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13122_ _06935_ _06936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_26088_ _06851_ _06852_ _06842_ _06853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15357__I _09074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17930_ _11007_ _11019_ _11074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13053_ _06865_ _06869_ _06870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16891__A1 _08062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25039_ _05757_ _05817_ _05822_ _05823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__14261__I rbzero.debug_overlay.facingX\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17861_ rbzero.debug_overlay.facingX\[-4\] _11004_ _11005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_79_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_245_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19600_ _12353_ _12370_ _12372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_206_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16812_ _07677_ _10243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_109_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17792_ _10934_ _10958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22716__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19531_ _12302_ _12303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16743_ _10182_ _10183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13955_ _07750_ _07765_ _07766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16188__I _09711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15092__I _08883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22192__A2 _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19462_ _10224_ _11099_ _12233_ _11390_ _12234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_16674_ _10075_ _10117_ _10118_ _10076_ _10119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_159_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24469__A1 _05252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13886_ _07683_ _07689_ _07692_ _07696_ _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_76_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18413_ rbzero.tex_g1\[25\] rbzero.tex_g1\[24\] _11512_ _11513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15625_ rbzero.spi_registers.buf_texadd1\[20\] _09281_ _09288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14957__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19393_ _12163_ _12164_ _12165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_16_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18344_ _07179_ _11468_ _11472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_201_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15556_ rbzero.spi_registers.texadd1\[3\] _09230_ _09236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14507_ _07501_ _08316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14709__B2 _08284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14436__I _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18275_ _11412_ _11416_ _11417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_155_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15487_ _09184_ _09185_ _09175_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17226_ _10574_ _10572_ _10575_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19648__A1 _12417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 net98 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14438_ _07511_ _08247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput21 i_reg_outs_enb net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__19648__B2 _12267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14880__B _08321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21455__A1 _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17157_ rbzero.pov.sclk_buffer\[2\] _09015_ _10523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14369_ _07701_ _08011_ _08017_ _08171_ _08178_ _08179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_123_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16108_ _09649_ _09650_ _09648_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17088_ _10469_ _10470_ _10462_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16039_ _08851_ _09544_ _09599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_21_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_243_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19820__A1 _08181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15437__A2 _09148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24172__A3 _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19729_ _12500_ _12501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13999__A2 _07807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13515__I _07325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22740_ _11169_ _03599_ _03601_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_189_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21930__A2 _10478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22671_ rbzero.wall_tracer.trackDistX\[-9\] _03533_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14948__A1 _06873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16826__I _10255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19202__I _12044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24410_ _05186_ _05073_ _05193_ _05163_ _05194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_21622_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] _02700_
+ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_177_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25390_ _06131_ _06173_ _06130_ _06174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24341_ _05120_ _05124_ _05125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21553_ _02628_ _02631_ _02637_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_74_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20504_ _12999_ _12645_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24272_ _04940_ _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27060_ _00970_ clknet_leaf_148_i_clk rbzero.tex_b1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21484_ _02447_ _02448_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_194_i_clk_I clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26011_ _06634_ _06787_ _06788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20249__A2 _12311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23223_ _04078_ _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20435_ rbzero.wall_tracer.size_full\[4\] _01430_ _01528_ _01529_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_200_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13923__A2 _07732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23154_ _03892_ _03893_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23595__S _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20366_ _01387_ _01393_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_160_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__23199__A1 _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22105_ rbzero.wall_tracer.rcp_fsm.i_data\[-11\] _03088_ _03098_ _03099_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23085_ _03940_ _03941_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20297_ _12210_ _12963_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_227_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22036_ _03046_ _03039_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26913_ _00823_ clknet_leaf_135_i_clk rbzero.tex_r1\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_101_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26844_ _00754_ clknet_leaf_194_i_clk rbzero.tex_r0\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_215_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_240_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15126__B _08909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26775_ _00685_ clknet_leaf_128_i_clk rbzero.tex_g1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23987_ rbzero.wall_tracer.rcp_fsm.operand\[4\] _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_205_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25726_ _06431_ _06464_ _06510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13740_ _07331_ _07551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22938_ _03794_ _03795_ _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_225_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17050__A1 _08159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21921__A2 _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25112__A2 _05408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25657_ _06439_ _06440_ _06441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_168_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13671_ _07481_ _07482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16736__I _08180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22869_ _03726_ _03727_ _02670_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_27_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15410_ rbzero.color_sky\[5\] _09129_ _09130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24608_ _05389_ _05391_ _05392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_183_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16390_ _09861_ _09862_ _09856_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25588_ _06321_ _06370_ _06372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20488__A2 _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15341_ _09076_ _09079_ _09073_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_27327_ _01232_ clknet_leaf_115_i_clk rbzero.traced_texa\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24539_ _05256_ _05319_ _05322_ _05323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_136_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18060_ _11201_ _11204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_27258_ _01163_ clknet_leaf_94_i_clk rbzero.wall_tracer.visualWallDist\[-2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15272_ rbzero.spi_registers.buf_otherx\[3\] _09021_ _09026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17011_ rbzero.pov.ready_buffer\[42\] _10412_ _10413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21437__A1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26209_ _00119_ clknet_leaf_239_i_clk rbzero.spi_registers.texadd1\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14223_ _07987_ _08032_ _08033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
XANTENNA__16471__I _08112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13914__A2 rbzero.map_overlay.i_othery\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_27189_ _01094_ clknet_leaf_78_i_clk rbzero.wall_tracer.size\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_21_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14154_ _07475_ _07961_ _07962_ _07963_ _07437_ _07964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_81_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13105_ rbzero.spi_registers.texadd1\[15\] _06918_ _06919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_2_i_clk clknet_5_1__leaf_i_clk clknet_leaf_2_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14085_ rbzero.tex_r1\[32\] _07894_ _07808_ _07895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18962_ rbzero.tex_g0\[18\] rbzero.tex_g0\[17\] _11851_ _11853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_211_i_clk clknet_5_16__leaf_i_clk clknet_leaf_211_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17913_ _11006_ _11055_ _11056_ _11057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18893_ rbzero.traced_texa\[6\] _07273_ _11807_ _11808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_119_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15815__I _09429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17844_ _10990_ _10849_ _10988_ _10991_ _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_28_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17775_ _10944_ rbzero.pov.ready_buffer\[48\] _10948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_156_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14987_ _08782_ _08788_ _08789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_226_i_clk clknet_5_2__leaf_i_clk clknet_leaf_226_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_19514_ _12265_ _12285_ _12286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16726_ _08875_ _10166_ _10167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_199_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13938_ _07745_ _07748_ _07749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14875__B _08308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19445_ _12183_ _12216_ _12217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16657_ _10097_ _10098_ _10101_ _10103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_157_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13869_ rbzero.debug_overlay.playerX\[0\] _07077_ _07680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15550__I _09208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15608_ _09274_ _09275_ _09267_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_186_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19376_ _12153_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__19869__A1 rbzero.wall_tracer.size\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16588_ _01029_ _10029_ _10037_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__23665__A2 _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18327_ _07760_ _11432_ _11457_ _11459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_84_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21676__A1 _10346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15539_ rbzero.spi_registers.buf_texadd0\[22\] _09030_ _09224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_211_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18258_ _11127_ _11128_ _11398_ _11401_ _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_154_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17209_ _10561_ _10559_ _10562_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18189_ rbzero.map_rom.d6 _11333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_130_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20220_ _12990_ _12891_ _12991_ _12992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_228_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15658__A2 _09306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20151_ _12900_ _12922_ _12923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_38_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21727__I _11134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20082_ _12822_ _12814_ _12821_ _12854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__20631__I _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_185_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23910_ _04717_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16607__B2 _10049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24890_ _05673_ _05674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_51_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_222_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23841_ _04568_ _04671_ _04446_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_240_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26560_ _00470_ clknet_5_21__leaf_i_clk rbzero.pov.spi_buffer\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23772_ _03603_ _04611_ _04560_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20984_ _02070_ _02072_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_212_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17032__A1 _08161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25511_ _06151_ _06158_ _06295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_177_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22723_ _03586_ _02167_ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_26491_ _00401_ clknet_leaf_56_i_clk rbzero.debug_overlay.facingY\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_193_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25442_ _06075_ _06001_ _06226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_165_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22654_ _03524_ _03525_ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21605_ rbzero.traced_texVinit\[10\] _02689_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25373_ _06133_ _06134_ _06157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_22585_ _09917_ _03473_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_36_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27112_ _01022_ clknet_leaf_142_i_clk rbzero.tex_b1\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24324_ _04957_ _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15346__A1 _07754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21536_ _02611_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_69_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24605__A1 _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21419__A1 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27043_ _00953_ clknet_leaf_159_i_clk rbzero.tex_g0\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24255_ _04898_ _05034_ _04953_ _05035_ _05036_ _05038_ _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_21467_ _02544_ _02552_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_229_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_177_Right_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_161_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17099__A1 _10478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20418_ _01510_ _01511_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22092__A1 _11393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23206_ _02540_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_21398_ _01948_ _02482_ _02351_ _02483_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_24186_ _04818_ _04820_ _04970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_31_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15649__A2 _09306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23137_ _03958_ _03993_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20349_ _01398_ _01443_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_242_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_242_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23068_ _03923_ _03924_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_207_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_158_Left_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22019_ _03032_ _03034_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14910_ rbzero.tex_b1\[62\] _08698_ _08603_ _08716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15890_ _09485_ _09486_ _09473_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26827_ _00737_ clknet_leaf_177_i_clk rbzero.tex_g1\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14841_ rbzero.tex_b1\[23\] _07633_ _08647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_243_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14085__A1 rbzero.tex_r1\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15821__A2 _09118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17560_ rbzero.tex_b0\[38\] rbzero.tex_b0\[37\] _10807_ _10809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26758_ _00668_ clknet_leaf_222_i_clk gpout0.vpos\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14772_ _08565_ _08575_ _08578_ _08579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_203_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16511_ rbzero.wall_tracer.rayAddendY\[-1\] _09965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__17023__A1 _08156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25709_ _06031_ _06051_ _05978_ _06493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_13723_ _07418_ _07534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__18220__B1 _11300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17491_ _10769_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17071__B _10436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25097__A1 _05880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26689_ _00599_ clknet_leaf_64_i_clk rbzero.pov.ready_buffer\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15370__I _09054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19230_ _12067_ _12062_ _12069_ _12070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_16442_ _09899_ _09900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_184_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13654_ _07464_ _07465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_167_Left_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19161_ _12004_ _12005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_27_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21658__A1 _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16373_ rbzero.spi_registers.spi_buffer\[11\] _09842_ _09850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_186_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13585_ _07366_ _07039_ _07044_ _07396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18112_ rbzero.map_rom.a6 _11256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__22417__B _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15324_ rbzero.spi_registers.buf_mapdx\[5\] _09038_ _09066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19092_ _11925_ _11935_ _11923_ _11936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18043_ _11160_ rbzero.wall_tracer.trackDistY\[4\] _11163_ _11164_ _11187_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_152_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15255_ _08818_ rbzero.pov.sclk_buffer\[0\] _09014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_227_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13899__A1 _07707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13899__B2 _07060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14206_ _07998_ _08015_ _08016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_10_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15186_ _08916_ _08960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_150_i_clk clknet_5_11__leaf_i_clk clknet_leaf_150_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__20633__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14137_ rbzero.tex_r1\[63\] _07938_ _07946_ _07947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19994_ _12764_ _12765_ _12766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_130_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_176_Left_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18945_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _11840_ _11843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14068_ _07483_ _07878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22386__A2 _08029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22630__I0 rbzero.wall_tracer.texu\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18876_ _11786_ _11793_ _11794_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_146_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_165_i_clk clknet_5_10__leaf_i_clk clknet_leaf_165_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_176_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_142_i_clk_I clknet_5_14__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17827_ _10980_ rbzero.pov.ready_buffer\[67\] _10981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14076__A1 _07803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17758_ _10843_ _10936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_221_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17014__A1 _08076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16709_ _09988_ _10151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17689_ _10890_ rbzero.pov.ready_buffer\[19\] _10891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_175_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_185_Left_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19428_ _12199_ _12200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19359_ rbzero.tex_b1\[55\] rbzero.tex_b1\[54\] _12141_ _12144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_103_i_clk clknet_5_30__leaf_i_clk clknet_leaf_103_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15328__A1 rbzero.map_overlay.i_mapdy\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22370_ _03306_ _03317_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21321_ _02256_ _02406_ _02407_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_67_i_clk_I clknet_5_21__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23937__I _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24040_ _04796_ _04822_ _04823_ rbzero.wall_tracer.rcp_fsm.operand\[4\] _04824_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_21252_ _12465_ _01944_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_118_i_clk clknet_5_19__leaf_i_clk clknet_leaf_118_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_229_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_194_Left_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20203_ _12966_ _12974_ _12975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_21183_ _02001_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_8__f_i_clk_I clknet_3_2_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_229_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_224_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20134_ _12277_ _12906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_224_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25991_ _06764_ _06767_ _06769_ _06770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__25563__A2 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15455__I _09150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20065_ _12836_ _12837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24942_ _05724_ _05719_ _05725_ _05687_ _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__22621__I0 rbzero.wall_tracer.texu\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24873_ _05654_ _05655_ _05657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__18766__I _11713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26612_ _00522_ clknet_leaf_168_i_clk rbzero.tex_b0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23824_ _04653_ _04656_ _04594_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_213_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17005__A1 _08071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26543_ _00453_ clknet_leaf_24_i_clk rbzero.pov.spi_buffer\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_198_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23755_ _03587_ _04596_ _04560_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_239_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20967_ _01933_ _01987_ _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_215_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_246_Right_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22706_ _11192_ _12243_ _03571_ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26474_ _00384_ clknet_leaf_208_i_clk rbzero.debug_overlay.playerY\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23686_ _04535_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20898_ _01933_ _01987_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_193_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25425_ _06204_ _06207_ _06208_ _06209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_81_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22637_ _03508_ _03512_ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_192_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22301__A2 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15319__A1 _07743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25356_ _06136_ _06104_ _06105_ _06140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_24_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13370_ _07179_ _07154_ _07158_ _07180_ _07159_ _07181_ _07182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_146_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22568_ _11282_ _03461_ _03462_ rbzero.traced_texa\[6\] _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14790__A2 _07932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24307_ _05090_ _05091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_180_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21519_ _02600_ _02603_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25287_ _06064_ _06070_ _06071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22499_ _03421_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_146_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15040_ _08823_ rbzero.spi_registers.spi_cmd\[2\] _08833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_27026_ _00936_ clknet_leaf_132_i_clk rbzero.tex_g0\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_239_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24238_ _05021_ _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22751__I _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24169_ _04730_ _04908_ _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_112_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_82_i_clk clknet_5_28__leaf_i_clk clknet_leaf_82_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16991_ rbzero.pov.ready_buffer\[37\] _10397_ _10398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_235_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17619__I0 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15942_ _09525_ _09507_ _09526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18730_ rbzero.tex_r1\[33\] rbzero.tex_r1\[32\] _11693_ _11694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24109__A3 _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18661_ _11654_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15873_ _09471_ _09472_ _09473_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_188_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17612_ _10822_ _10838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14824_ rbzero.tex_b1\[31\] _08252_ _08630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_192_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_97_i_clk clknet_5_26__leaf_i_clk clknet_leaf_97_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_18592_ rbzero.tex_r0\[38\] rbzero.tex_r0\[37\] _11613_ _11615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17543_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _10796_ _10799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14755_ rbzero.tex_b0\[31\] _07499_ _08562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_169_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13706_ _07510_ _07512_ _07514_ _07516_ _07495_ _07517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_169_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17474_ _10759_ _10760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_213_Right_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14686_ rbzero.color_sky\[4\] rbzero.color_floor\[4\] _07966_ _08493_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_20_i_clk clknet_5_5__leaf_i_clk clknet_leaf_20_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_129_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16425_ _08903_ _09886_ _09888_ _08894_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_19213_ rbzero.wall_tracer.mapY\[8\] _12016_ _12055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_15_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13637_ _07443_ _07448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25490__A1 _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19144_ _11973_ _11987_ _11988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_171_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16356_ _09836_ _09837_ _09833_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20303__A1 _12982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14781__A2 _08300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13568_ _07362_ _06873_ _07376_ _07377_ _06863_ _07378_ _07379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XANTENNA__13584__A3 _07039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15307_ rbzero.spi_registers.buf_mapdx\[1\] _09045_ _09053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19075_ rbzero.wall_tracer.rayAddendY\[6\] _11919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_132_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16287_ rbzero.spi_registers.spi_buffer\[13\] _09782_ _09786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_35_i_clk clknet_5_5__leaf_i_clk clknet_leaf_35_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13499_ _07284_ _07309_ _07310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22056__A1 rbzero.wall_tracer.stepDistY\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18026_ rbzero.wall_tracer.trackDistY\[0\] _11170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_152_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15238_ _09000_ _09001_ _09002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15169_ rbzero.spi_registers.spi_buffer\[6\] _08946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19977_ _12746_ _12748_ _12749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_165_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15275__I _08876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18928_ _11833_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_197_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_18859_ rbzero.traced_texa\[0\] rbzero.texV\[0\] _11780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_206_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17786__A2 rbzero.pov.ready_buffer\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15797__A1 rbzero.spi_registers.buf_texadd3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21870_ _10482_ _08142_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_143_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20821_ _01854_ _01885_ _01910_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13272__A2 _07026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23540_ _04372_ _04392_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20752_ rbzero.wall_tracer.stepDistY\[7\] _01838_ _01839_ _01842_ _01843_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_147_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20683_ _01773_ _01774_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23471_ _03979_ _04214_ _04175_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_63_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_217_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25210_ _05880_ _05987_ _05994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22422_ _03354_ _03357_ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26190_ _00100_ clknet_leaf_237_i_clk rbzero.spi_registers.texadd0\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25141_ _05924_ _05925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_150_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22353_ _03210_ _03302_ _03303_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_143_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22047__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21304_ _02384_ _02389_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25072_ _05854_ _05855_ _05856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_22284_ _11174_ _03243_ _03244_ _03246_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_170_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15721__A1 rbzero.spi_registers.buf_texadd2\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22598__A2 _11394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24023_ _04794_ rbzero.wall_tracer.rcp_fsm.operand\[1\] _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21235_ _02252_ _02265_ _02321_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_229_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_245_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_21166_ _01996_ _01859_ _02137_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_20117_ _12410_ _12274_ _12889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25974_ _05261_ _06753_ _05087_ _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_21097_ _02183_ _02184_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20048_ _12812_ _12813_ _12820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24925_ _05672_ _05674_ _05709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_137_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15913__I _09428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17777__A2 rbzero.pov.ready_buffer\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24856_ _05320_ _05640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_212_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23807_ _04640_ _04634_ _04641_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_237_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24787_ _05287_ _05271_ _05361_ _05571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_21999_ _02991_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13433__I gpout0.vpos\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14540_ _08339_ _08347_ _08348_ _08349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_26526_ _00436_ clknet_leaf_213_i_clk rbzero.pov.spi_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23738_ _11191_ _03050_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_233_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14471_ _07489_ _08280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26457_ _00367_ clknet_leaf_206_i_clk rbzero.debug_overlay.playerX\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23669_ rbzero.wall_tracer.stepDistX\[10\] _04519_ _04520_ _04521_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16210_ _09726_ _09727_ _09723_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_12_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25408_ _06186_ _06190_ _06191_ _06192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_13422_ rbzero.trace_state\[0\] _07233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17190_ _10538_ _10545_ _10548_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14763__A2 _08448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26388_ _00298_ clknet_leaf_20_i_clk rbzero.spi_registers.buf_texadd2\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__19151__A1 rbzero.wall_tracer.rayAddendY\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16141_ _09591_ _09676_ _09677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25339_ _06079_ _06080_ _06081_ _05724_ _06123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_13353_ net23 _07165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16072_ _09600_ _09624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22481__I _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13284_ _07050_ _07094_ _07097_ _07074_ _07098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_121_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19900_ _12608_ _12671_ _12672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_224_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15023_ _08806_ _08818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_27009_ _00919_ clknet_leaf_189_i_clk rbzero.tex_g0\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__19454__A2 _12006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19831_ _12510_ _12532_ _12603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15095__I _08810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13608__I _07418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19762_ _12461_ _12505_ _12533_ _12534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_78_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16974_ rbzero.pov.ready_buffer\[34\] _10383_ _10384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18713_ rbzero.tex_r1\[26\] rbzero.tex_r1\[25\] _11682_ _11684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_217_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15925_ rbzero.spi_registers.buf_othery\[0\] _09507_ _09478_ _09513_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19693_ _12464_ _12465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_30_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16919__I _10336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 i_gpout1_sel[0] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_15_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15856_ rbzero.spi_registers.buf_floor\[0\] _09459_ _08909_ _09461_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18644_ _11628_ _11644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_189_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16440__A2 _08869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14807_ _07802_ _08552_ _08613_ _08614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_125_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18575_ rbzero.tex_r0\[31\] rbzero.tex_r0\[30\] _11602_ _11605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15787_ _09117_ _09409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13343__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17526_ _10789_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14738_ _08540_ _08542_ _08544_ _08284_ _08245_ _08545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_47_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17457_ _10745_ _10746_ _10747_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14669_ _07480_ _08471_ _08476_ _08477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__24266__A2 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17940__A2 _11076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16408_ _09818_ _09876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15951__A1 _09515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14754__A2 _08554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17388_ _10542_ _10696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19142__A1 _08152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19127_ _11924_ _11969_ _11970_ _11971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16339_ rbzero.spi_registers.buf_texadd3\[2\] _09816_ _09825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24092__B _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22029__A1 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19058_ rbzero.tex_g0\[60\] rbzero.tex_g0\[59\] _11903_ _11907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18009_ rbzero.wall_tracer.trackDistX\[7\] _11150_ rbzero.wall_tracer.trackDistX\[6\]
+ _11151_ _11152_ _11153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_51_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19445__A2 _12216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21020_ _01962_ _01985_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_140_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13518__I _07328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22201__A1 _11282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22971_ _03820_ _03828_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__16829__I _07687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24710_ _05444_ _05449_ _05494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_207_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21922_ _10040_ _02961_ _02962_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25690_ _06445_ _06473_ _06474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_222_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24641_ _05368_ _05369_ _05425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_136_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14349__I rbzero.debug_overlay.facingY\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21853_ _02880_ _02881_ _02897_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_219_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_195_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27360_ _01265_ clknet_leaf_103_i_clk rbzero.wall_tracer.trackDistX\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20804_ _01784_ _01890_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24572_ _05229_ _05356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_148_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__26038__I _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21784_ _02829_ _02832_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19381__A1 _11456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26311_ _00221_ clknet_leaf_235_i_clk rbzero.spi_registers.buf_vshift\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23523_ _04373_ _04374_ _04375_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_20735_ _01824_ _01825_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_27291_ _01196_ clknet_leaf_211_i_clk rbzero.row_render.size\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22268__A1 rbzero.wall_tracer.visualWallDist\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26242_ _00152_ clknet_leaf_21_i_clk rbzero.spi_registers.texadd2\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_232_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23454_ _04150_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15942__A1 _09525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20666_ _01756_ _01757_ _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_98_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22405_ _03193_ _03350_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26173_ _00083_ clknet_leaf_223_i_clk rbzero.color_floor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14084__I _07831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20597_ _01596_ _01601_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23385_ _04236_ _04239_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25124_ _05872_ _05907_ _05908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_6_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20294__A3 _12666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22336_ _03200_ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25055_ _05520_ _05308_ _05839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22267_ rbzero.wall_tracer.trackDistY\[-6\] _03226_ _03232_ _03233_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19436__A2 _12207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_210_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24006_ rbzero.wall_tracer.rcp_fsm.i_data\[9\] _04773_ _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21218_ _02171_ _02305_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_247_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22198_ _03154_ _03175_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_228_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21149_ _02231_ _02236_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_228_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25957_ _06737_ _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13971_ _07777_ _07780_ _07781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_232_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16739__I _10178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18798__I1 rbzero.tex_r1\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15710_ _09257_ _09352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_214_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24908_ _05691_ _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16690_ _09990_ _10133_ _10134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_189_i_clk_I clknet_5_9__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25888_ _06667_ _06670_ _06671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_214_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15641_ rbzero.spi_registers.buf_texadd2\[0\] _09293_ _09300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24839_ _05302_ _05324_ _05623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_17_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18360_ rbzero.tex_g1\[2\] rbzero.tex_g1\[1\] _11481_ _11483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_201_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15572_ _09247_ _09248_ _09242_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15799__B _09417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17311_ rbzero.pov.spi_buffer\[32\] _10638_ _10635_ _10639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18175__A2 _11308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14523_ _08245_ _08328_ _08331_ _08332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_26509_ _00419_ clknet_leaf_59_i_clk rbzero.debug_overlay.vplaneX\[-2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_230_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16186__A1 _08973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18291_ _11402_ _11429_ _11430_ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_194_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Left_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17242_ rbzero.pov.spi_buffer\[14\] _10587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_241_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14454_ _08257_ _08259_ _08261_ _08255_ _08262_ _08263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__15933__A1 _09518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14736__A2 _07919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25996__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19785__I _12500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13405_ _07199_ _07216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_187_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17173_ _10532_ _10531_ _10534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14385_ _07185_ _08195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_153_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16124_ _09008_ _09657_ _09663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13336_ _07065_ _07150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_84_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16055_ rbzero.spi_registers.buf_texadd0\[4\] _09610_ _09611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13267_ _06865_ _07080_ _07081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15006_ _08805_ _08806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13172__A1 rbzero.spi_registers.texadd1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22431__A1 _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13198_ rbzero.spi_registers.texadd0\[19\] _07008_ _07011_ _07012_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_209_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19814_ _12585_ _12586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16110__A1 _08997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19745_ rbzero.wall_tracer.stepDistY\[-2\] _12256_ _12294_ _12517_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16957_ _08066_ _10182_ _10369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_155_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14672__A1 _08357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13475__A2 rbzero.spi_registers.vshift\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15908_ rbzero.spi_registers.buf_otherx\[1\] _09495_ _09500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19676_ _12275_ _12448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_79_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16888_ rbzero.debug_overlay.playerY\[-5\] _10303_ _10310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_220_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18627_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _11634_ _11635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_140_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15839_ _09442_ _09447_ _09448_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_188_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22498__A1 _12514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18558_ _11595_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18166__A2 _11308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17509_ _10779_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18489_ rbzero.tex_g1\[58\] rbzero.tex_g1\[57\] _11554_ _11556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20520_ _01611_ _01612_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14727__A2 _08248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_214_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20451_ _01446_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_144_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19666__A2 _11998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23170_ _03912_ _03957_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_20382_ _01473_ _01475_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_179_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22121_ _03088_ _03107_ _03112_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_242_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_22052_ rbzero.wall_tracer.stepDistY\[-1\] _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_58_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21003_ rbzero.wall_tracer.size_full\[9\] _01976_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26860_ _00770_ clknet_leaf_187_i_clk rbzero.tex_r0\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_195_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25811_ _06593_ _06594_ _06595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_215_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25911__A2 _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26791_ _00701_ clknet_leaf_197_i_clk rbzero.tex_g1\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_214_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22725__A2 _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14663__B2 _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25742_ _06519_ _06525_ _06526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22954_ _01580_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_190_i_clk_I clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21905_ _02941_ _02942_ _02945_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_25673_ _06453_ _06339_ _06456_ _06457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_195_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14079__I _07608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22885_ _03706_ _03743_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13218__A2 _07026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24478__A2 _05216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25675__A1 _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27412_ _01317_ clknet_leaf_109_i_clk rbzero.wall_tracer.stepDistX\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_194_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24624_ _05407_ _05408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_214_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21836_ _02880_ _02881_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_211_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27343_ _01248_ clknet_leaf_36_i_clk rbzero.texu_hot\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24555_ _05327_ _05338_ _05339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_93_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21767_ _02812_ _02814_ _02818_ _09953_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_194_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23506_ _04258_ _04261_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20718_ _01802_ _01808_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14718__A2 _08227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27274_ _01179_ clknet_leaf_46_i_clk rbzero.wall_tracer.texu\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24486_ _05207_ _05219_ _05229_ _05270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_21698_ _11307_ _02729_ _02759_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26225_ _00135_ clknet_leaf_6_i_clk rbzero.spi_registers.texadd1\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23437_ _04182_ _04290_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20649_ _01739_ _01652_ _01740_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_22_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_19__f_i_clk clknet_3_4_0_i_clk clknet_5_19__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_26156_ _00066_ clknet_leaf_218_i_clk rbzero.map_overlay.i_mapdy\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14170_ _07203_ _07790_ _07979_ _07980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23368_ _03714_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13941__A3 rbzero.map_overlay.i_mapdy\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25107_ _05301_ _05889_ _05890_ _05891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13121_ rbzero.side_hot _06933_ _06935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22319_ _11163_ _03270_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26087_ _05022_ _06811_ _06837_ _06852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__16340__A1 _08915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23299_ _04038_ _04152_ _04153_ _04043_ _04036_ _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__23855__I _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25038_ _05755_ _05818_ _05821_ _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_13052_ _06868_ _06869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17860_ rbzero.wall_tracer.rayAddendX\[4\] _11004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17840__A1 _10857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16811_ _10236_ _10237_ _10242_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_109_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16469__I _09925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17791_ _10951_ _10704_ _10954_ _10957_ _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_26989_ _00899_ clknet_leaf_131_i_clk rbzero.tex_g0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13457__A2 rbzero.spi_registers.vshift\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19530_ rbzero.wall_tracer.visualWallDist\[-11\] _12301_ _12302_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13954_ _07764_ _07765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16742_ _10181_ _10182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__20727__A1 _12885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16673_ _10073_ _10089_ _08096_ _10118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_89_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19461_ _07701_ _11098_ _12233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_198_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13885_ _07213_ _07693_ _07677_ _07102_ _07695_ _07696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_88_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18412_ _11501_ _11512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_202_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15624_ rbzero.spi_registers.texadd1\[20\] _09279_ _09287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_189_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19392_ _07237_ _07239_ _12164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14957__A2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15555_ _09234_ _09235_ _09229_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18343_ _11445_ _11470_ _11444_ _11471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__25418__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13621__I rbzero.row_render.side vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14506_ _07329_ _08315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18274_ _11413_ _11415_ _11416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15906__A1 _08946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15486_ rbzero.spi_registers.buf_texadd0\[8\] _09178_ _09185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13917__B1 _07721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14437_ _08240_ _08242_ _08244_ _07463_ _08245_ _08246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_17225_ rbzero.pov.spi_buffer\[10\] _10568_ _10565_ _10575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput11 net85 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15382__A2 _09108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput22 i_reg_sclk net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17156_ _10515_ _10520_ _10521_ _10522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13777__B _07587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14368_ _08173_ _08174_ _08177_ _08178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_123_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16107_ _08994_ _09646_ _09650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18320__A2 _11449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13319_ rbzero.spi_registers.texadd2\[1\] _07036_ _07133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17087_ rbzero.pov.ready_buffer\[17\] _10460_ _10470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14299_ rbzero.debug_overlay.vplaneY\[-5\] _08109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_122_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24370__B _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16038_ rbzero.spi_registers.buf_texadd0\[0\] _09597_ _09598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22404__A1 rbzero.wall_tracer.texu\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19820__A2 _12160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24157__A1 _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16379__I _08932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17989_ _11132_ _11133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14645__A1 _07841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15283__I _09035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23904__A1 _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19728_ _12499_ _12245_ _12331_ _12332_ _12500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__23714__B _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19659_ _12402_ _12431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_189_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_175_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22670_ rbzero.wall_tracer.trackDistX\[-9\] _03533_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14948__A2 _07101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21621_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] _02700_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_177_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_158_Right_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24340_ _04953_ _05090_ _05123_ _05124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__17898__A1 rbzero.debug_overlay.facingX\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21552_ _02632_ _02636_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20503_ _01590_ _01595_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__17938__I _11081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24271_ _05026_ _05054_ _05005_ _05020_ _05055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_118_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16570__A1 _09998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21483_ _02308_ _02567_ _02568_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_137_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26010_ _06786_ _06670_ _06666_ _06787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23222_ _03935_ _03955_ _04077_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13384__A1 _07189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20434_ _12912_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21446__A2 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23153_ rbzero.wall_tracer.stepDistX\[6\] _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20365_ _01387_ _01393_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22104_ _12185_ _03093_ _03094_ _03097_ _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_113_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20296_ _01389_ _01390_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_23084_ _02262_ _03817_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_227_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_244_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22035_ rbzero.wall_tracer.stepDistY\[-6\] _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26912_ _00822_ clknet_leaf_134_i_clk rbzero.tex_r1\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_228_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26843_ _00753_ clknet_leaf_196_i_clk rbzero.tex_r0\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13439__A2 _06859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25896__A1 _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20709__A1 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26774_ _00684_ clknet_leaf_197_i_clk rbzero.tex_g1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23986_ _04777_ _04778_ _04767_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_199_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23624__B _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14030__C _07839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25725_ _06508_ _06509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_242_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_205_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22937_ _03656_ _02349_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_196_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16389__A1 rbzero.spi_registers.spi_buffer\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15921__I _09494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25656_ _05333_ _06000_ _06440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_13670_ _07321_ _07338_ _07481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22868_ _12960_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24607_ _05376_ _05390_ _05391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_211_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21819_ _02856_ _02858_ _02864_ _02866_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_25587_ _06321_ _06370_ _06371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__14537__I _07551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22799_ _03655_ _03657_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_27326_ _01231_ clknet_leaf_117_i_clk rbzero.traced_texa\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15340_ rbzero.spi_registers.buf_mapdy\[2\] _09078_ _09079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24538_ _05320_ _05321_ _05322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27257_ _01162_ clknet_leaf_94_i_clk rbzero.wall_tracer.visualWallDist\[-3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_15271_ rbzero.map_overlay.i_otherx\[3\] _09019_ _09025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24469_ _05252_ _05196_ _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_149_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15364__A2 _09095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17010_ _10378_ _10412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26208_ _00118_ clknet_leaf_9_i_clk rbzero.spi_registers.texadd0\[23\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14222_ _07985_ _07990_ _07993_ _08032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__22634__A1 _09944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21437__A2 _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18689__I0 rbzero.tex_r1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27188_ _01093_ clknet_leaf_77_i_clk rbzero.wall_tracer.size\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_145_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14153_ _07432_ _07473_ _07440_ _07434_ _07963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_26139_ _00049_ clknet_leaf_215_i_clk rbzero.map_overlay.i_otherx\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13104_ _06917_ _06918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14084_ _07831_ _07894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18961_ _11852_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16864__A2 _08048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17912_ _08087_ rbzero.wall_tracer.rayAddendX\[3\] _11056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_18892_ rbzero.traced_texa\[5\] _07279_ _11806_ _11807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17843_ rbzero.pov.ready_buffer\[73\] _10852_ _10991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_206_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17774_ _10946_ _10947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14986_ _07246_ _08785_ _08787_ _08788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_19513_ _12276_ _12284_ _12285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16725_ _10161_ _10166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13937_ _07741_ _07678_ _07423_ _07743_ _07747_ _07748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_198_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17041__A2 _10434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19444_ rbzero.wall_tracer.rayAddendX\[-2\] _12216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_16656_ _10097_ _10098_ _10101_ _10102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_157_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13868_ _07244_ _07676_ _07677_ _07678_ _07679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_157_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24311__A1 _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15607_ rbzero.spi_registers.buf_texadd1\[15\] _09270_ _09275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19375_ rbzero.tex_b1\[62\] rbzero.tex_b1\[61\] _12151_ _12153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16587_ _10031_ _09977_ _10035_ _10036_ _10037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_146_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13799_ rbzero.tex_r0\[11\] _07584_ _07610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24365__B _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18326_ _11456_ _11458_ _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15538_ _09222_ _09223_ _09217_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__26064__A1 _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14891__B _08214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_211_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17758__I _10843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15469_ _07119_ _09124_ _09172_ _09126_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_18257_ rbzero.wall_tracer.mapX\[6\] _11400_ _11401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17208_ rbzero.pov.spi_buffer\[6\] _10556_ _10552_ _10562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18188_ _11331_ _11332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15278__I _09030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17139_ _10506_ _10507_ _10508_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19906__C _12352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20150_ _12902_ _12903_ _12921_ _12922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__14115__C _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14866__A1 _08321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22928__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20081_ _12847_ _12851_ _12852_ _12853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_185_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23050__A1 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_185_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21987__I0 rbzero.wall_tracer.rcp_fsm.o_data\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16607__A2 _10040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24320__S _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14618__A1 _07842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_227_Right_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23840_ _11143_ _03076_ _04670_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_222_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25215__I _05998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_63_i_clk_I clknet_5_21__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23771_ _04530_ _04609_ _04610_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_178_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20983_ _02071_ _01953_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13841__A2 _07459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15741__I _09352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25510_ _06159_ _06294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_178_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22722_ _02732_ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26490_ _00400_ clknet_leaf_48_i_clk rbzero.debug_overlay.facingX\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25441_ _06222_ _06224_ _06225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_177_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22653_ _11212_ _12214_ _03525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_149_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21604_ _10019_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25372_ _06153_ _06155_ _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22584_ _07234_ _03471_ _03472_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15897__B _09491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_27111_ _01021_ clknet_leaf_142_i_clk rbzero.tex_b1\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_91_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24323_ _04952_ _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_35_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21535_ _02506_ _02618_ _02619_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_145_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16543__A1 _09982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24605__A2 _05388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27042_ _00952_ clknet_leaf_159_i_clk rbzero.tex_g0\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_50_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24254_ _05037_ _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__21419__A2 _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21466_ _02545_ _02551_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_90_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_229_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23205_ _03946_ _03949_ _04060_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_105_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20417_ _12568_ _12644_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24185_ _04888_ _04944_ _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22092__A2 _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21397_ _02350_ _02353_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23136_ _03962_ _03992_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_219_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20348_ _01402_ _01442_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_242_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23067_ _03656_ _03792_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20279_ _12977_ _13032_ _01373_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__21978__I0 rbzero.wall_tracer.rcp_fsm.o_data\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_207_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22018_ _03033_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_216_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26826_ _00736_ clknet_leaf_176_i_clk rbzero.tex_g1\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14840_ rbzero.tex_b1\[22\] _07595_ _08646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_215_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14085__A2 _07894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14771_ _08335_ _08576_ _08577_ _08578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_23969_ _04764_ _04758_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26757_ _00667_ clknet_leaf_221_i_clk gpout0.vpos\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_86_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16747__I _09067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13832__A2 _07641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13372__S net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16510_ _09924_ _09963_ _09964_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13722_ rbzero.tex_r0\[35\] _07532_ _07533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18220__A1 _11344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25708_ _06037_ _05969_ _06453_ _06492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_168_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17490_ rbzero.tex_b0\[8\] rbzero.tex_b0\[7\] _10765_ _10769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_26688_ _00598_ clknet_leaf_26_i_clk rbzero.pov.ready_buffer\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16441_ _09897_ _09898_ _09899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13653_ _07332_ _07464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25639_ _06375_ _06421_ _06423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13171__I _06918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16782__A1 rbzero.debug_overlay.playerX\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19160_ _12003_ _12004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_155_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16372_ rbzero.spi_registers.buf_texadd3\[11\] _09840_ _09849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21658__A2 _08628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13584_ _07366_ rbzero.row_render.size\[0\] _07039_ _07395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15323_ _09064_ _09065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18111_ rbzero.map_rom.b6 _11255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_27309_ _01214_ clknet_leaf_112_i_clk rbzero.traced_texa\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_152_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19091_ _11926_ _11933_ _11934_ _11935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_152_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16482__I _09938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17582__I0 rbzero.tex_b0\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18042_ _11171_ _11183_ _11185_ _11186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15254_ _09013_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13899__A2 _07706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14205_ _08001_ _08014_ _08015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_111_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15185_ rbzero.spi_registers.spi_buffer\[10\] _08959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_10_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20094__A1 _12775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14136_ _07488_ _07946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_39_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19993_ _12456_ _12534_ _12393_ _12765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__14848__A1 _07889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23032__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18944_ _11842_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14067_ rbzero.tex_r1\[2\] _07876_ _07877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19787__A1 _12471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13520__A1 _07305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18875_ _11791_ _11792_ _11794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_193_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21594__A1 _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17826_ _10856_ _10980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_146_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14886__B _08603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17757_ _10934_ _10935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14969_ _08766_ _08769_ _08770_ _08771_ _08747_ _08772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__13823__A2 _07633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15561__I _08931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19033__I _11892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16708_ rbzero.wall_tracer.rayAddendY\[10\] _10150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17688_ _10874_ _10890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19427_ _12198_ _12199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_187_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23099__A1 _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16639_ _09897_ _09971_ _10086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13081__I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22608__B _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19358_ _12143_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23894__I0 rbzero.wall_tracer.rcp_fsm.o_data\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16606__B _09899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18309_ _07181_ _08753_ _11446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15510__B _09202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19289_ _12093_ _12104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_127_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21320_ _02259_ _02263_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21251_ _02071_ _02336_ _02192_ _02337_ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_187_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20202_ _12970_ _12972_ _12973_ _12974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_21182_ _02152_ _02153_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_40_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_245_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_224_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20133_ _12386_ _12587_ _12905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25990_ _06768_ _06769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_229_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20064_ _12835_ _12836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24941_ _05641_ _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24872_ _05654_ _05655_ _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14067__A2 _07876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24523__A1 _05304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24374__I1 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23823_ _04654_ _04655_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26611_ _00521_ clknet_leaf_170_i_clk rbzero.tex_b0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_213_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21337__A1 _12522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16567__I _09938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_202_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18202__A1 _11331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26542_ _00452_ clknet_leaf_24_i_clk rbzero.pov.spi_buffer\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_240_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23754_ _04592_ _04593_ _04595_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19250__I0 rbzero.tex_b1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_239_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15016__A1 _08811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20966_ _01988_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_198_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_239_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22705_ _11220_ rbzero.wall_tracer.stepDistX\[-5\] _03565_ _03571_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19950__A1 _12432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26473_ _00383_ clknet_leaf_206_i_clk rbzero.debug_overlay.playerY\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23685_ _04526_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20897_ _01961_ _01986_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_32_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_1_i_clk clknet_5_1__leaf_i_clk clknet_leaf_1_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25424_ _06008_ _06016_ _06004_ _06208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_22636_ _03493_ _03510_ _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_210_i_clk clknet_5_7__leaf_i_clk clknet_leaf_210_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_81_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25355_ _06138_ _06100_ _06139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22567_ _03463_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24306_ _05062_ _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21518_ _02601_ _02602_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25286_ _06066_ _06069_ _06070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_146_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__26803__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22498_ _12514_ _03417_ _03418_ _07378_ _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_27025_ _00935_ clknet_leaf_132_i_clk rbzero.tex_g0\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24237_ _05020_ _05021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_225_i_clk clknet_5_2__leaf_i_clk clknet_leaf_225_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_21449_ _02528_ _02534_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20076__A1 _12841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24168_ _04943_ _04945_ _04951_ _04929_ _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_112_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23119_ _03867_ _03873_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_112_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24099_ rbzero.wall_tracer.rcp_fsm.operand\[9\] _04846_ _04847_ _04883_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_16990_ _10396_ _10397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_247_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15941_ rbzero.spi_registers.spi_buffer\[4\] _09525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18660_ rbzero.tex_r1\[3\] rbzero.tex_r1\[2\] _11651_ _11654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_216_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15872_ _09429_ _09473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17611_ _10837_ _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_243_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26809_ _00719_ clknet_leaf_179_i_clk rbzero.tex_g1\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14823_ _08629_ net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_153_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18591_ _11614_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_231_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13805__A2 _07592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17542_ _10798_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14754_ rbzero.tex_b0\[29\] _08554_ _07955_ _08561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_230_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13705_ rbzero.tex_r0\[56\] _07515_ _07492_ _07516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17473_ _10758_ _10759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14685_ _07186_ _08491_ _08492_ net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_19212_ rbzero.wall_tracer.mapY\[8\] _12054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16424_ _09443_ _09887_ _09888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13636_ _07435_ _07446_ _07447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_172_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25490__A2 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19143_ _11939_ _11958_ _11987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16507__A1 _09945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14725__I _07935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16355_ _08939_ _09831_ _09837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13567_ rbzero.row_render.size\[6\] _07378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_137_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15306_ _07741_ _09043_ _09052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19074_ _08151_ rbzero.wall_tracer.rayAddendY\[7\] _11918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_11_i_clk_I clknet_5_4__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16286_ rbzero.spi_registers.buf_texadd2\[13\] _09780_ _09785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13498_ _07306_ _07308_ _07309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17180__A1 rbzero.pov.mosi vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18025_ rbzero.wall_tracer.trackDistX\[0\] _11169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15237_ _08951_ _09001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20067__A1 _12667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15168_ _08944_ _08940_ _08945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13785__B _07462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14119_ rbzero.tex_r1\[48\] _07629_ _07929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23005__A1 _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19976_ _12747_ _12740_ _12748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_165_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15099_ rbzero.spi_registers.spi_counter\[0\] _08889_ _08890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_182_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18927_ rbzero.tex_g0\[3\] rbzero.tex_g0\[2\] _11830_ _11833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21567__A1 _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_236_i_clk_I clknet_5_6__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18858_ _11737_ _11779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14049__A2 _07591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17809_ _10965_ _10723_ _10968_ _10969_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_238_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18789_ rbzero.tex_r1\[59\] rbzero.tex_r1\[58\] _11724_ _11727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15291__I _08987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20820_ _01798_ _01853_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_194_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20751_ _12173_ _01841_ _01525_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15549__A2 _09230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16746__A1 rbzero.pov.ready_buffer\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23470_ _04173_ _04174_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_174_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20682_ _01558_ _01658_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__25481__A2 _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_217_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22421_ _01776_ _03353_ _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_234_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25140_ _05896_ _05923_ _05924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22352_ _11278_ _03290_ _03299_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_21303_ _02384_ _02389_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_171_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25071_ _05794_ _05795_ _05582_ _05855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22283_ _11175_ _03245_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19999__A1 _12761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24022_ _04768_ _04805_ _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_103_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21234_ _02320_ _02264_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Left_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_229_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21165_ _02139_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_20116_ _12886_ _12623_ _12887_ _12888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25973_ _06749_ _06752_ _06704_ _06753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_217_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_21096_ _02084_ _02104_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_233_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20047_ _12815_ _12818_ _12819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24924_ _05707_ _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_176_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16297__I _09746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24855_ _05267_ _05639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_217_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23806_ _11161_ _03065_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24786_ _05407_ _05254_ _05570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_21998_ rbzero.wall_tracer.rcp_fsm.o_data\[6\] _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_157_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14460__A2 _07816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19923__A1 _12689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23737_ _11226_ _04554_ _04580_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26525_ _00435_ clknet_leaf_39_i_clk rbzero.pov.spi_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20949_ _01901_ _02028_ _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19401__I _12172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14470_ _07835_ _08279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23668_ rbzero.wall_tracer.stepDistX\[10\] _04519_ _11134_ _04520_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26456_ _00366_ clknet_leaf_206_i_clk rbzero.debug_overlay.playerX\[-3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_181_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13421_ _07231_ _07232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_25407_ _06075_ _06001_ _06189_ _06191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_12_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22619_ rbzero.wall_tracer.texu\[0\] rbzero.texu_hot\[0\] _03476_ _03501_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22286__A2 _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26387_ _00297_ clknet_leaf_14_i_clk rbzero.spi_registers.buf_texadd2\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23599_ _04449_ _04450_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23858__I _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19151__A2 rbzero.wall_tracer.rayAddendY\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20297__A1 _12210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16140_ _09675_ _09676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25338_ _06091_ _06120_ _06121_ _06122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13352_ gpout0.vinf _07164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_164_i_clk clknet_5_10__leaf_i_clk clknet_leaf_164_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_107_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_185_i_clk_I clknet_5_3__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16071_ rbzero.spi_registers.buf_texadd0\[8\] _09622_ _09623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25269_ _06049_ _06052_ _06053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13283_ _07095_ _07096_ _07097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15022_ _08817_ _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27008_ _00918_ clknet_leaf_190_i_clk rbzero.tex_g0\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_121_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21797__A1 rbzero.debug_overlay.vplaneX\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19830_ _12546_ _12566_ _12601_ _12602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xclkbuf_leaf_179_i_clk clknet_5_8__leaf_i_clk clknet_leaf_179_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19761_ _12508_ _12510_ _12532_ _12533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_16973_ _10378_ _10383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21549__A1 _12728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_235_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18712_ _11683_ _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15924_ _09511_ _09512_ _09505_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_223_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19692_ _12462_ _12463_ _12464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_102_i_clk clknet_5_27__leaf_i_clk clknet_leaf_102_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_30_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 i_gpout1_sel[1] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_160_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18643_ _11643_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15855_ _09459_ _09460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_231_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20772__A2 _12261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25160__A1 _05871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14806_ _07888_ _08581_ _08612_ _08357_ _08613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_18574_ _11604_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_125_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__18178__B1 _11106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15786_ rbzero.spi_registers.texadd3\[13\] _09407_ _09408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21841__I _09989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14451__A2 _07818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_117_i_clk clknet_5_19__leaf_i_clk clknet_leaf_117_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17525_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _10786_ _10789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14737_ rbzero.tex_b0\[37\] _08526_ _08543_ _08544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_197_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14883__C _08334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17456_ rbzero.pov.spi_buffer\[69\] _10743_ _10740_ _10747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_200_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14668_ _08472_ _08473_ _08475_ _07955_ _07913_ _08476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_52_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17940__A3 _11078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16407_ rbzero.spi_registers.buf_texadd3\[20\] _09874_ _09875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13619_ rbzero.floor_leak\[5\] _07326_ _07352_ _07429_ _07430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__14455__I _07479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17387_ rbzero.pov.spi_buffer\[51\] _10695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14599_ rbzero.tex_g1\[9\] _07857_ _07646_ _08407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19126_ _08161_ _10038_ _11970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16338_ _09823_ _09824_ _09822_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19057_ _11906_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15703__A2 _09338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16269_ _09761_ _09773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18008_ _11147_ rbzero.wall_tracer.trackDistY\[8\] _11152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15286__I _09037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19959_ _12729_ _12730_ _12731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_227_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_145_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22970_ _03822_ _03827_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__20141__B _12912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21921_ _02952_ _02696_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_241_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21960__A1 rbzero.wall_tracer.size\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24640_ _05422_ _05423_ _05424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_171_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21852_ _02883_ _02884_ _02882_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_65_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18169__B1 rbzero.map_rom.i_row\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19905__A1 _12675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14442__A2 _08250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20803_ _01893_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_195_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24571_ _05351_ _05352_ _05354_ _05355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_78_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21783_ _02829_ _02832_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16845__I _10271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26310_ _00220_ clknet_leaf_235_i_clk rbzero.spi_registers.buf_vshift\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23522_ _04291_ _04297_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20734_ _12569_ _01436_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27290_ _01195_ clknet_leaf_205_i_clk rbzero.row_render.side vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_175_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_81_i_clk clknet_5_28__leaf_i_clk clknet_leaf_81_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26241_ _00151_ clknet_leaf_21_i_clk rbzero.spi_registers.texadd2\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_232_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23453_ _04170_ _04187_ _04306_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_175_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20665_ _12472_ _01377_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23678__I _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22404_ rbzero.wall_tracer.texu\[0\] _03323_ _03348_ _03349_ _03350_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_26172_ _00082_ clknet_leaf_223_i_clk rbzero.color_sky\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23384_ _04237_ _04238_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17144__A1 _10067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20596_ _01590_ _01595_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25123_ _05873_ _05906_ _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22335_ _03287_ _03275_ _03288_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18892__A1 rbzero.traced_texa\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20294__A4 _12700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_96_i_clk clknet_5_26__leaf_i_clk clknet_leaf_96_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Left_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25054_ _05782_ _05790_ _05837_ _05838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_143_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22266_ _03231_ _03221_ _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21779__A1 rbzero.debug_overlay.vplaneX\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15196__I rbzero.spi_registers.spi_buffer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24005_ rbzero.wall_tracer.rcp_fsm.operand\[9\] _04722_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13709__I _07335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21217_ _02303_ _02304_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_218_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22197_ _03162_ _03164_ _03174_ _03109_ rbzero.wall_tracer.rcp_fsm.i_data\[5\] _03175_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__22440__A2 _07701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_247_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21148_ _02234_ _02235_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__20830__I _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25956_ _05033_ _06737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13970_ _07227_ _06874_ _07780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21079_ rbzero.traced_texVinit\[6\] _01551_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24907_ _05689_ _05690_ _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15145__B _08887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16958__A1 rbzero.pov.ready_buffer\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25887_ _06643_ _06668_ _06669_ _06670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__20754__A2 _12206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_61_Left_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_34_i_clk clknet_5_22__leaf_i_clk clknet_leaf_34_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_241_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_197_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15640_ rbzero.spi_registers.texadd2\[0\] _09291_ _09299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24838_ _05417_ _05426_ _05622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_17_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25693__A2 _06440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15571_ rbzero.spi_registers.buf_texadd1\[6\] _09245_ _09248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24769_ _05509_ _05551_ _05552_ _05553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__21703__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17310_ _10602_ _10638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14522_ _08321_ _08329_ _08330_ _08331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_26508_ _00418_ clknet_leaf_30_i_clk rbzero.debug_overlay.vplaneX\[-3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_18290_ rbzero.wall_tracer.mapX\[10\] _11424_ _11430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_49_i_clk clknet_5_17__leaf_i_clk clknet_leaf_49_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17241_ _10585_ _10583_ _10586_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26439_ _00349_ clknet_leaf_55_i_clk rbzero.wall_tracer.rayAddendY\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14275__I rbzero.debug_overlay.facingX\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14453_ _07333_ _08262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_83_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13404_ gpout0.vpos\[9\] gpout0.vpos\[8\] _07214_ _07215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__13944__A1 _07214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14384_ _07222_ _07973_ _08193_ _08194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_52_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17172_ _10532_ _10531_ _10533_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22492__I _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17135__A1 _10024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13112__C _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16123_ rbzero.spi_registers.buf_texadd0\[21\] _09655_ _09662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13335_ _07148_ _07149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_106_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18883__A1 rbzero.traced_texa\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21219__B1 _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23759__A2 _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24956__A1 _05696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16054_ _09596_ _09610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13266_ _07078_ _07079_ _07080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_51_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22967__B1 _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15005_ _06896_ _08805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_13197_ _07003_ _07010_ _07011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19813_ _12584_ _12585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_236_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25381__A1 _05948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24184__A2 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19744_ _12252_ _12513_ _12515_ _12516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14878__C _08346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__18210__I _11256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16956_ _10166_ _10366_ _10314_ _10368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__22195__A1 _11283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14672__A2 _08430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23931__A2 _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15907_ _09496_ _09499_ _09491_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19675_ _12437_ _12443_ _12446_ _12447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_205_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16949__A1 rbzero.pov.ready_buffer\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16887_ _10271_ _10309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__20745__A2 _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18626_ _11628_ _11634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_140_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15838_ _09429_ _09448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_140_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18557_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _11592_ _11595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15769_ _09393_ _09394_ _09395_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_177_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17508_ rbzero.tex_b0\[16\] rbzero.tex_b0\[15\] _10775_ _10779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18488_ _11555_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_185_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23447__A1 _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17439_ rbzero.pov.spi_buffer\[64\] _10734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_214_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_214_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20450_ _01462_ _01464_ _01543_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_28_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17126__A1 rbzero.pov.ready_buffer\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19109_ _11952_ _11953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_127_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20381_ _12969_ _01474_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_242_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22670__A2 _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22120_ rbzero.wall_tracer.rcp_fsm.i_data\[-9\] _03109_ _03111_ _03112_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22051_ _03057_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_58_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21002_ _01528_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25810_ _06578_ _06587_ _06594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26790_ _00700_ clknet_leaf_129_i_clk rbzero.tex_g1\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_71_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input28_I i_vec_mosi vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_133_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25741_ _06520_ _06524_ _06525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22953_ _02262_ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21904_ _02941_ _02942_ _02945_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_223_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25672_ _06389_ _06454_ _06455_ _06456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22884_ _03708_ _03742_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27411_ _01316_ clknet_leaf_107_i_clk rbzero.wall_tracer.stepDistX\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24623_ _05219_ _05407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21835_ rbzero.debug_overlay.vplaneX\[-1\] _08131_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_214_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24554_ _05330_ _05333_ _05336_ _05337_ _05338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27342_ _01247_ clknet_leaf_37_i_clk rbzero.texu_hot\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21766_ _08143_ _12185_ _02817_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_182_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23505_ _04252_ _04356_ _04357_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20717_ _01806_ _01807_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_135_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24485_ _05268_ _05269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_27273_ _01178_ clknet_leaf_93_i_clk rbzero.wall_tracer.side vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21697_ _12046_ _02758_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23989__A2 _08814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26224_ _00134_ clknet_leaf_6_i_clk rbzero.spi_registers.texadd1\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23436_ _04181_ _04184_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20648_ _01629_ _01639_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_78_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_78_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26155_ _00065_ clknet_leaf_218_i_clk rbzero.map_overlay.i_mapdy\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_190_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23367_ _03736_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18865__A1 _11779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20579_ _01646_ _01651_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_58_i_clk_I clknet_5_23__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13120_ rbzero.side_hot _06933_ _06934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25106_ _05311_ _05890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_22318_ _03220_ _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__20672__A1 _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26086_ _06811_ _06812_ _06850_ _06691_ _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23298_ _03922_ _04042_ _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25037_ _05819_ _05820_ _05821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13051_ _06867_ _06868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_22249_ _03209_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19554__C _12325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16810_ rbzero.pov.ready_buffer\[68\] _10228_ _10229_ _10241_ _10242_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__25363__A1 _06003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17790_ _10952_ rbzero.pov.ready_buffer\[54\] _10957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_109_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26988_ _00898_ clknet_leaf_146_i_clk rbzero.tex_g0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14654__A2 _07940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16741_ _10162_ _10181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25939_ _06696_ _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13953_ _07755_ _07759_ _07763_ _07764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__19593__A2 _12363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19460_ _12225_ _12227_ _12230_ _12231_ _12232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_89_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16672_ _10074_ _10090_ _10117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13884_ _07694_ _06874_ _07695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_89_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15603__A1 rbzero.spi_registers.texadd1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18411_ _11511_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_186_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15623_ _09285_ _09286_ _09278_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19391_ rbzero.trace_state\[2\] _12163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_201_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18342_ _07176_ _07779_ _11450_ _11470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_186_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15554_ rbzero.spi_registers.buf_texadd1\[2\] _09232_ _09235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25418__A2 _06102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14505_ _08264_ _08286_ _08296_ _08303_ _08313_ _08314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_18273_ _11403_ _11405_ _11414_ _11415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15906__A2 _09498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15485_ rbzero.spi_registers.texadd0\[8\] _09176_ _09184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__26091__A2 _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17224_ rbzero.pov.spi_buffer\[9\] _10574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_182_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14436_ _07333_ _08245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_24_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 i_gpout2_sel[0] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_226_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput23 i_reset net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_25_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17155_ _07167_ rbzero.pov.ss_buffer\[1\] _10521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22652__A2 _12395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14367_ _08175_ _08065_ _08060_ _08176_ _07218_ _08177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_24_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16106_ rbzero.spi_registers.buf_texadd0\[17\] _09644_ _09649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13318_ rbzero.spi_registers.texadd3\[1\] _07111_ _07030_ rbzero.spi_registers.texadd1\[1\]
+ _07132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_14298_ _08106_ _08039_ _08044_ _08107_ _08108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_17086_ _08143_ _10458_ _10469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_208_Right_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16037_ _09596_ _09597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13249_ _07062_ _07063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14893__A2 _07484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_199_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16095__A1 _08980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24157__A2 _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22168__A1 _11293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17988_ _11131_ _11132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_236_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19727_ rbzero.wall_tracer.stepDistX\[-7\] _12499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_16939_ _08057_ _10348_ _10354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13084__I _06898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19658_ _12429_ _12430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25657__A2 _06440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18609_ _11624_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16395__I _09855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19589_ _12360_ _12361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_177_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23668__A1 rbzero.wall_tracer.stepDistX\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_177_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21620_ _02695_ _02699_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__21143__A2 _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14129__B _07917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21551_ _02634_ _02635_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_20502_ _01593_ _01594_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_24270_ _05015_ _05051_ _05053_ _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_16_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21482_ rbzero.traced_texVinit\[9\] _01551_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24117__I _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23221_ _03938_ _03954_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_133_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15739__I _09349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20433_ rbzero.wall_tracer.size_full\[4\] _01430_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18847__A1 rbzero.traced_texa\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23956__I _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23152_ rbzero.wall_tracer.trackDistX\[6\] _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20364_ _01375_ _01395_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22103_ _09948_ _03095_ _03096_ _12834_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_23083_ _02258_ _03815_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20295_ _12971_ _12704_ _12688_ _12967_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_73_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22034_ _03030_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26911_ _00821_ clknet_leaf_134_i_clk rbzero.tex_r1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_244_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15474__I _09150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_209_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26842_ _00752_ clknet_leaf_190_i_clk rbzero.tex_r0\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13439__A3 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26773_ _00683_ clknet_leaf_197_i_clk rbzero.tex_g1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23985_ rbzero.wall_tracer.rcp_fsm.i_data\[3\] _04770_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21906__A1 _10121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25724_ _06472_ _06507_ _06508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22936_ _03654_ _02481_ _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_104_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25655_ _06436_ _06437_ _06438_ _06439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__22100__I _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25112__A4 _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22867_ _03725_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24606_ _05378_ _05379_ _05390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_168_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13072__A1 _06884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21818_ _10015_ _02865_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25586_ _06322_ _06369_ _06370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22798_ _03656_ _02481_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_195_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22331__A1 _11283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13611__A3 _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27325_ _01230_ clknet_leaf_115_i_clk rbzero.traced_texa\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24537_ _05273_ _05321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21749_ _02708_ _02801_ _02802_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_182_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20893__A1 _12836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27256_ _01161_ clknet_leaf_90_i_clk rbzero.wall_tracer.visualWallDist\[-4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_15270_ _09023_ _09024_ _09018_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24468_ _05238_ _05251_ _05252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26207_ _00117_ clknet_leaf_239_i_clk rbzero.spi_registers.texadd0\[22\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14221_ _08030_ _08031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_23419_ _04162_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_27187_ _01092_ clknet_leaf_77_i_clk rbzero.wall_tracer.size\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24399_ _05121_ _04910_ _05131_ _05130_ _05060_ _05079_ _05183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__18689__I1 rbzero.tex_r1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14152_ _07458_ _07447_ _07455_ _07436_ _07962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_26138_ _00048_ clknet_leaf_218_i_clk rbzero.map_overlay.i_otherx\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19565__B _12310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_28__f_i_clk_I clknet_3_7_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13103_ _06916_ _06917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14083_ rbzero.tex_r1\[33\] _07635_ _07893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18960_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _11851_ _11852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26069_ _06777_ _06837_ _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_219_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17911_ _11045_ _11053_ _11054_ _11055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14875__A2 _08250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18891_ _11803_ _11805_ _11806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16077__A1 _08962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17842_ rbzero.pov.spi_buffer\[73\] _10990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_234_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17773_ _09034_ _10946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14985_ _07178_ _08786_ _07712_ _07191_ _08787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_19512_ _12283_ _12284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16724_ _10164_ _10165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13936_ _07737_ _07373_ _07678_ _07741_ _07746_ _07747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__22570__A1 _11281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19443_ rbzero.wall_tracer.size_full\[-10\] _12173_ _12215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22570__B2 rbzero.traced_texa\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16655_ _10099_ _10100_ _10101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13867_ _07101_ _07678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_157_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15606_ rbzero.spi_registers.texadd1\[15\] _09268_ _09274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19374_ _12152_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_232_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16586_ _09973_ _10036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22322__A1 _11290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13798_ _07608_ _07609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18325_ _11432_ _11457_ _11458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15537_ rbzero.spi_registers.buf_texadd0\[21\] _09220_ _09223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__26064__A2 rbzero.wall_tracer.rcp_fsm.o_data\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_211_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18256_ _11399_ _11400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_15468_ rbzero.spi_registers.buf_texadd0\[3\] _09137_ _09172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_154_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17207_ rbzero.pov.spi_buffer\[5\] _10561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_135_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14419_ rbzero.tex_g0\[20\] _08227_ _08220_ _08228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18187_ rbzero.map_rom.f4 _11331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15399_ rbzero.color_sky\[2\] _09115_ _09122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17138_ _10491_ _10508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_90_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13079__I _06894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17069_ _10455_ _10432_ _10456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22389__A1 _12907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20080_ _12845_ _12846_ _12852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_0_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16068__A1 _08950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14412__B _08220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21987__I1 rbzero.wall_tracer.size\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_191_Right_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25878__A2 _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23889__A1 _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_222_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_222_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19557__A2 _11078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23770_ _04605_ _04608_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_178_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20982_ _12464_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_192_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22721_ _11173_ _12511_ _03584_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_149_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25440_ _06220_ _06223_ _06224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22652_ rbzero.wall_tracer.trackDistX\[-11\] _12395_ _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22855__I _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22313__A1 _11165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16791__A2 _10224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21603_ _02571_ _02687_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_168_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25371_ _06154_ _05998_ _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_22583_ rbzero.wall_tracer.w\[2\] rbzero.wall_tracer.w\[1\] rbzero.wall_tracer.w\[0\]
+ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_76_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27110_ _01020_ clknet_leaf_142_i_clk rbzero.tex_b1\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24322_ _04987_ _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_21534_ _02508_ _02513_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20375__I _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24253_ _05012_ _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_27041_ _00951_ clknet_leaf_159_i_clk rbzero.tex_g0\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21465_ _02549_ _02550_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22616__A2 _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23686__I _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23204_ _02271_ _04059_ _03947_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_20416_ _12494_ _12585_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19493__A1 _12261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24184_ _04920_ _04921_ _04901_ _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__18296__A2 _07707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21396_ _02481_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_160_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23135_ _03964_ _03991_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_247_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20347_ _01404_ _01441_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_105_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23066_ _03654_ _03652_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20278_ _12979_ _13031_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_235_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21978__I1 _12514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22017_ _03029_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14609__A2 _07579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25869__A2 _06628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26825_ _00735_ clknet_leaf_178_i_clk rbzero.tex_g1\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_242_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26756_ _00666_ clknet_leaf_222_i_clk gpout0.vpos\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14770_ rbzero.tex_b0\[18\] _08342_ _08577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13293__A1 _07065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23968_ rbzero.wall_tracer.rcp_fsm.operand\[0\] _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22552__A1 _11293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25707_ _06438_ _06489_ _06490_ _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_169_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13721_ _07531_ _07532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22919_ _03646_ _03675_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14548__I _07326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26687_ _00597_ clknet_leaf_26_i_clk rbzero.pov.ready_buffer\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23899_ _03893_ _04704_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16440_ _07241_ _08869_ _09898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25638_ _06375_ _06421_ _06422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_151_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13652_ _07462_ _07463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_168_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14242__B1 _08040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16371_ _09847_ _09848_ _09844_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25569_ _06280_ _06289_ _06353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_186_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13583_ rbzero.row_render.size\[5\] _07386_ _07394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18110_ rbzero.debug_overlay.playerX\[3\] _11249_ _11251_ rbzero.debug_overlay.playerY\[4\]
+ _11253_ _11254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_82_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27308_ _01213_ clknet_leaf_112_i_clk rbzero.traced_texa\[-10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15322_ _08877_ _09064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19090_ _08155_ _10030_ _11934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_152_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18041_ rbzero.wall_tracer.trackDistX\[2\] _11184_ _11167_ _11168_ _11185_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_136_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14545__A1 _08304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27239_ _01144_ clknet_leaf_92_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15253_ _08818_ net29 _09013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13401__B _06859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14204_ _08002_ _08013_ _08014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_152_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15184_ _08956_ _08958_ _08954_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_10_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16298__A1 _08990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20094__A2 _12864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14135_ rbzero.tex_r1\[62\] _07645_ _07945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19992_ _12757_ _12762_ _12763_ _12764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_120_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18943_ rbzero.tex_g0\[10\] rbzero.tex_g0\[9\] _11840_ _11842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14066_ _07511_ _07876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_167_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21043__A1 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18874_ _11791_ _11792_ _11793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_234_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17825_ _10848_ _10979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_33_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17756_ _10847_ _10934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14968_ _07180_ _08749_ _08760_ gpout0.vpos\[0\] _08756_ _07179_ _08771_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__13284__A1 _07050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16707_ _10072_ _10144_ _10148_ _10049_ _10149_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_89_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13919_ rbzero.map_overlay.i_otherx\[4\] _06868_ _07730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__18211__A2 _11308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17687_ _10872_ _10889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14899_ rbzero.tex_b1\[49\] _07577_ _08214_ _08705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19426_ _12197_ _12198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16638_ _10081_ _10084_ _10085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_231_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19357_ rbzero.tex_b1\[54\] rbzero.tex_b1\[53\] _12141_ _12143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16569_ _10008_ _10020_ _10021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23894__I1 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26037__A2 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18308_ _11444_ _08788_ _11445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_57_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_232_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_0__f_i_clk clknet_3_0_0_i_clk clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_99_Left_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_19288_ _12103_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18239_ _11382_ _11383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_170_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13311__B _07028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14536__A1 _08334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13339__A2 _07146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20609__A1 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14126__C _07935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21250_ _02190_ _02191_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_187_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23271__A2 _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20201_ _12933_ _12700_ _12973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21181_ _02148_ _02267_ _02268_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_20132_ _12525_ _12646_ _12904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_224_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24331__S _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14142__B _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20063_ _12834_ _12301_ _12835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24940_ _05640_ _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_24871_ _05418_ _05466_ _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16461__A1 _09895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26610_ _00520_ clknet_leaf_168_i_clk rbzero.tex_b0\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_213_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23822_ _03287_ _03069_ _04649_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_202_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_202_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26541_ _00451_ clknet_leaf_24_i_clk rbzero.pov.spi_buffer\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_240_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23753_ _04592_ _04593_ _04594_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18202__A2 _11343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20965_ _02052_ _02053_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_239_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15016__A2 _08814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_198_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_239_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22704_ _03570_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26472_ _00382_ clknet_leaf_207_i_clk rbzero.debug_overlay.playerY\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20896_ _01962_ _01985_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_23684_ _04524_ _04529_ _04534_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__17679__I _08809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25423_ _06193_ _06205_ _06206_ _06207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_119_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22635_ _03509_ _03510_ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25354_ _06063_ _06094_ _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24039__A1 _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22566_ _11283_ _03461_ _03462_ rbzero.traced_texa\[5\] _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19894__I _12369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15199__I _08933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24429__I3 _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21517_ _01948_ _02097_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24305_ _05088_ _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_106_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25285_ _06067_ _06068_ _06069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22497_ _03420_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_27024_ _00934_ clknet_leaf_132_i_clk rbzero.tex_g0\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_90_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24236_ _05019_ _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21448_ _02529_ _02533_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_146_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24167_ _04922_ _04948_ _04949_ _04950_ _04942_ _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_21379_ _02339_ _02346_ _02344_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23118_ _03973_ _03974_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_112_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24098_ _04881_ _04882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_101_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_236_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23049_ _03847_ _03855_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15940_ rbzero.spi_registers.buf_othery\[4\] _09494_ _09524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15871_ _08937_ _09459_ _09472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_204_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_216_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17610_ rbzero.tex_b0\[60\] rbzero.tex_b0\[59\] _10833_ _10837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16452__A1 rbzero.debug_overlay.vplaneY\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26808_ _00718_ clknet_leaf_179_i_clk rbzero.tex_g1\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14822_ reg_rgb\[4\] _08628_ _08195_ _08629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_18590_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _11613_ _11614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_181_i_clk_I clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17541_ rbzero.tex_b0\[30\] rbzero.tex_b0\[29\] _10796_ _10798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14753_ rbzero.tex_b0\[28\] _08494_ _08560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26739_ _00649_ clknet_leaf_40_i_clk rbzero.pov.ready_buffer\[69\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_230_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22709__B _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13704_ _07340_ _07515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17472_ _10757_ _10758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_196_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14684_ _08195_ reg_rgb\[3\] _08492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19211_ _12048_ _12049_ _12050_ _12053_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_168_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16423_ _09885_ _09887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13635_ rbzero.row_render.texu\[3\] rbzero.row_render.texu\[2\] rbzero.row_render.texu\[1\]
+ _07328_ _07445_ _07446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_156_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13910__I rbzero.map_overlay.i_othery\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19142_ _08152_ _10089_ _11975_ _11986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_15_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16354_ rbzero.spi_registers.buf_texadd3\[6\] _09829_ _09836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13566_ rbzero.row_render.size\[5\] _06884_ _07100_ _07363_ _07377_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_165_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15305_ _09050_ _09051_ _09042_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19073_ _08159_ rbzero.wall_tracer.rayAddendY\[8\] _11917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_54_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16285_ _09781_ _09783_ _09784_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13497_ _07307_ _07308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_132_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18024_ rbzero.wall_tracer.trackDistX\[1\] _11168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_152_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15236_ rbzero.spi_registers.spi_buffer\[19\] _09000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15191__A1 rbzero.spi_registers.spi_buffer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15167_ rbzero.spi_registers.spi_buffer\[7\] _08944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14118_ _07349_ _07928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_239_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19975_ _12682_ _12720_ _12747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15098_ _08856_ _08862_ _08867_ _08889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_120_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18926_ _11832_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14049_ rbzero.tex_r1\[11\] _07591_ _07859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_197_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I i_debug_trace_overlay vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21567__A2 _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18857_ _08750_ _08751_ _11774_ _11777_ _11778_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_235_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17808_ _10966_ rbzero.pov.ready_buffer\[60\] _10969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18788_ _11726_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13257__A1 _06906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22516__A1 rbzero.wall_tracer.texu\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17739_ _10921_ rbzero.pov.ready_buffer\[36\] _10924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13092__I _06905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20750_ _01840_ _01717_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_203_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16746__A2 _10183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19409_ _12180_ _12181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_20681_ _01561_ _01657_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22420_ _01892_ _03363_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_163_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_217_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19696__A1 _12369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_234_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14137__B _07946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22351_ _11142_ _03243_ _03301_ _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21302_ _02385_ _02388_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22354__B _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25070_ _05838_ _05853_ _05854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19448__A1 rbzero.wall_tracer.stepDistY\[-10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22282_ _03205_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23244__A2 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24021_ _04802_ _04803_ _04804_ _04794_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_21233_ _02255_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14651__I _07337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18120__A1 rbzero.debug_overlay.playerX\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21164_ _02249_ _02251_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20115_ _12471_ _12885_ _12562_ _12501_ _12887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__25941__A1 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25972_ _06702_ _06752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21095_ _02063_ _02083_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20046_ _12816_ _12817_ _12818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24923_ _05705_ _05706_ _05707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_99_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24854_ _05628_ _05603_ _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_213_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23805_ _11161_ _03065_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19889__I _12660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14996__A1 _07175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18793__I _11713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13799__A2 _07584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24785_ _05512_ _05515_ _05568_ _05569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_21997_ _03017_ _03011_ _03018_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19923__A2 _12691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26524_ _00434_ clknet_leaf_39_i_clk rbzero.pov.spi_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23736_ _04542_ _04579_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20948_ _01895_ _02031_ _02036_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_83_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21730__A2 _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26455_ _00365_ clknet_leaf_45_i_clk rbzero.debug_overlay.playerX\[-4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_23667_ _11140_ _04518_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20879_ _01723_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13730__I _07444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25406_ _06075_ _06001_ _06189_ _06190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13420_ _07223_ _07225_ _07230_ _07231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_181_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22618_ _03490_ _03499_ _03500_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_12_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19687__A1 _12425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26386_ _00296_ clknet_leaf_14_i_clk rbzero.spi_registers.buf_texadd2\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23598_ _04431_ _04439_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24463__C _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25337_ _06009_ _06089_ _06083_ _06121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__19151__A3 _11993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13351_ clknet_leaf_226_i_clk _07158_ net14 _07163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22549_ _03452_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_128_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15173__A1 _08948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16070_ _09596_ _09622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25268_ _06051_ _06033_ _06052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24035__I _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13282_ _06906_ _06970_ _07096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15021_ _08807_ rbzero.spi_registers.mosi_buffer\[0\] _08817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27007_ _00917_ clknet_leaf_200_i_clk rbzero.tex_g0\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24219_ _04932_ _04917_ _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__14920__A1 _08355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25199_ _05982_ _05983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18968__I _11850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13177__I _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14279__A3 _07719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19760_ _12530_ _12531_ _12532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16972_ _08084_ _10381_ _10382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21549__A2 _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15923_ _08965_ _09508_ _09512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18711_ rbzero.tex_r1\[25\] rbzero.tex_r1\[24\] _11682_ _11683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_19691_ _11388_ _12419_ _12463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16488__I _09896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15392__I _08882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20221__A2 _12258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18642_ rbzero.tex_r0\[60\] rbzero.tex_r0\[59\] _11639_ _11643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15854_ _09444_ _09458_ _09459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_232_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_231_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14805_ _08586_ _08594_ _08611_ _07478_ _08612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_204_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25160__A2 _05908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18573_ rbzero.tex_r0\[30\] rbzero.tex_r0\[29\] _11602_ _11604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15785_ _09037_ _09407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18178__A1 rbzero.map_overlay.i_otherx\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18178__B2 _09027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17524_ _10788_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14736_ rbzero.tex_b0\[36\] _07919_ _08543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_52_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17455_ _10712_ _10746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14667_ rbzero.tex_g1\[50\] _07919_ _08474_ _08475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_184_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16406_ _09814_ _09874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13618_ gpout0.vinf _07428_ _07429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_45_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17940__A4 _11083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13411__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17386_ _10692_ _10688_ _10694_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14598_ rbzero.tex_g1\[8\] _07855_ _08406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19125_ _11960_ _11967_ _11968_ _11969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_82_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16337_ _08913_ _09820_ _09824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13549_ _06883_ _07358_ _07359_ _07360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19056_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _11903_ _11906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16268_ _08948_ _09771_ _09772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18007_ rbzero.wall_tracer.trackDistY\[6\] _11151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_140_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15567__I _09208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15219_ _08986_ _08987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_164_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16199_ _09670_ _09719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22902__B _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22985__A1 _12760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_i_clk clknet_5_1__leaf_i_clk clknet_leaf_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_19958_ _12328_ _12730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_145_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18909_ _11779_ _11820_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19889_ _12660_ _12661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_241_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21920_ _10022_ _02954_ _02958_ _02960_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_207_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__26802__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21851_ _02895_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_222_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_224_i_clk clknet_5_2__leaf_i_clk clknet_leaf_224_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__18169__A1 rbzero.map_overlay.i_mapdy\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18169__B2 _07754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19502__I _12273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19905__A2 _12676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20802_ rbzero.traced_texVinit\[4\] _01778_ _01892_ _01662_ _01893_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_236_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24570_ _05353_ _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21782_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] _02831_
+ _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_195_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23521_ _04291_ _04297_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20733_ _12999_ _13024_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26240_ _00150_ clknet_leaf_14_i_clk rbzero.spi_registers.texadd2\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20664_ _12968_ _01468_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23452_ _04284_ _04186_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_239_i_clk clknet_5_1__leaf_i_clk clknet_leaf_239_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22403_ _03340_ _03345_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_23383_ _04016_ _04114_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26171_ _00081_ clknet_leaf_224_i_clk rbzero.color_sky\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20595_ _01587_ _01602_ _01677_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__18341__A1 _11462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25122_ _05877_ _05905_ _05906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_60_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22334_ _11156_ _03270_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22265_ rbzero.wall_tracer.trackDistX\[-6\] _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_170_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25053_ _05777_ _05781_ _05837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14902__B2 _08564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24004_ _04790_ _04791_ _04786_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_21216_ _02174_ _02302_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22196_ _03165_ _03173_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_247_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21147_ _12787_ _02111_ _02233_ _12192_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13469__A1 rbzero.traced_texVinit\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25955_ _06726_ _06735_ _05007_ _06736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_21078_ _02037_ _02040_ _02166_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_245_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20029_ _12786_ _12800_ _12801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24906_ _05286_ _05493_ _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25886_ _06631_ _06639_ _06669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_54_i_clk_I clknet_5_25__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24837_ _05611_ _05619_ _05620_ _05621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_17_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15570_ rbzero.spi_registers.texadd1\[6\] _09243_ _09247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24768_ _05511_ _05516_ _05552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_197_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14521_ rbzero.tex_g0\[50\] _07834_ _08330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26507_ _00417_ clknet_leaf_59_i_clk rbzero.debug_overlay.vplaneX\[-4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23719_ _11196_ _03046_ _04564_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_139_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24699_ _05481_ _05482_ _05483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17240_ rbzero.pov.spi_buffer\[14\] _10580_ _10577_ _10586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_120_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26438_ _00348_ clknet_leaf_55_i_clk rbzero.wall_tracer.rayAddendY\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14452_ rbzero.tex_g0\[14\] _08258_ _08260_ _08261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_187_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13403_ _07213_ _07214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17171_ _10532_ _10531_ _10521_ _10533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14383_ _08192_ _08193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26369_ _00279_ clknet_leaf_4_i_clk rbzero.spi_registers.buf_texadd1\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16122_ _09656_ _09658_ _09661_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13334_ _07060_ _07057_ _06905_ _07148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__24405__A1 _05186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18883__A2 rbzero.texV\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15697__A2 _09338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16053_ _09608_ _09609_ _09603_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16894__A1 rbzero.pov.ready_buffer\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21219__B2 _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13265_ _06886_ _07079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23818__B _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15004_ _08804_ _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22967__A1 _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22967__B2 _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13196_ rbzero.spi_registers.texadd3\[19\] _06997_ _07009_ rbzero.spi_registers.texadd2\[19\]
+ _06998_ rbzero.spi_registers.texadd1\[19\] _07010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_209_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19812_ _12574_ _12583_ _12584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19743_ _12514_ _12171_ _12515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14121__A2 _07930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16955_ _10365_ _10367_ _10214_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_223_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15906_ _08946_ _09498_ _09499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19674_ _12417_ _12418_ _12419_ _12445_ _12368_ _12446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_16886_ _10272_ _10308_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13880__A1 rbzero.debug_overlay.playerX\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_205_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_204_Left_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15837_ _08920_ _09446_ _09447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18625_ _11633_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_205_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18556_ _11594_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15768_ _09383_ _09395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_177_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23695__A2 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17507_ _10778_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14719_ _07537_ _08526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__24319__S1 _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18487_ rbzero.tex_g1\[57\] rbzero.tex_g1\[56\] _11554_ _11555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15699_ _09342_ _09343_ _09337_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17438_ _10731_ _10724_ _10733_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23447__A2 _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13303__C _07057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_214_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_214_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13935__A2 _06873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17369_ _10658_ _10682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_160_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19108_ _11948_ _11951_ _11952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15137__A1 _08915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_213_Left_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20380_ _12957_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19039_ _11896_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16885__A1 _08041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23728__B _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22050_ rbzero.wall_tracer.rcp_fsm.o_data\[-2\] _03056_ _03051_ _03057_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21001_ rbzero.wall_tracer.size_full\[9\] _01976_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_227_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21630__A1 _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24255__S0 _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14112__A2 _07919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25740_ _05979_ _06522_ _06523_ _06524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_242_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_222_Left_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22952_ _03800_ _03673_ _03809_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_163_i_clk clknet_5_10__leaf_i_clk clknet_leaf_163_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_3_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17062__A1 rbzero.pov.ready_buffer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21903_ _02906_ _02943_ _02944_ _02907_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_25671_ _05982_ _06013_ _06387_ _06455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_22883_ _03721_ _03724_ _03741_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_27410_ _01315_ clknet_leaf_107_i_clk rbzero.wall_tracer.stepDistX\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_214_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__19232__I _11478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24622_ _05384_ _05392_ _05405_ _05406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_21834_ _08125_ _08127_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27341_ _01246_ clknet_leaf_36_i_clk rbzero.texu_hot\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24553_ _05313_ _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_178_i_clk clknet_5_8__leaf_i_clk clknet_leaf_178_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_21765_ _08133_ rbzero.wall_tracer.rayAddendX\[-4\] _02816_ _02817_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23504_ _04342_ _04345_ _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_20716_ _12433_ _01803_ _01805_ _12426_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27272_ _01177_ clknet_leaf_204_i_clk rbzero.wall_tracer.wall\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24484_ _05206_ _05218_ _05228_ _05268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_19_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21696_ _07693_ _02733_ _02756_ _02757_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_93_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17687__I _10872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26223_ _00133_ clknet_leaf_6_i_clk rbzero.spi_registers.texadd1\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23435_ _04285_ _04288_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_46_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_231_Left_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_191_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20647_ _01640_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_101_i_clk clknet_5_27__leaf_i_clk clknet_leaf_101_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_22_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26154_ _00064_ clknet_leaf_218_i_clk rbzero.map_overlay.i_mapdy\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23366_ _04219_ _04220_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20578_ _01646_ _01651_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25105_ _05314_ _05889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16876__A1 _08042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22317_ _03201_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_5_18__f_i_clk_I clknet_3_4_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26085_ _06672_ _06787_ _06850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23297_ _04151_ _04040_ _04041_ _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_104_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25036_ _05636_ _05685_ _05820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13050_ _06866_ _06867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_22248_ _11207_ _03204_ _03216_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_116_i_clk clknet_5_19__leaf_i_clk clknet_leaf_116_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22179_ _11954_ _03095_ _03105_ _11291_ _03115_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_245_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_245_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26987_ _00897_ clknet_leaf_146_i_clk rbzero.tex_g0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_109_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_28__f_i_clk clknet_3_7_0_i_clk clknet_5_28__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__19578__B1 _12347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16740_ _10179_ _10180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25938_ _06694_ _02990_ _06661_ _06718_ _06719_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_13952_ _07684_ rbzero.map_overlay.i_mapdy\[4\] _07751_ _07760_ _07762_ _07763_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__21672__I _12035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16671_ _08096_ _10107_ _10116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_25869_ _06650_ _06628_ _06652_ _06653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_89_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13883_ rbzero.debug_overlay.playerX\[2\] _07694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_214_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15622_ rbzero.spi_registers.buf_texadd1\[19\] _09281_ _09286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18410_ rbzero.tex_g1\[24\] rbzero.tex_g1\[23\] _11507_ _11511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16800__A1 _07708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19390_ _12159_ _12162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__20288__I _12448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18341_ _11462_ _11468_ _11469_ _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_15553_ rbzero.spi_registers.texadd1\[2\] _09230_ _09234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14504_ _08304_ _08312_ _08313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_204_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18272_ _11407_ _11414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_166_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15484_ _06958_ _09180_ _09183_ _09182_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__20360__A1 _09901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16715__B _09934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17223_ _10570_ _10572_ _10573_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_155_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14435_ rbzero.tex_g0\[5\] _08241_ _08243_ _08244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13917__A2 rbzero.map_overlay.i_othery\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18305__A1 _07102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 i_gpout2_sel[1] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 i_tex_in[0] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17154_ rbzero.pov.spi_counter\[3\] _10513_ _10517_ _10519_ _10520_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__14590__A2 _08226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14366_ rbzero.debug_overlay.playerX\[-4\] _08176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_137_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16105_ _09645_ _09647_ _09648_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16867__A1 _08029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13317_ rbzero.spi_registers.texadd0\[0\] _07127_ _07130_ _07040_ _07131_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__16006__I _09550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17085_ _10447_ _10467_ _10468_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_172_Right_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_161_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14297_ rbzero.debug_overlay.vplaneY\[-7\] _08107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25319__I _06102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16036_ _09595_ _09596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13248_ gpout0.hpos\[2\] _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__24223__I _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14889__C _08595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13179_ rbzero.spi_registers.texadd3\[16\] _06922_ _06992_ rbzero.spi_registers.texadd2\[16\]
+ _06918_ rbzero.spi_registers.texadd1\[16\] _06993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_202_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80_i_clk clknet_5_30__leaf_i_clk clknet_leaf_80_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17987_ _11130_ _11131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_53_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19726_ _12497_ _12498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22678__I _11409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20179__A1 _12950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16938_ _08057_ _10348_ _10353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__21915__A2 _10474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17044__A1 _08152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19657_ _12424_ _12429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16676__I _09897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16869_ _10281_ _10293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_205_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23117__A1 _12950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_95_i_clk clknet_5_26__leaf_i_clk clknet_leaf_95_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_149_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18608_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _11623_ _11624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_189_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19588_ rbzero.debug_overlay.playerX\[-6\] _11096_ _12359_ _12158_ _12360_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_88_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14948__A4 _07225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18539_ _11584_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22340__A2 _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Left_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__18395__I1 rbzero.tex_g1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15358__A1 rbzero.mapdyw\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21550_ _12777_ _02114_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20926__I _12713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22891__A3 _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20501_ _12422_ _12586_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21481_ _02446_ _02566_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_133_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25290__A1 _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14030__B2 _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20432_ _01429_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_23220_ _03975_ _04074_ _04075_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14581__A2 _07822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23840__A2 _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16858__A1 _08049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23151_ _03618_ _04005_ _04007_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20363_ _01365_ _01452_ _01456_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_33_i_clk clknet_5_22__leaf_i_clk clknet_leaf_33_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_31_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25229__I _06012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22102_ _03090_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23082_ _03726_ _03812_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20294_ _12660_ _01388_ _12666_ _12700_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_140_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15755__I _09349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22033_ _03044_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26910_ _00820_ clknet_leaf_126_i_clk rbzero.tex_r1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_246_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_244_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_244_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_48_i_clk clknet_5_17__leaf_i_clk clknet_leaf_48_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_26841_ _00751_ clknet_leaf_190_i_clk rbzero.tex_r0\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_209_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19671__B _12442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_227_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26772_ _00682_ clknet_leaf_198_i_clk rbzero.tex_g1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_215_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23984_ _04775_ _04776_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17035__A1 _08162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25723_ _06476_ _06504_ _06506_ _06507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_138_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22935_ _03651_ _03792_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16586__I _09973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25654_ _05889_ _05973_ _06438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_104_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22866_ _02530_ _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_104_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_119_Left_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24605_ _05385_ _05388_ _05378_ _05389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_27_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21817_ _02859_ _02860_ _02863_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25585_ _06325_ _06368_ _06369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_38_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22797_ _02340_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_27324_ _01229_ clknet_leaf_117_i_clk rbzero.traced_texa\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24536_ _05276_ _05320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21748_ _10449_ _09982_ _09921_ rbzero.wall_tracer.rayAddendX\[-5\] _02802_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27255_ _01160_ clknet_leaf_90_i_clk rbzero.wall_tracer.visualWallDist\[-5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_0_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24467_ _05244_ _05245_ _05246_ _05250_ _05251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_21679_ _02743_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26206_ _00116_ clknet_leaf_9_i_clk rbzero.spi_registers.texadd0\[21\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14220_ _07983_ _07995_ _08030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_23418_ _03800_ _03930_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22095__A1 _08374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27186_ _01091_ clknet_leaf_73_i_clk rbzero.wall_tracer.size\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_24398_ _05143_ _05165_ _05170_ _05181_ _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_190_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23831__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16849__A1 _08175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20645__A2 _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14151_ rbzero.row_render.texu\[4\] _07570_ _07961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26137_ _00047_ clknet_leaf_218_i_clk rbzero.map_overlay.i_otherx\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23349_ _03845_ _02482_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_145_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_128_Left_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__21667__I _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13102_ _06915_ _06916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_120_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26068_ _06663_ _06684_ _06837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_238_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14082_ rbzero.tex_r1\[35\] _07855_ _07613_ _07892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25019_ _05758_ _05801_ _05803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_17910_ _08085_ _11017_ _11054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_237_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18890_ rbzero.traced_texa\[5\] _07279_ _11805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17841_ _10845_ _10755_ _10988_ _10989_ _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_246_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_206_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15824__A2 _09118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14984_ gpout0.vpos\[8\] _08786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17772_ _10943_ _10684_ _10939_ _10945_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_234_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19511_ _12282_ _12283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_191_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13935_ rbzero.map_overlay.i_mapdx\[2\] _06873_ _07746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_16723_ _10160_ _10163_ _09028_ _10164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_233_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_137_Left_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19442_ rbzero.wall_tracer.stepDistX\[-10\] _12214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_16654_ _08094_ _08103_ _10100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_159_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13866_ rbzero.debug_overlay.playerX\[1\] _07677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_198_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15605_ _09272_ _09273_ _09267_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_157_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16585_ _10033_ _10034_ _10035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_19373_ rbzero.tex_b1\[61\] rbzero.tex_b1\[60\] _12151_ _12152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13797_ _07468_ _07608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_241_Right_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18324_ _11434_ _08753_ _11450_ _11457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_15536_ rbzero.spi_registers.texadd0\[21\] _09218_ _09222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18255_ _11397_ _11399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_211_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15467_ _07123_ _09124_ _09171_ _09126_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_155_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18216__I _11301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17206_ _10558_ _10559_ _10560_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_182_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22086__A1 _08379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14418_ _08226_ _08227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14563__A2 _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18186_ _11299_ _11314_ _11329_ _11330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15398_ _07967_ _09065_ _09121_ _09068_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__23822__A2 _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_146_Left_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_176_i_clk_I clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17137_ rbzero.pov.ready_buffer\[8\] _10472_ _10507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14349_ rbzero.debug_overlay.facingY\[0\] _08159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_90_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17068_ _08129_ _10455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22389__A2 _08049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16019_ _09547_ _09583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_55_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_226_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25327__A2 _05998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_222_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17017__A1 _08160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22010__A1 _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19709_ _12480_ _12481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_192_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20981_ _02067_ _02069_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_204_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22720_ _11175_ _12374_ _03583_ _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_189_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22651_ _02789_ _03521_ _03523_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_24_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23510__A1 _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21602_ _02573_ _02686_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_25370_ _05890_ _06154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22582_ _12170_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24321_ _04977_ _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_21533_ _02514_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_145_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_27040_ _00950_ clknet_leaf_159_i_clk rbzero.tex_g0\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24252_ _04976_ _04986_ _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_173_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26490__D _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21464_ _02547_ _02548_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19666__B _10323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23813__A2 _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23203_ _04058_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20415_ _12626_ _12918_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21395_ _01967_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24183_ _04966_ _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23134_ _03975_ _03978_ _03990_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20346_ _01421_ _01440_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22624__I0 rbzero.wall_tracer.texu\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23065_ _03921_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20277_ _01370_ _12974_ _01371_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_101_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22016_ rbzero.wall_tracer.stepDistY\[-11\] _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__25869__A3 _06652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26824_ _00734_ clknet_leaf_178_i_clk rbzero.tex_g1\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__22001__A1 _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26755_ _00665_ clknet_leaf_222_i_clk gpout0.vpos\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_23967_ _04762_ _04763_ _04752_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_169_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14490__A1 rbzero.tex_g0\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25706_ _06436_ _06437_ _06490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13720_ _07482_ _07531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_86_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22918_ _03703_ _03744_ _03701_ _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26686_ _00596_ clknet_leaf_25_i_clk rbzero.pov.ready_buffer\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23898_ _04685_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25637_ _06420_ _06376_ _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__24466__C _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13651_ _07421_ _07462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_85_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22849_ _02620_ _02639_ _03707_ _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_14_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14242__A1 _08029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19420__I _12191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14242__B2 _08041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16370_ _08959_ _09842_ _09848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25568_ _06328_ _06276_ _06352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13582_ _07363_ _07392_ _07393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_183_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27307_ _01212_ clknet_leaf_112_i_clk rbzero.traced_texa\[-11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15321_ _09062_ _09063_ _09055_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24519_ _05283_ _05303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25499_ _05725_ _06012_ _06283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_152_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18040_ rbzero.wall_tracer.trackDistY\[2\] _11184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_152_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22068__A1 _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27238_ _01143_ clknet_leaf_82_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15252_ _09010_ _09012_ _09003_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__23804__A2 _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14203_ _08012_ _08008_ _08013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15183_ _08957_ _08952_ _08958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27169_ _01074_ clknet_leaf_51_i_clk rbzero.wall_tracer.rayAddendX\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14134_ _07507_ _07936_ _07943_ _07944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__26699__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19991_ _12752_ _12753_ _12763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_123_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13908__I gpout0.vpos\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18942_ _11841_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14065_ _07870_ _07871_ _07874_ _07838_ _07604_ _07875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__23826__B _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_219_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13520__A3 _07330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18873_ rbzero.traced_texa\[1\] rbzero.texV\[1\] _11790_ _11792_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_219_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17824_ _10972_ _10739_ _10975_ _10978_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_146_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14967_ _07175_ _08755_ net6 _08770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17755_ _10927_ _10670_ _10930_ _10933_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_206_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16706_ _10140_ _10087_ _10149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13918_ _07196_ rbzero.map_overlay.i_othery\[1\] _07729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22956__I _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14898_ rbzero.tex_b1\[48\] _08631_ _08704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17686_ _10881_ _10598_ _10885_ _10888_ _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_76_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19425_ _11381_ _12197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_187_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16637_ _10082_ _10083_ _10084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13849_ _07656_ _07657_ _07658_ _07659_ _07603_ _07660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__25493__A1 _06271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17970__A2 _11099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19356_ _12142_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14784__A2 _07629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16568_ _10019_ _10020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18307_ _08869_ _11444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15519_ rbzero.spi_registers.buf_texadd0\[16\] _09209_ _09210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16499_ _09948_ _09940_ _09955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19287_ rbzero.tex_b1\[24\] rbzero.tex_b1\[23\] _12099_ _12103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_154_Left_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23787__I _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18238_ _07233_ _11381_ _11382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__13339__A3 _07152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15733__A1 rbzero.spi_registers.buf_texadd2\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18169_ rbzero.map_overlay.i_mapdy\[2\] _11300_ rbzero.map_rom.i_row\[4\] _07754_
+ _11312_ _11313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_187_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20200_ _12432_ _12971_ _12972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21180_ _02150_ _02155_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_229_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20131_ _12628_ _12880_ _12903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_187_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24220__A2 _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_224_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_241_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20062_ rbzero.wall_tracer.visualWallDist\[-11\] _12834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_163_Left_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_225_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_206_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24870_ _05303_ _05464_ _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23821_ _03287_ _03069_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_202_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26540_ _00450_ clknet_leaf_23_i_clk rbzero.pov.spi_buffer\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23752_ _12035_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_68_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18202__A3 _11344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20964_ _01990_ _02026_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_239_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22703_ _03568_ _11220_ _03569_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_239_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26471_ _00381_ clknet_leaf_45_i_clk rbzero.debug_overlay.playerY\[-3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23683_ _03520_ _04532_ _04533_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20895_ _01965_ _01984_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__24287__A2 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25422_ _06194_ _06195_ _06197_ _06206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_22634_ _09944_ _03483_ _03473_ _03484_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_49_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14775__A2 _08494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_172_Left_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_81_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25353_ _06104_ _06105_ _06136_ _06137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__20848__A2 _12647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22565_ _09939_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18910__A1 rbzero.traced_texa\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24304_ _05079_ _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_134_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21516_ _01952_ _02349_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25284_ _06051_ _06040_ _06068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14527__A2 _07901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22496_ rbzero.wall_tracer.size\[5\] _03417_ _03418_ rbzero.row_render.size\[5\]
+ _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27023_ _00933_ clknet_leaf_132_i_clk rbzero.tex_g0\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
X_24235_ _05008_ _05018_ _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21447_ _02531_ _02532_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_133_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24166_ _04821_ _04824_ _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_21378_ _02338_ _02347_ _02463_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_247_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13728__I _07443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23117_ _12950_ _03965_ _03972_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20329_ _13001_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16104__I _09614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24097_ _04839_ _04881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_112_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24211__A2 _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_181_Left_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__21945__I _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_229_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_23048_ _03847_ _03855_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_244_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22773__A2 _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15870_ rbzero.spi_registers.buf_floor\[4\] _09463_ _09471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20784__A1 _12472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14821_ _07770_ _08627_ _07231_ _08628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_231_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_216_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26807_ _00717_ clknet_leaf_174_i_clk rbzero.tex_g1\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA_clkbuf_leaf_124_i_clk_I clknet_5_18__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24999_ _05526_ _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14463__A1 _08264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14752_ _08553_ _08555_ _08557_ _08558_ _08334_ _08559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_17540_ _10797_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__20536__A1 _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26738_ _00648_ clknet_leaf_40_i_clk rbzero.pov.ready_buffer\[68\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21680__I _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13703_ rbzero.tex_r0\[57\] _07513_ _07514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17471_ _07052_ _06876_ _06860_ _10757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_14683_ _07222_ _08490_ _08193_ _08491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_26669_ _00579_ clknet_leaf_40_i_clk rbzero.pov.ready vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19210_ _12048_ _12051_ _12052_ _12053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_157_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16422_ _09885_ _09886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13634_ _07443_ _07444_ _07445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19141_ _11977_ _11984_ _11985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_156_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16353_ _09834_ _09835_ _09833_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13412__B _07222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13565_ _07363_ _07100_ _07375_ _07376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__18901__A1 rbzero.traced_texa\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15304_ rbzero.spi_registers.buf_mapdx\[0\] _09045_ _09051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19072_ _11914_ _11915_ _11916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16284_ _09761_ _09784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14518__A2 _07890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13496_ _07282_ _07283_ _07307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_136_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16723__B _09028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18023_ rbzero.wall_tracer.trackDistY\[1\] _11167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_140_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15235_ rbzero.spi_registers.spi_buffer\[20\] _08992_ _08999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_49_i_clk_I clknet_5_17__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20245__B _12182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15166_ _08941_ _08943_ _08934_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22461__A1 _07147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13638__I _07444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14117_ _07889_ _07904_ _07926_ _07927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19974_ _12745_ _12746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15097_ _08864_ _08888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_182_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18925_ rbzero.tex_g0\[2\] rbzero.tex_g0\[1\] _11830_ _11832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14048_ rbzero.tex_r1\[9\] _07857_ _07646_ _07858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_182_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22764__A2 _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18856_ _11774_ _11777_ _11778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_158_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17807_ _10946_ _10968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_222_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18787_ rbzero.tex_r1\[58\] rbzero.tex_r1\[57\] _11724_ _11726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15999_ _09525_ _09562_ _09569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24910__B1 _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17738_ _10915_ _10923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19393__A1 _12163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17669_ _10875_ rbzero.pov.ready_buffer\[12\] _10878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19060__I _11892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19408_ _12179_ _12180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_148_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20680_ _01666_ _01771_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15954__A1 _09518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19145__A1 _08162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19339_ _12132_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25218__A1 _05996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_234_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19696__A2 _12465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22350_ _11145_ _03245_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14509__A2 _08317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21301_ _02386_ _02387_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22281_ _03200_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19448__A2 _12169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24020_ _04764_ rbzero.wall_tracer.rcp_fsm.operand\[-1\] _04757_ rbzero.wall_tracer.rcp_fsm.operand\[-3\]
+ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_142_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21232_ _02246_ _02287_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21163_ _02250_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20114_ _12471_ _12481_ _12557_ _12885_ _12886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_25971_ _06745_ _06746_ _06750_ _06695_ _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_21094_ _02180_ _02125_ _02181_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20045_ _12789_ _12817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_24922_ _05666_ _05668_ _05659_ _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_198_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24853_ _05636_ _05637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_240_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23804_ _03283_ _03067_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__20518__A1 _12283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24784_ _05513_ _05514_ _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21996_ rbzero.wall_tracer.size_full\[5\] _03005_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19384__A1 rbzero.hsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26523_ _00433_ clknet_leaf_54_i_clk rbzero.debug_overlay.vplaneY\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23735_ _04568_ _04578_ _03574_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20947_ _02030_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__21191__A1 _12713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26454_ _00364_ clknet_leaf_46_i_clk rbzero.debug_overlay.playerX\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23666_ _04515_ _04516_ _04517_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14748__A2 _08554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20878_ _12697_ _12699_ _01966_ _01967_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_113_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25405_ _06187_ _06188_ _06189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22617_ _11129_ _03489_ _09927_ _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26385_ _00295_ clknet_leaf_14_i_clk rbzero.spi_registers.buf_texadd2\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__19687__A2 _12447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23597_ _04364_ _04430_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13420__A2 _07225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25336_ _06010_ _06088_ _06083_ _06120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13350_ _07147_ _07158_ _07159_ _07150_ _07160_ _07161_ _07162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_183_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19151__A4 _11994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22548_ _11287_ _03449_ _03450_ rbzero.traced_texa\[-2\] _03452_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25267_ _06050_ _06051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15173__A2 _08940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13281_ _06957_ _06969_ _07095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18314__I _11444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16370__A1 _08959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22479_ _03408_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_50_i_clk_I clknet_5_17__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15020_ _08816_ _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_27006_ _00916_ clknet_leaf_200_i_clk rbzero.tex_g0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24218_ _04940_ _04992_ _04995_ _05001_ _05002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_25198_ _05321_ _05982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24149_ _04843_ _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_130_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21675__I _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16971_ _10374_ _10381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22746__A2 rbzero.wall_tracer.stepDistX\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18710_ _11671_ _11682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15922_ rbzero.spi_registers.buf_otherx\[4\] _09510_ _09511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19690_ _12417_ _12418_ _12462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_232_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18641_ _11642_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15853_ _09457_ _08827_ _09458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_160_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14804_ _07803_ _08602_ _08610_ _08611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_207_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18572_ _11603_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14987__A2 _08788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15784_ _09404_ _09405_ _09406_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17523_ rbzero.tex_b0\[22\] rbzero.tex_b0\[21\] _10786_ _10788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14735_ rbzero.tex_b0\[38\] _08541_ _08316_ _08542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13921__I rbzero.map_overlay.i_othery\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_7__f_i_clk_I clknet_3_1_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14666_ rbzero.tex_g1\[51\] _07583_ _08474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14739__A2 _08233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17454_ rbzero.pov.spi_buffer\[68\] _10745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_200_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16405_ _09872_ _09873_ _09867_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13617_ _07415_ _07416_ _07427_ _07428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_157_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14597_ _07480_ _08386_ _08391_ _08396_ _08404_ _08405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_17385_ rbzero.pov.spi_buffer\[51\] _10685_ _10693_ _10694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13411__A2 _07212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19124_ rbzero.debug_overlay.facingY\[-6\] _10030_ _11968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16336_ rbzero.spi_registers.buf_texadd3\[1\] _09816_ _09823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13548_ _07354_ _07357_ _07353_ _07359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19055_ _11905_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16267_ _09747_ _09771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_164_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13479_ _07288_ _07289_ _07290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18006_ rbzero.wall_tracer.trackDistY\[7\] _11150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15218_ _07166_ _08986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16198_ _09717_ _09718_ _09712_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14911__A2 _07876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13368__I gpout0.vpos\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15149_ _08906_ _08929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16113__A1 _09000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19957_ _12315_ _12318_ _12729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15583__I _08882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18099__C _11200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18908_ rbzero.traced_texa\[9\] _07259_ _11819_ _11820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_226_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19888_ _12659_ _12660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_184_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18839_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] _11763_ _11764_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_223_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21850_ _08126_ _08134_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_223_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18169__A2 _11300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20801_ _01781_ _01891_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_65_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_219_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_236_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21781_ _02830_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_236_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13831__I _07343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23520_ _04289_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_20732_ _12487_ _01535_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_186_Right_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23451_ _04210_ _04303_ _04304_ _04228_ _04208_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_175_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20663_ _01753_ _01754_ _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_135_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22365__B _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22402_ _03340_ _03346_ _03347_ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26170_ _00080_ clknet_leaf_233_i_clk rbzero.color_sky\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_98_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23382_ _04019_ _04113_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20594_ _01681_ _01685_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25121_ _05884_ _05904_ _05905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22333_ rbzero.wall_tracer.trackDistY\[6\] _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16352__A1 _08935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4_0_i_clk clknet_0_i_clk clknet_3_4_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_131_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24414__A2 _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23975__I _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13166__A1 _06927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25052_ _05833_ _05835_ _05836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14363__B1 _08045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22264_ _03225_ _03228_ _03230_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24003_ rbzero.wall_tracer.rcp_fsm.i_data\[8\] _04773_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21215_ _02174_ _02302_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22195_ _11283_ _03166_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_130_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_247_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21146_ _12191_ _12403_ _02111_ _02233_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_245_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13469__A2 rbzero.spi_registers.vshift\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22728__A2 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15493__I _08986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25954_ _06729_ _06731_ _06734_ _06707_ _05261_ _06735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__23924__B _10508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21077_ _02041_ _02045_ _02165_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_20028_ _12792_ _12793_ _12800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24905_ _05688_ _05642_ _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25885_ _06548_ _06571_ _06668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_214_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17080__A2 _10445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24836_ _05612_ _05618_ _05620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_100_Left_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24767_ _05511_ _05516_ _05551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21979_ _03007_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14520_ rbzero.tex_g0\[51\] _08317_ _08329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23718_ _04557_ _04562_ _04563_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26506_ _00416_ clknet_leaf_30_i_clk rbzero.debug_overlay.vplaneX\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24698_ _05475_ _05479_ _05480_ _05468_ _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_56_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14451_ rbzero.tex_g0\[15\] _07818_ _08260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_23649_ _04441_ _04444_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26437_ _00347_ clknet_leaf_52_i_clk rbzero.wall_tracer.rayAddendY\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_120_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_153_Right_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_166_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13402_ gpout0.vpos\[7\] _07213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17170_ rbzero.pov.spi_counter\[5\] _10532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14382_ _07225_ _07230_ _08191_ _08192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_26368_ _00278_ clknet_leaf_5_i_clk rbzero.spi_registers.buf_texadd1\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16121_ _09660_ _09661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25319_ _06102_ _06103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13333_ _07046_ _07147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16343__A1 _08922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26299_ _00209_ clknet_leaf_217_i_clk rbzero.spi_registers.buf_otherx\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__25602__A1 _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16052_ _09522_ _09601_ _09609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21219__A2 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13264_ _07077_ _07078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16894__A2 _10252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15003_ _06900_ rbzero.wall_tracer.rcp_fsm.state\[2\] _08804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_122_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13195_ _06992_ _07009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__20523__B _12906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19811_ _12575_ _12582_ _12267_ _12583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_209_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15617__B _09278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24264__S1 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22719__A2 rbzero.wall_tracer.stepDistX\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14657__B2 _07955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19742_ rbzero.wall_tracer.size\[6\] _12514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_194_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16954_ rbzero.pov.ready_buffer\[57\] _10260_ _10366_ _10266_ _10293_ _10367_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_224_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15905_ _09497_ _09498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19673_ _12444_ _12445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16885_ _08041_ _10301_ _10307_ _10308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18624_ rbzero.tex_r0\[52\] rbzero.tex_r0\[51\] _11629_ _11633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_205_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15836_ _09445_ _09446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_204_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18555_ rbzero.tex_r0\[22\] rbzero.tex_r0\[21\] _11592_ _11594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14747__I _07811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15767_ rbzero.spi_registers.buf_texadd3\[8\] _09387_ _09394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_231_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17506_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _10775_ _10778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15909__A1 _08950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14718_ rbzero.tex_b0\[40\] _08227_ _08525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18486_ _11543_ _11554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20902__A1 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15698_ rbzero.spi_registers.buf_texadd2\[14\] _09340_ _09343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17437_ rbzero.pov.spi_buffer\[64\] _10732_ _10729_ _10733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14649_ rbzero.tex_g1\[56\] _07599_ _08457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_60_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_214_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20484__I _12301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_231_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17368_ rbzero.pov.spi_buffer\[46\] _10681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_144_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19107_ _11949_ _11950_ _11951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_82_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16319_ _09808_ _09809_ _09807_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17299_ _10618_ _10630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_207_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19038_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _11893_ _11896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_93_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14896__A1 _07624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21000_ _02087_ _02088_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23907__A1 _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_242_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_242_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22951_ _03668_ _03672_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_223_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13871__A2 _07681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21902_ _02904_ _11069_ _08123_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25670_ _05983_ _06013_ _06387_ _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_3_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17062__A2 _10445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22882_ _03729_ _03740_ _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24621_ _05396_ _05404_ _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__24332__B2 _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21833_ _11020_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21146__A1 _12191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27340_ _01245_ clknet_leaf_36_i_clk rbzero.texu_hot\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24552_ _05335_ _05336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21764_ _02815_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__19669__B _10217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__25250__I _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23503_ _04346_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_20715_ _12426_ _12787_ _01803_ _01805_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_27271_ _01176_ clknet_leaf_204_i_clk rbzero.wall_tracer.wall\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24483_ _05266_ _05267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15376__A2 _09104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21695_ _12036_ _12027_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_26222_ _00132_ clknet_leaf_6_i_clk rbzero.spi_registers.texadd1\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23434_ _04286_ _04287_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_19_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22646__A1 _12775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20646_ _01679_ _01737_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_223_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17189__B _10174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26153_ _00063_ clknet_leaf_221_i_clk rbzero.map_overlay.i_mapdy\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_22_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14392__I _07928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23365_ _03734_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_78_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20577_ _01628_ _01653_ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_190_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25104_ _05336_ _05267_ _05311_ _05888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_15_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22316_ _03253_ _03272_ _03273_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14325__C gpout0.vpos\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26084_ _06846_ _03022_ _06844_ _06849_ _11825_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_15_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16876__A2 _10283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23296_ _12676_ _04150_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25035_ _05685_ _05748_ _05752_ _05819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__26014__C _05242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22247_ _11206_ _03206_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22178_ _11039_ _03117_ _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21129_ _02215_ _02216_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_246_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_26986_ _00896_ clknet_leaf_171_i_clk rbzero.tex_g0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_109_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24571__A1 _05351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25937_ _10987_ _06719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_219_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22050__S _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13951_ _07219_ _07757_ _07751_ _07760_ _07761_ _07762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XPHY_EDGE_ROW_222_Right_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16670_ _08096_ _10107_ _10115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__20569__I _09973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13882_ rbzero.debug_overlay.playerY\[4\] _07693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_25868_ _06651_ _06371_ _06652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_198_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15621_ rbzero.spi_registers.texadd1\[19\] _09279_ _09285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_122_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24819_ _05318_ _05600_ _05602_ _05603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_158_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25799_ _06557_ _06558_ _06480_ _06523_ _06583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_154_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14811__B2 _08364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18340_ _11466_ _11465_ _07176_ _11469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15552_ _09231_ _09233_ _09229_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14503_ _08245_ _08307_ _08311_ _08312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__15900__B _09491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15483_ rbzero.spi_registers.buf_texadd0\[7\] _09030_ _09183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18271_ _11403_ _11405_ _11413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15367__A2 _09097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20360__A2 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16715__C _10067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17222_ rbzero.pov.spi_buffer\[9\] _10568_ _10565_ _10573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14434_ rbzero.tex_g0\[4\] _08206_ _08243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_126_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_172_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput14 i_gpout2_sel[2] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput25 i_tex_in[1] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17153_ _10518_ rbzero.pov.spi_counter\[5\] rbzero.pov.spi_counter\[4\] _10519_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_14365_ rbzero.debug_overlay.playerX\[5\] _08175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_137_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13316_ _07127_ _07128_ _07129_ _07130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_16104_ _09614_ _09648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14327__B1 _08017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16867__A2 _10283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17084_ rbzero.pov.ready_buffer\[16\] _10445_ _10468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14296_ _08105_ _08106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_223_i_clk clknet_5_2__leaf_i_clk clknet_leaf_223_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16035_ _08851_ _09544_ _09595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13247_ _07047_ _07058_ _07060_ _07061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_58_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22024__I _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13178_ _06925_ _06992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_237_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17986_ _11129_ _08373_ _07775_ _07235_ _11130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__22959__I _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_238_i_clk clknet_5_4__leaf_i_clk clknet_leaf_238_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_224_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19725_ _12496_ _12497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_53_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16937_ rbzero.debug_overlay.playerY\[2\] _10352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__20179__A2 _12728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19656_ _12414_ _12428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_205_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_172_i_clk_I clknet_5_9__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16868_ _10272_ _10292_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_220_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24314__A1 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18607_ _11607_ _11623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15819_ _09431_ _09432_ _09430_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_220_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19587_ _12320_ _12322_ _10197_ _12325_ _12359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_177_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14802__A1 _07601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16799_ _10231_ _10232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18538_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _11581_ _11584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15810__B _09417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18469_ rbzero.tex_g1\[49\] rbzero.tex_g1\[48\] _11544_ _11545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_173_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20500_ _01591_ _01592_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_145_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21480_ _02449_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_16_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20431_ _12906_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19936__C _12223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23150_ _03892_ _04006_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20362_ _01369_ _01451_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14869__A1 _08316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22101_ _03085_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_97_i_clk_I clknet_5_26__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23081_ _03936_ _03937_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20293_ rbzero.wall_tracer.visualWallDist\[1\] _12228_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_73_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22032_ rbzero.wall_tracer.rcp_fsm.o_data\[-7\] _03043_ _03030_ _03044_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_244_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_244_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26840_ _00750_ clknet_leaf_190_i_clk rbzero.tex_r0\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_209_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19671__C _12191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15294__A1 rbzero.map_overlay.i_othery\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23983_ _04721_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26771_ _00681_ clknet_leaf_198_i_clk rbzero.tex_g1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_215_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19243__I _12072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25722_ _06505_ _06475_ _06506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22934_ _02098_ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_138_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25653_ _05980_ _06014_ _06437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22865_ _03723_ _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_104_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16794__A1 _07709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24604_ _05387_ _05388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21816_ _02859_ _02860_ _02863_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_25584_ _06330_ _06367_ _06368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_27_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__26058__A1 _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22796_ _03654_ _02075_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_195_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__17698__I _10872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24535_ _05259_ _05266_ _05319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27323_ _01228_ clknet_leaf_117_i_clk rbzero.traced_texa\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_66_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21747_ _10463_ rbzero.wall_tracer.rayAddendX\[-5\] _02800_ _02801_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_241_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24466_ _05083_ _05248_ _05249_ _05004_ _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_27254_ _01159_ clknet_leaf_90_i_clk rbzero.wall_tracer.visualWallDist\[-6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21678_ _11349_ _02742_ _02728_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23417_ _04269_ _04270_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26205_ _00115_ clknet_leaf_8_i_clk rbzero.spi_registers.texadd0\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_27185_ _01090_ clknet_leaf_73_i_clk rbzero.wall_tracer.size\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_20629_ rbzero.wall_tracer.stepDistX\[6\] _11387_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24397_ _05171_ _05178_ _05180_ _05057_ _05086_ _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_190_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15011__I _08809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14309__B1 _08023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14150_ _07802_ _07887_ _07959_ _07960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26136_ _00046_ clknet_leaf_219_i_clk rbzero.map_overlay.i_otherx\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23348_ _03851_ _01969_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24324__I _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13101_ rbzero.wall_hot\[0\] _06914_ _06915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_26067_ _06772_ _06812_ _06836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14081_ rbzero.tex_r1\[34\] _07890_ _07891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23279_ _04025_ _04112_ _04110_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25018_ _05758_ _05801_ _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_219_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20802__B1 _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17840_ _10857_ rbzero.pov.ready_buffer\[72\] _10989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19581__C _12352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23347__A2 _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17771_ _10944_ rbzero.pov.ready_buffer\[47\] _10945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14983_ _07979_ _07707_ _08785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13296__B1 _07109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21358__A1 _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26969_ _00879_ clknet_leaf_118_i_clk rbzero.texV\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_19510_ _11386_ _12279_ _12281_ _12282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_156_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16722_ rbzero.pov.ready _10162_ _10163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_13934_ _06869_ _07744_ _07745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_156_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19441_ _12193_ _12212_ _12213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_199_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16653_ _08095_ _08118_ _10099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14297__I rbzero.debug_overlay.vplaneY\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13865_ rbzero.debug_overlay.playerY\[0\] _07676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_187_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_157_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15604_ rbzero.spi_registers.buf_texadd1\[14\] _09270_ _09273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_202_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22858__A1 _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19372_ _12135_ _12151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_174_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16584_ _10009_ _10014_ _10034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13796_ _07574_ _07606_ _07607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_186_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13063__A3 _06879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14260__A2 _08052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18323_ _10271_ _11456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_186_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15535_ _09219_ _09221_ _09217_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_139_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20333__A2 _12325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18254_ _11134_ _11397_ _11398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_15466_ rbzero.spi_registers.buf_texadd0\[2\] _09137_ _09171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_127_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_211_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17205_ rbzero.pov.spi_buffer\[5\] _10556_ _10552_ _10560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14417_ _07511_ _08226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22086__A2 _08374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18185_ _11298_ _11323_ _11328_ _11329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_170_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15397_ rbzero.spi_registers.buf_sky\[1\] _09080_ _09121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_119_i_clk_I clknet_5_18__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17136_ _10131_ _10485_ _10506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_162_i_clk clknet_5_10__leaf_i_clk clknet_leaf_162_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14348_ _08155_ _08040_ _08045_ _08156_ _08157_ _08035_ _08158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_12_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14279_ _07216_ _07200_ _07719_ _08089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_90_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17067_ _10453_ _10454_ _10436_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_228_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16018_ _09581_ _09582_ _09576_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_55_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_177_i_clk clknet_5_8__leaf_i_clk clknet_leaf_177_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_237_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17969_ _11112_ _11100_ _11113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13826__A2 _07635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19708_ _12479_ _12480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_100_i_clk clknet_5_26__leaf_i_clk clknet_leaf_100_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_20980_ _02068_ _12919_ _01704_ _02066_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_178_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19639_ _12410_ _12411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_204_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22650_ rbzero.wall_tracer.trackDistX\[-11\] _03522_ _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19714__A1 _12314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_115_i_clk clknet_5_19__leaf_i_clk clknet_leaf_115_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21601_ _02574_ _02685_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_177_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22581_ _07440_ _10072_ _03470_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_168_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24320_ _05040_ _04959_ _05037_ _05104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21532_ _02588_ _02616_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_7_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14003__A2 _07810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24251_ _04944_ _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21463_ _02547_ _02548_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_161_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15751__A2 _09375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23202_ _02115_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20414_ _01503_ _01507_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24182_ _04952_ _04957_ _04965_ _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_161_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21394_ _02361_ _02362_ _02479_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_160_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23133_ _03981_ _03989_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20345_ _01423_ _01425_ _01439_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_113_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23064_ _12676_ _02485_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_20276_ _12949_ _12963_ _12975_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_22015_ _03030_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__20260__A1 _12979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16464__B1 _09921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26823_ _00733_ clknet_leaf_177_i_clk rbzero.tex_g1\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_227_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26754_ _00664_ clknet_leaf_222_i_clk gpout0.vpos\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_230_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23966_ rbzero.wall_tracer.rcp_fsm.i_data\[-1\] _04755_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15019__A1 _08807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14490__A2 _08298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25705_ _06436_ _06437_ _06489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_86_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22917_ _03771_ _03774_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_168_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23897_ _04710_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26685_ _00595_ clknet_leaf_25_i_clk rbzero.pov.ready_buffer\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15006__I _08805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25636_ _06377_ _06419_ _06420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22848_ _02623_ _02638_ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13650_ _07460_ _07461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_151_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14242__A2 _08036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13581_ _07372_ _07385_ _07392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25567_ _06328_ _06276_ _06351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20315__A2 _12258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22779_ _03634_ _03637_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__17221__I _10571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15320_ rbzero.spi_registers.buf_mapdx\[4\] _09060_ _09063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27306_ _01211_ clknet_leaf_201_i_clk rbzero.row_render.texu\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24518_ _05298_ _05301_ _05302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25498_ _06030_ _06050_ _06005_ _06012_ _06282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_109_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_152_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27237_ _01142_ clknet_leaf_81_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15251_ _09011_ _09001_ _09012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24449_ _05232_ _05233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15742__A2 _09375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_120_i_clk_I clknet_5_18__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14202_ _07373_ _07981_ _08012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_117_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15182_ rbzero.spi_registers.spi_buffer\[8\] _08957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_27168_ _01073_ clknet_leaf_51_i_clk rbzero.wall_tracer.rayAddendX\[-3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15676__I _09302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14133_ _07937_ _07939_ _07942_ _07923_ _07924_ _07943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_10_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26119_ _00029_ clknet_leaf_4_i_clk rbzero.spi_registers.spi_buffer\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19990_ _12752_ _12753_ _12762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_94_i_clk clknet_5_19__leaf_i_clk clknet_leaf_94_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_27099_ _01009_ clknet_leaf_140_i_clk rbzero.tex_b1\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_123_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold41_I i_gpout1_sel[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18941_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _11840_ _11841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14064_ rbzero.tex_r1\[6\] _07872_ _07873_ _07874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_130_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18872_ rbzero.traced_texa\[2\] rbzero.texV\[2\] _11791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__15258__A1 _08811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17823_ _10973_ rbzero.pov.ready_buffer\[66\] _10978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_50_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13808__A2 _07577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_12__f_i_clk clknet_3_3_0_i_clk clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17754_ _10928_ rbzero.pov.ready_buffer\[42\] _10933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_221_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14966_ net27 _08755_ _08756_ net19 _08768_ _08769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_89_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_180_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14481__A2 _08288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16705_ _10127_ _10145_ _10136_ _10147_ _10148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_226_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13917_ _07684_ rbzero.map_overlay.i_othery\[4\] _07721_ _07686_ _07727_ _07728_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA_clkbuf_leaf_45_i_clk_I clknet_5_16__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17685_ _10882_ rbzero.pov.ready_buffer\[18\] _10888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_187_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14897_ _07609_ _08690_ _08702_ _08703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__19611__I _12382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_32_i_clk clknet_5_22__leaf_i_clk clknet_leaf_32_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_19424_ rbzero.debug_overlay.playerY\[-1\] _12006_ _12195_ _12196_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__22458__B _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16636_ _10065_ _08117_ _10083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13848_ rbzero.tex_r0\[20\] _07599_ _07448_ _07659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__24229__I _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25493__A2 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19355_ rbzero.tex_b1\[53\] rbzero.tex_b1\[52\] _12141_ _12142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_146_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16567_ _09938_ _10019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13779_ _07578_ _07581_ _07585_ _07588_ _07589_ _07590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_85_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18306_ _11440_ _11442_ _11443_ _11441_ _10992_ _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_72_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15518_ _09208_ _09209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19286_ _12102_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16498_ _09943_ _09947_ _09952_ _09953_ _09954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_47_i_clk clknet_5_17__leaf_i_clk clknet_leaf_47_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__25488__C _05605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18237_ _11380_ _11381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15449_ rbzero.spi_registers.buf_vshift\[3\] _09154_ _09159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18168_ rbzero.map_overlay.i_mapdy\[0\] _11301_ _11312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_187_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_187_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17119_ _09942_ _10487_ _10495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18099_ _11139_ rbzero.wall_tracer.trackDistX\[10\] _11146_ _11200_ _11243_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_229_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20130_ _12638_ _12648_ _12901_ _12902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_40_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_241_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20061_ _12193_ _12224_ _12807_ _12699_ _12833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_225_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_206_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24508__A1 _05252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13834__I _07341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17306__I _10611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23820_ _03292_ _03072_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_240_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__19935__A1 _12705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23751_ _11179_ _03056_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__23731__A2 _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20963_ _01914_ _01989_ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_205_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_68_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14209__C1 _08017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22702_ _02766_ _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_239_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_239_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23682_ _04527_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26470_ _00380_ clknet_leaf_45_i_clk rbzero.debug_overlay.playerY\[-4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__24139__I _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20894_ _01974_ _01983_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_198_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14224__A2 _08033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24287__A3 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25421_ _06194_ _06195_ _06197_ _06205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_138_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22633_ _03508_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_177_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23495__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25352_ _06130_ _06132_ _06135_ _06136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_36_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13983__A1 _07244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22564_ _09973_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24303_ _05086_ _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21515_ _12789_ _02213_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25283_ _06030_ _06047_ _06067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22495_ _03419_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__24444__C2 _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24234_ _05011_ _05015_ _05017_ _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_27022_ _00932_ clknet_leaf_149_i_clk rbzero.tex_g0\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23798__A2 rbzero.wall_tracer.stepDistY\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24995__A1 _05304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21446_ _01483_ _01608_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15496__I _09150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24165_ _04868_ _04889_ _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21377_ _02348_ _02354_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23116_ _12949_ _03965_ _03972_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_20328_ _13015_ _13026_ _01422_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_24096_ _04827_ _04840_ _04851_ _04879_ _04880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_112_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23047_ _03841_ _03876_ _03903_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20259_ _12982_ _13030_ _13031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_235_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21981__A1 rbzero.wall_tracer.size\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20784__A2 _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13744__I _07468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17216__I _10555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26806_ _00716_ clknet_leaf_174_i_clk rbzero.tex_g1\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14820_ _07243_ _08621_ _08626_ _08627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_192_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24998_ _05777_ _05781_ _05782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_162_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14751_ _07917_ _08558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_26737_ _00647_ clknet_leaf_40_i_clk rbzero.pov.ready_buffer\[67\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_203_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23949_ rbzero.wall_tracer.rcp_fsm.operand\[-4\] _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_13702_ _07508_ _07513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17470_ _10755_ _10547_ _10756_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26668_ _00578_ clknet_leaf_155_i_clk rbzero.tex_b0\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14682_ _08379_ net2 _07243_ _08489_ _08490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_16421_ rbzero.spi_registers.sclk_buffer\[1\] _08866_ _08904_ _09885_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_25619_ _06400_ _06401_ _06402_ _06403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_13633_ _07305_ _07322_ _07330_ _07444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_183_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26599_ _00509_ clknet_leaf_42_i_clk rbzero.pov.spi_buffer\[68\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19140_ _11943_ _11956_ _11984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13974__A1 _07720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16352_ _08935_ _09831_ _09835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22792__I _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13564_ _07364_ _06885_ _07371_ _07374_ _07375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_54_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15303_ _07737_ _09043_ _09050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19071_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] _11915_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16283_ rbzero.spi_registers.spi_buffer\[12\] _09782_ _09783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13495_ _07290_ _07305_ _07306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16912__A1 _07698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18022_ _11163_ _11164_ _11165_ rbzero.wall_tracer.trackDistY\[2\] _11166_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_23_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15234_ _08996_ _08998_ _08988_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18114__B1 _11256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15165_ _08942_ _08929_ _08943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22461__A2 _07150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24738__A1 _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14116_ _07555_ _07914_ _07925_ _07926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19973_ _12703_ _12743_ _12744_ _12745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15096_ _08880_ _08886_ _08887_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_201_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14151__A1 rbzero.row_render.texu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18924_ _11831_ _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22213__A2 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14047_ _07518_ _07857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_182_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19090__A1 _08155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18855_ _11775_ _11776_ _11777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_147_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13654__I _07464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17806_ _10965_ _10720_ _10961_ _10967_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_234_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18786_ _11725_ _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_207_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15998_ rbzero.spi_registers.buf_mapdy\[0\] _09560_ _09568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_222_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24910__A1 _05640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_167_Right_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17737_ _10920_ _10648_ _10916_ _10922_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__24910__B2 _05298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14949_ _08750_ _08751_ _08752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_17668_ _10850_ _10877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19407_ _07774_ _07233_ _07238_ _12179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16619_ _10066_ _10067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14485__I _07819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17599_ rbzero.tex_b0\[55\] rbzero.tex_b0\[54\] _10828_ _10831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19338_ rbzero.tex_b1\[46\] rbzero.tex_b1\[45\] _12130_ _12132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24277__I0 _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19269_ _12092_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_155_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21300_ _12704_ _02111_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22280_ _03220_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22207__I _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21231_ _02248_ _02286_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24729__A1 _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21162_ _01608_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20113_ _12884_ _12885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25970_ _06700_ _06709_ _06748_ _06749_ _06750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_21093_ _02060_ _02105_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14693__A2 _07930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13350__C1 _07160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20044_ _12788_ _12816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_24921_ _05694_ _05700_ _05701_ _05702_ _05704_ _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_217_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_24852_ _05599_ _05631_ _05636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14445__A2 _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23803_ _03283_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_3_0_0_i_clk clknet_0_i_clk clknet_3_0_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21995_ rbzero.wall_tracer.rcp_fsm.o_data\[5\] _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_24783_ _05472_ _05307_ _05567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_68_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26522_ _00432_ clknet_leaf_56_i_clk rbzero.debug_overlay.vplaneY\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_240_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23734_ _11226_ _03050_ _04577_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20946_ _02035_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14609__B _07580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_26453_ _00363_ clknet_leaf_46_i_clk rbzero.debug_overlay.playerX\[-6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_20877_ _01845_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_193_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23665_ _11141_ _04351_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25404_ _06047_ _06188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13956__A1 _07149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22616_ _03471_ _03105_ _03498_ _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_23596_ _04448_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26384_ _00294_ clknet_leaf_14_i_clk rbzero.spi_registers.buf_texadd2\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_22_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13420__A3 _07230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25335_ _05996_ _06118_ _06119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22547_ _03451_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18895__A1 rbzero.traced_texa\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13280_ _06950_ _06971_ _07094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25266_ _05725_ _06050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_22478_ _03342_ _02034_ _10040_ _07433_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_114_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27005_ _00915_ clknet_leaf_200_i_clk rbzero.tex_g0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_106_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24217_ _04996_ _05000_ _04893_ _05001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_21429_ _02506_ _02514_ _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14381__A1 _07976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25197_ _05980_ _05981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16115__I _09595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24148_ _04931_ _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_209_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24196__A2 _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24079_ _04742_ rbzero.wall_tracer.rcp_fsm.operand\[-7\] _04863_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_16970_ _10376_ _10380_ _10214_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_235_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_31_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15921_ _09494_ _09510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_200_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13892__B1 _07700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_218_i_clk_I clknet_5_3__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18640_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _11639_ _11642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15852_ _08826_ _09457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_231_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14803_ _07839_ _08606_ _08609_ _08610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_18571_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _11602_ _11603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15783_ _09383_ _09406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16785__I _07166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_125_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17522_ _10787_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14734_ _07566_ _08541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_231_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17453_ _10742_ _10735_ _10744_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_184_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23459__A1 _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14665_ rbzero.tex_g1\[49\] _07916_ _07636_ _08473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16404_ rbzero.spi_registers.spi_buffer\[19\] _09865_ _09873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13947__A1 _07244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13616_ _07417_ _07422_ _07425_ _07426_ _07427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_55_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17384_ _10658_ _10693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21640__B _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14596_ _07507_ _08403_ _08404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19123_ _11961_ _11965_ _11966_ _11967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__16734__B _10174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16335_ _09817_ _09821_ _09822_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_216_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13547_ _07353_ _07354_ _07357_ _07358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_125_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18505__I _11564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19054_ rbzero.tex_g0\[58\] rbzero.tex_g0\[57\] _11903_ _11905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16266_ rbzero.spi_registers.buf_texadd2\[8\] _09769_ _09770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13478_ rbzero.texV\[5\] _07280_ _07289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_18005_ _11147_ rbzero.wall_tracer.trackDistY\[8\] _11148_ rbzero.wall_tracer.trackDistY\[7\]
+ _11149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__13649__I _07459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15217_ _08983_ _08984_ _08985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16197_ _08983_ _09709_ _09718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24242__I _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15148_ rbzero.spi_registers.spi_buffer\[3\] _08928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_236_Right_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19956_ _12700_ _12728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15079_ _07719_ _08870_ _08871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18907_ _11817_ _11818_ _11819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_184_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19887_ _12658_ _12659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__25136__A1 _05408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18838_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] _11762_ _11763_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13317__C _07040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14427__A2 _08210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18769_ rbzero.tex_r1\[50\] rbzero.tex_r1\[49\] _11714_ _11716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13635__B1 _07328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20800_ _01784_ _01890_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21780_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] _02824_
+ _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_236_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_236_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20731_ _01816_ _01821_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22646__B _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23450_ _04212_ _04227_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20662_ _12237_ _01744_ _01752_ _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__17129__A1 rbzero.pov.ready_buffer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22401_ _03322_ _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23381_ _04023_ _04235_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18877__A1 rbzero.traced_texa\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23870__A1 _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22673__A2 _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20593_ _01683_ _01684_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_61_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25120_ _05903_ _05904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22332_ _03274_ _03285_ _03286_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25051_ _05784_ _05789_ _05834_ _05835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_116_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22263_ rbzero.wall_tracer.visualWallDist\[-7\] _03218_ _03229_ _03230_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__23622__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24002_ rbzero.wall_tracer.rcp_fsm.operand\[8\] _04722_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21214_ _02175_ _02178_ _02301_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_22194_ _03154_ _03172_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_76_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_203_Right_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__20987__A2 _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_247_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21145_ _02232_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15863__A1 _09462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14666__A2 _07583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25953_ _06627_ _06621_ _06732_ _06733_ _06632_ _06703_ _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_21076_ _02051_ _02054_ _02164_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_20027_ _12796_ _12798_ _12799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24904_ _05687_ _05639_ _05688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25884_ _06666_ _06667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_225_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24835_ _05612_ _05618_ _05619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24766_ _05502_ _05518_ _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21978_ rbzero.wall_tracer.rcp_fsm.o_data\[-2\] _12514_ _03002_ _03007_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__22361__A1 rbzero.mapdxw\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26505_ _00415_ clknet_leaf_30_i_clk rbzero.debug_overlay.vplaneX\[-6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23717_ rbzero.wall_tracer.trackDistY\[-7\] _03043_ _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20929_ _12683_ _01378_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24697_ _05468_ _05475_ _05479_ _05480_ _05481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_139_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26436_ _00346_ clknet_leaf_52_i_clk rbzero.wall_tracer.rayAddendY\[-3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14450_ rbzero.tex_g0\[12\] _08258_ _08220_ _08259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23648_ _04470_ _04498_ _04499_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_83_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13401_ _07207_ _07211_ _06859_ _07212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_14_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26367_ _00277_ clknet_leaf_5_i_clk rbzero.spi_registers.buf_texadd1\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14381_ _07976_ _07978_ _08190_ _07222_ _08191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_92_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22664__A2 _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23579_ _04337_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16120_ _09659_ _09660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_92_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25318_ _06033_ _06102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13332_ _07061_ _07082_ _07103_ _07145_ _06879_ _07146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_106_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26298_ _00208_ clknet_leaf_229_i_clk rbzero.spi_registers.buf_leak\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16051_ rbzero.spi_registers.buf_texadd0\[3\] _09597_ _09608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25249_ _06032_ _06033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_40_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13263_ _06885_ _07077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20427__A1 _12282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15002_ _08803_ net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13194_ _07003_ _07008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19810_ _12576_ _12578_ _12581_ _12166_ _12582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_102_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19741_ _12289_ _11986_ _12290_ _12512_ _12513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_159_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16953_ _07685_ _10359_ _10353_ _10366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_127_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19596__A2 _12202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15904_ _08821_ _08858_ _09497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_19672_ _12399_ _12444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_205_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16884_ _10293_ _10302_ _10306_ _10307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_95_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18623_ _11632_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15835_ _08826_ _09443_ _09444_ _09445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_91_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18554_ _11593_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15766_ rbzero.spi_registers.texadd3\[8\] _09385_ _09393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_204_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22352__A1 _11278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17505_ _10777_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_177_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14717_ _07609_ _08516_ _08523_ _08524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_87_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18485_ _11553_ _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15909__A2 _09498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15697_ rbzero.spi_registers.texadd2\[14\] _09338_ _09342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17436_ _10696_ _10732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14648_ rbzero.tex_g1\[58\] _07932_ _07946_ _08456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__24237__I _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22104__A1 _12185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_214_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_231_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17367_ _10679_ _10677_ _10680_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_231_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14579_ rbzero.tex_g1\[16\] _07816_ _08387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19106_ _08148_ _10150_ _11950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19520__A2 _11989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16318_ _09008_ _09804_ _09809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17298_ rbzero.pov.spi_buffer\[28\] _10629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19037_ _11895_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22407__A2 _08062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16249_ _09742_ _09757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14712__B _08289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16098__A1 _08983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14648__A2 _07932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19939_ _12708_ _12709_ _12711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__20005__I _12691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22950_ _03688_ _03696_ _03807_ _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_71_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22591__A1 _07028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23316__I _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21901_ _02905_ _02918_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__22220__I _09989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22881_ _03732_ _03739_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14938__I net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24620_ _05400_ _05403_ _05404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_195_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21832_ _01029_ _02874_ _02878_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_93_i_clk_I clknet_5_24__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21146__A2 _12403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18854__B _11772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14159__B _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24551_ _05269_ _05334_ _05335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_21763_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] _02805_
+ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16022__A1 _09518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23502_ _11145_ _04351_ _04354_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20714_ _01804_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27270_ _01175_ clknet_leaf_116_i_clk rbzero.wall_tracer.visualWallDist\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24482_ _05265_ _05266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21694_ _12017_ _12026_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16573__A2 _08107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26221_ _00131_ clknet_leaf_6_i_clk rbzero.spi_registers.texadd1\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20645_ _01686_ _01736_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_23433_ _03868_ _04054_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22646__A2 _12864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23364_ _03852_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26152_ _00062_ clknet_leaf_217_i_clk rbzero.map_overlay.i_mapdy\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20576_ _01570_ _01655_ _01667_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25103_ _05845_ _05852_ _05886_ _05887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22315_ _11291_ _03264_ _03257_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26083_ _06847_ _06848_ _06842_ _06849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_23295_ _04039_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_131_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14887__A2 _07561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22246_ _03202_ _03214_ _03215_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_25034_ _05809_ _05810_ net73 _05818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_104_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_22177_ rbzero.wall_tracer.rcp_fsm.i_data\[2\] _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_79_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21128_ _12696_ _02097_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26985_ _00895_ clknet_leaf_171_i_clk rbzero.tex_g0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_100_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_109_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19704__I _12475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19578__A2 _12271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25936_ _06695_ _06706_ _06717_ _05006_ _06718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_21059_ _02018_ _02019_ _02147_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13950_ gpout0.vpos\[4\] rbzero.map_overlay.i_mapdy\[1\] _07761_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_17_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22130__I _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25867_ _06318_ _06319_ _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13881_ _07690_ _07691_ _07692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_202_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15620_ _09283_ _09284_ _09278_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_198_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24818_ _05309_ _05601_ _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_122_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25798_ _06562_ _06564_ _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__18389__I0 rbzero.tex_g1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15551_ rbzero.spi_registers.buf_texadd1\[1\] _09232_ _09233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24749_ _05531_ _05532_ _05477_ _05478_ _05533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_159_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__26076__A2 _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14502_ _08308_ _08309_ _08310_ _08311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_18270_ rbzero.wall_tracer.mapX\[8\] _11404_ _11412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_204_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15482_ _06962_ _09180_ _09181_ _09182_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_83_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17221_ _10571_ _10572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_42_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14433_ rbzero.tex_g0\[7\] _08241_ _07867_ _08242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26419_ _00329_ clknet_leaf_18_i_clk rbzero.spi_registers.buf_texadd3\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13701__B _07488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27399_ _01304_ clknet_leaf_76_i_clk rbzero.wall_tracer.stepDistX\[-3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17152_ rbzero.pov.spi_counter\[6\] _10518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput15 i_gpout2_sel[3] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14364_ rbzero.debug_overlay.playerX\[-5\] _08064_ _08174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput26 i_tex_in[2] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_137_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16103_ _08990_ _09646_ _09647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13315_ rbzero.spi_registers.texadd3\[0\] _07111_ _07129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17083_ _10466_ _10443_ _10467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_220_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14295_ rbzero.debug_overlay.vplaneY\[-6\] _08105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_122_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16034_ _09593_ _09594_ _09587_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13246_ _07059_ _07060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_126_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17816__A2 rbzero.pov.ready_buffer\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13177_ _06913_ _06991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_236_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17985_ _07237_ _11129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_229_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19614__I _12282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19724_ _12495_ _12496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16936_ _10345_ _10347_ _10351_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_53_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20179__A3 _12936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_115_i_clk_I clknet_5_19__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19655_ _12426_ _12427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14758__I _07603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16867_ _08029_ _10283_ _10291_ _10292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16252__A1 _08926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15818_ rbzero.spi_registers.buf_texadd3\[21\] _09118_ _09432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18606_ _11622_ _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19586_ _12357_ _12358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_172_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21128__A2 _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16798_ rbzero.debug_overlay.playerX\[-1\] _10230_ _10231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_189_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_220_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18537_ _11583_ _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15749_ _09379_ _09380_ _09372_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19741__A2 _11986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24078__A1 _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18468_ _11543_ _11544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14566__A1 _08374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_17419_ _10717_ _10713_ _10719_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18399_ rbzero.tex_g1\[19\] rbzero.tex_g1\[18\] _11502_ _11505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20430_ _12280_ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21300__A2 _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20361_ _01449_ _01367_ _01447_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_141_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22100_ _03087_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23080_ _03800_ _03803_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20292_ _01385_ _12973_ _01386_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_141_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25954__C _05261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14442__B _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13837__I _07526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22031_ rbzero.wall_tracer.stepDistY\[-7\] _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__21064__A1 _12713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23755__B _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_244_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_244_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_209_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16491__A1 _09945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26770_ _00680_ clknet_leaf_123_i_clk rbzero.tex_g1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23982_ rbzero.wall_tracer.rcp_fsm.operand\[3\] _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_138_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input26_I i_tex_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25721_ _06384_ _06391_ _06460_ _06505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_22933_ _03655_ _03657_ _03783_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_39_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25652_ _05983_ _06006_ _06436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_196_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22864_ _02662_ _02673_ _03722_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_196_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24603_ _05363_ _05386_ _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21815_ _02846_ _02861_ _02862_ _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25583_ _06331_ _06366_ _06367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22795_ _02343_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__26058__A2 rbzero.wall_tracer.rcp_fsm.o_data\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27322_ _01227_ clknet_leaf_117_i_clk rbzero.traced_texa\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24534_ _05312_ _05316_ _05317_ _05318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_148_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21746_ _02711_ _02798_ _02799_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_27253_ _01158_ clknet_leaf_90_i_clk rbzero.wall_tracer.visualWallDist\[-7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24465_ _05197_ _05180_ _05249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21677_ _02736_ _02738_ _02741_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26204_ _00114_ clknet_leaf_8_i_clk rbzero.spi_registers.texadd0\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23416_ _04031_ _04165_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20628_ rbzero.wall_tracer.stepDistY\[6\] _01525_ _01526_ _01719_ _01720_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_27184_ _01089_ clknet_leaf_74_i_clk rbzero.wall_tracer.size_full\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24396_ _05153_ _05179_ _05088_ _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14309__B2 _08118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26135_ _00045_ clknet_leaf_218_i_clk rbzero.map_overlay.i_otherx\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23347_ _03846_ _03652_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20559_ _01643_ _01646_ _01651_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_105_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13100_ rbzero.wall_hot\[1\] _06914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_26066_ _06835_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14080_ _07632_ _07890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_23278_ _04015_ _04130_ _04132_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_219_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25017_ _05760_ _05800_ _05801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_22229_ _03199_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__20802__A1 rbzero.traced_texVinit\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20802__B2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17770_ _10936_ _10944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26968_ _00878_ clknet_leaf_117_i_clk rbzero.texV\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14982_ _08775_ _08777_ _08783_ _08784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13296__A1 rbzero.spi_registers.texadd2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21358__A2 _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16721_ _08875_ _10161_ _10162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_25919_ _06683_ _06687_ _06698_ _06700_ _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_13933_ _07740_ _07742_ _07743_ _07744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_233_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26899_ _00809_ clknet_leaf_132_i_clk rbzero.tex_r1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_19440_ _12211_ _12212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16652_ _10079_ _10080_ _10084_ _10098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22795__I _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13864_ _07199_ rbzero.debug_overlay.playerY\[2\] _07675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_232_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15603_ rbzero.spi_registers.texadd1\[14\] _09268_ _09272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_186_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19371_ _12150_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_202_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16583_ _10032_ _10031_ _10033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22858__A2 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13795_ _07590_ _07605_ _07606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_186_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18322_ _11454_ _11455_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15534_ rbzero.spi_registers.buf_texadd0\[20\] _09220_ _09221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21204__I _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18253_ _09925_ _11379_ _11396_ _11397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_139_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15465_ _09169_ _09170_ _09162_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_211_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17204_ _10544_ _10559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14416_ rbzero.tex_g0\[21\] _08202_ _08225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_231_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18184_ _11324_ _11325_ _11326_ _11327_ _11328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24480__A1 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22086__A3 _07775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15396_ _09114_ _09116_ _09120_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_108_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17135_ _10024_ _10397_ _10505_ _09441_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_14347_ rbzero.debug_overlay.facingY\[-8\] _08157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_41_i_clk_I clknet_5_16__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17066_ rbzero.pov.ready_buffer\[12\] _10434_ _10454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_204_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14278_ rbzero.debug_overlay.facingX\[-4\] _08088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13657__I _07328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16017_ _08962_ _09574_ _09582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13229_ _07034_ _07042_ _07043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_55_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21597__A2 _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_226_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15872__I _09429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17968_ rbzero.map_rom.f3 _11112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22546__A1 _11288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22546__B2 rbzero.traced_texa\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19707_ _12439_ _12440_ _12442_ _12479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_240_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16919_ _10336_ _10337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_192_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17899_ rbzero.debug_overlay.facingX\[-3\] _11025_ _11043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_79_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19638_ _12409_ _12410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_204_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14787__A1 _08304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19569_ _12320_ _12322_ _10190_ _12325_ _12341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_193_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_21600_ _02575_ _02684_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_34_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22580_ rbzero.wall_tracer.wall\[1\] _09974_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21531_ _02606_ _02615_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_168_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24250_ _04733_ _04903_ _05034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_21462_ _12522_ _01378_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23274__A2 _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20413_ _01504_ _01505_ _01506_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_23201_ _04051_ _04056_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21393_ _02214_ _02363_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24181_ _04958_ _04961_ _04962_ _04964_ _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__14951__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18150__A1 _11290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20344_ _01426_ _01427_ _01438_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_23132_ _03983_ _03988_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__23026__A2 _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24361__S _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23063_ _03794_ _03795_ _03916_ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__13514__A2 _07324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20275_ _12966_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22014_ _03029_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__25256__I _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16464__A1 _09915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26822_ _00732_ clknet_leaf_178_i_clk rbzero.tex_g1\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13278__A1 _06906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14398__I _08206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26753_ _00663_ clknet_leaf_219_i_clk rbzero.hsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_98_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23965_ _04761_ _04758_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19253__I1 rbzero.tex_b1\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15019__A2 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25704_ _06435_ _06441_ _06488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_242_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22916_ _03772_ _03709_ _03720_ _03773_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_169_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26684_ _00594_ clknet_leaf_26_i_clk rbzero.pov.ready_buffer\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23896_ rbzero.wall_tracer.rcp_fsm.o_data\[4\] _03764_ _04693_ _04710_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17964__A1 _11106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16827__B _10256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25635_ _06383_ _06418_ _06419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_190_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22847_ _02656_ _03704_ _03705_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_222_i_clk clknet_5_2__leaf_i_clk clknet_leaf_222_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_168_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25566_ _06336_ _06345_ _06349_ _06350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_13580_ _07389_ _07390_ _07391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22778_ _03635_ _03636_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27305_ _01210_ clknet_leaf_189_i_clk rbzero.row_render.texu\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24517_ _05300_ _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_164_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21729_ _02744_ _02785_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25497_ _06034_ _06087_ _06281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17192__A2 _10547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27236_ _01141_ clknet_leaf_84_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15250_ rbzero.spi_registers.spi_buffer\[22\] _09011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__20863__I _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24448_ _05231_ _05232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_237_i_clk clknet_5_6__leaf_i_clk clknet_leaf_237_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__24462__A1 _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23265__A2 _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14201_ _08010_ _08011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_117_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13753__A2 _07563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15181_ _08955_ _08940_ _08956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27167_ _01072_ clknet_leaf_51_i_clk rbzero.wall_tracer.rayAddendX\[-4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24379_ _05017_ _05163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_134_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18141__A1 _11281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14132_ rbzero.tex_r1\[52\] _07940_ _07941_ _07942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26118_ _00028_ clknet_leaf_4_i_clk rbzero.spi_registers.spi_buffer\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__24214__A1 _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27098_ _01008_ clknet_leaf_140_i_clk rbzero.tex_b1\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_160_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14082__B _07613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21028__A1 _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26049_ _06785_ _06819_ _06820_ _06756_ _06821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_18940_ _11829_ _11840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14063_ rbzero.tex_r1\[7\] _07835_ _07873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_37_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_148_Right_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_167_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18871_ _11786_ _11789_ _11790_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_218_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15692__I _09302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19164__I _12007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17822_ _10972_ _10737_ _10975_ _10977_ _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__22528__A1 _12595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14965_ net6 _08767_ _08768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17753_ _10927_ _10668_ _10930_ _10932_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_89_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_221_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16704_ _10127_ _10146_ _10136_ _10147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13916_ rbzero.map_overlay.i_otherx\[3\] _06864_ _07727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17684_ _10881_ _10596_ _10885_ _10887_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_18_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14896_ _07624_ _08695_ _08701_ _08702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__16758__A2 _08180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Left_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16635_ _08104_ _09928_ _10082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19423_ _10337_ _10338_ _12015_ _12195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_18_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13847_ rbzero.tex_r0\[21\] _07576_ _07658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13940__I rbzero.map_overlay.i_mapdy\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16566_ _10004_ _10006_ _10014_ _10017_ _10018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_146_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19354_ _12135_ _12141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13778_ _07449_ _07589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__22700__A1 _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15517_ _08883_ _09208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18305_ _07102_ _07423_ _07992_ _11443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_19285_ rbzero.tex_b1\[23\] rbzero.tex_b1\[22\] _12099_ _12102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16497_ _09926_ _09953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18236_ _08379_ rbzero.trace_state\[2\] rbzero.trace_state\[1\] _11380_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_15448_ rbzero.spi_registers.vshift\[3\] _09151_ _09158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14941__A1 rbzero.vga_sync.vsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18167_ _07757_ _11306_ _11307_ rbzero.map_overlay.i_mapdy\[4\] _11310_ _11311_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_170_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15379_ _09105_ _09106_ _09100_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_187_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_187_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_68_Left_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17118_ _10493_ _10494_ _10492_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18098_ _11217_ _11215_ _11227_ _11241_ _11242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_128_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16694__A1 _09953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17049_ _10439_ _10440_ _10436_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22767__A1 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20060_ _12809_ _12811_ _12832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_241_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15816__B _09430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14720__B _08308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15249__A2 _08917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16446__A1 rbzero.debug_overlay.vplaneY\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20242__A2 _12917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_206_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Left_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_240_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19935__A2 _12706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23750_ _04590_ _04591_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14011__I _07341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14209__B1 _08011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20962_ _02047_ _02050_ _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_68_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14209__C2 _08018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22701_ _03556_ _03566_ _03567_ _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_27__f_i_clk_I clknet_3_6_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_239_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23681_ _04530_ _04531_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20893_ _12836_ _01982_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_178_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25420_ _06181_ _06188_ _06204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22632_ rbzero.wall_tracer.w\[0\] _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__17549__I1 rbzero.tex_b0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25351_ _06133_ _06134_ _06135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_181_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22563_ _03460_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__19677__C _12448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24302_ _05085_ _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_21514_ _02592_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25282_ _06065_ _05999_ _06066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24444__A1 _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22494_ rbzero.wall_tracer.size\[4\] _03417_ _03418_ _07363_ _03419_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27021_ _00931_ clknet_leaf_150_i_clk rbzero.tex_g0\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_44_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Left_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24233_ _04939_ _05016_ _05009_ _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_21445_ _02000_ _02530_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18153__I _11296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24164_ _04946_ _04947_ _04941_ _04948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_21376_ _02356_ _02366_ _02461_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22058__I0 rbzero.wall_tracer.rcp_fsm.o_data\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20327_ _12692_ _12919_ _13013_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_23115_ _03966_ _03971_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__24747__A2 _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24095_ _04874_ _04868_ _04871_ _04878_ _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XTAP_TAPCELL_ROW_112_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23046_ _03838_ _03877_ _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20258_ _12984_ _13029_ _13030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__22222__A3 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16437__A1 rbzero.vga_sync.vsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21430__A1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20189_ _12960_ _12961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_243_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26805_ _00715_ clknet_leaf_174_i_clk rbzero.tex_g1\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XPHY_EDGE_ROW_95_Left_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_204_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14999__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24997_ _05775_ _05780_ _05781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_162_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14750_ rbzero.tex_b0\[24\] _08499_ _08556_ _08557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_clkbuf_leaf_9_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26736_ _00646_ clknet_leaf_41_i_clk rbzero.pov.ready_buffer\[66\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20858__I _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23948_ _04747_ _04748_ _04736_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_153_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_161_i_clk clknet_5_10__leaf_i_clk clknet_leaf_161_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_212_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13701_ rbzero.tex_r0\[58\] _07511_ _07488_ _07512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26667_ _00577_ clknet_leaf_154_i_clk rbzero.tex_b0\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14681_ _07717_ _08381_ _08488_ _07258_ _08489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_212_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23879_ rbzero.wall_tracer.rcp_fsm.o_data\[-4\] _04689_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17232__I _10555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16420_ _09883_ _09884_ _09878_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25618_ _06340_ _06341_ _06402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13632_ _07442_ _07443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_156_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26598_ _00508_ clknet_leaf_42_i_clk rbzero.pov.spi_buffer\[67\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_16351_ rbzero.spi_registers.buf_texadd3\[5\] _09829_ _09834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25549_ _06035_ _06088_ _06282_ _06284_ _06333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_183_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13974__A2 _07139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13563_ _07372_ _07373_ _07059_ _07365_ _07374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_176_i_clk clknet_5_8__leaf_i_clk clknet_leaf_176_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__19587__C _12325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15302_ _07732_ _09031_ _09049_ _09036_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_183_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19070_ _08148_ rbzero.wall_tracer.rayAddendY\[9\] _11914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_214_i_clk_I clknet_5_6__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16282_ _09747_ _09782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_217_Right_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13494_ _07295_ _07303_ _07304_ _07305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_192_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18021_ rbzero.wall_tracer.trackDistX\[2\] _11165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_180_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27219_ _01124_ clknet_leaf_109_i_clk rbzero.wall_tracer.stepDistY\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15233_ _08997_ _08984_ _08998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14923__A1 _07433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18114__A1 rbzero.debug_overlay.playerY\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18114__B2 _10358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15164_ _08935_ _08942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14115_ _07915_ _07918_ _07922_ _07923_ _07924_ _07925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__24738__A2 _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19972_ _12712_ _12719_ _12744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15095_ _08810_ _08887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_238_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14151__A2 _07570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18923_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _11830_ _11831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14046_ rbzero.tex_r1\[8\] _07855_ _07856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_114_i_clk clknet_5_31__leaf_i_clk clknet_leaf_114_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_197_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_223_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21421__A1 _12780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18854_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] _11772_ _11776_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_219_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17805_ _10966_ rbzero.pov.ready_buffer\[59\] _10967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18785_ rbzero.tex_r1\[57\] rbzero.tex_r1\[56\] _11724_ _11725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15997_ _09566_ _09567_ _09565_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_237_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15651__A2 _09303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24910__A2 _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14948_ _06873_ _07101_ _07424_ _07225_ _08751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_129_i_clk clknet_5_13__leaf_i_clk clknet_leaf_129_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_17736_ _10921_ rbzero.pov.ready_buffer\[35\] _10922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_222_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20768__I _12594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_201_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14879_ rbzero.tex_b1\[38\] _08250_ _08685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17667_ _10873_ _10579_ _10868_ _10876_ _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_148_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19406_ _12177_ _12178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_159_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16618_ _10065_ _10066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17598_ _10830_ _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16549_ _08111_ _08098_ _10001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19337_ _12131_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_234_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24426__A1 _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23229__A2 _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19268_ rbzero.tex_b1\[16\] rbzero.tex_b1\[15\] _12088_ _12092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14914__A1 rbzero.tex_b1\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18219_ _11337_ _11360_ _11303_ _11120_ _11363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_19199_ _11131_ _12038_ _11329_ _11376_ _12043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_103_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21230_ _02315_ _02316_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21161_ _12237_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__21660__A1 _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14006__I _07804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_229_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20112_ _12409_ _12884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__19605__A1 rbzero.wall_tracer.size\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14142__A2 _07916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21092_ _02106_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14450__B _08220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20043_ _12750_ _12791_ _12815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24920_ _05703_ _05701_ _05704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__17092__A1 _10471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24851_ _05634_ _05635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_198_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23802_ _04637_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_24782_ _05561_ _05565_ _05566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_163_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21994_ _03016_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26521_ _00431_ clknet_leaf_56_i_clk rbzero.debug_overlay.vplaneY\[-1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23733_ _04575_ _04576_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20945_ rbzero.traced_texVinit\[5\] _01778_ _02033_ _02034_ _02035_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_221_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_93_i_clk clknet_5_24__leaf_i_clk clknet_leaf_93_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_26452_ _00362_ clknet_leaf_46_i_clk rbzero.debug_overlay.playerX\[-7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23664_ _04354_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_20876_ _01834_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_25403_ _06010_ _06187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22615_ _11131_ _12225_ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26383_ _00293_ clknet_leaf_247_i_clk rbzero.spi_registers.buf_texadd2\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23595_ _04447_ _11141_ _02767_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__18344__A1 _07179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25334_ _06117_ _06118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_12_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22546_ _11288_ _03449_ _03450_ rbzero.traced_texa\[-3\] _03451_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13708__A2 _07518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25265_ _06030_ _06041_ _06049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22477_ _03402_ _03407_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_161_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27004_ _00914_ clknet_leaf_200_i_clk rbzero.tex_g0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24216_ net60 _04997_ net68 _04999_ _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_162_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21428_ _02508_ _02513_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25196_ _05921_ _05980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19844__A1 _12556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16658__A1 _10015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_248_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_88_i_clk_I clknet_5_24__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21651__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24147_ _04787_ _04835_ _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclkbuf_leaf_31_i_clk clknet_5_22__leaf_i_clk clknet_leaf_31_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_21359_ _02312_ _02441_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24078_ _04852_ _04854_ _04860_ net49 _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13755__I _07486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15920_ _09506_ _09509_ _09505_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23029_ _03767_ _03759_ _03886_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__13892__A1 _07191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13892__B2 _07041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17083__A1 _10466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_i_clk clknet_5_19__leaf_i_clk clknet_leaf_46_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_129_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15851_ _09455_ _09456_ _09448_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14802_ _07601_ _08607_ _08608_ _08609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_18570_ _11586_ _11602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15782_ rbzero.spi_registers.buf_texadd3\[12\] _09398_ _09405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_243_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17521_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _10786_ _10787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14733_ rbzero.tex_b0\[39\] _08233_ _08540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26719_ _00629_ clknet_leaf_29_i_clk rbzero.pov.ready_buffer\[49\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17452_ rbzero.pov.spi_buffer\[68\] _10743_ _10740_ _10744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14664_ rbzero.tex_g1\[48\] _07460_ _08472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16403_ rbzero.spi_registers.buf_texadd3\[19\] _09863_ _09872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13615_ _07325_ _07348_ _07426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13947__A2 rbzero.map_overlay.i_mapdy\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17383_ rbzero.pov.spi_buffer\[50\] _10692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14595_ _07827_ _08399_ _08402_ _08403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_95_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18335__A1 _11462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19122_ rbzero.debug_overlay.facingY\[-7\] _10007_ _11966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16334_ _09806_ _09822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_216_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13546_ _07355_ _07356_ _07357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__24408__A1 _05186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_216_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19053_ _11904_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16897__A1 _10295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16265_ _09742_ _09769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13477_ _07287_ _07288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18004_ rbzero.wall_tracer.trackDistX\[7\] _11148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15216_ _08951_ _08984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16196_ rbzero.spi_registers.buf_texadd1\[15\] _09707_ _09717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15147_ _08926_ _08918_ _08927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21642__A1 _08099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14124__A2 _07932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19955_ _12715_ _12716_ _12726_ _12727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15078_ _07190_ _07191_ _07192_ _08870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_248_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14029_ _07541_ _07839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_18906_ rbzero.traced_texa\[8\] rbzero.texV\[8\] _11815_ _11818_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_19886_ rbzero.wall_tracer.visualWallDist\[0\] _12301_ _12656_ _12657_ _12658_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_18837_ _11759_ _11761_ _11762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_241_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18768_ _11715_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17719_ _10904_ _10632_ _10908_ _10910_ _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_19_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18699_ rbzero.tex_r1\[20\] rbzero.tex_r1\[19\] _11672_ _11676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_236_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_236_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_195_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22370__A2 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20730_ _01819_ _01820_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_19_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20661_ _12236_ _01744_ _01752_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_18_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18326__A1 _11456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14060__A1 rbzero.tex_r1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22400_ _03345_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23380_ _04134_ _04234_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20592_ _12403_ _01578_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18877__A2 rbzero.texV\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22331_ _11283_ _03264_ _03278_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14348__C1 _08157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25050_ _05787_ _05788_ _05834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22262_ _03110_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14363__A2 _08040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24001_ _04788_ _04789_ _04786_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_21213_ _02290_ _02300_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22193_ _03162_ _03164_ _03171_ _03109_ rbzero.wall_tracer.rcp_fsm.i_data\[4\] _03172_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_76_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21144_ rbzero.wall_tracer.visualWallDist\[10\] _01577_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_247_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14180__B _07976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25952_ _06637_ _06733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_21075_ _02162_ _02163_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_245_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20026_ _12682_ _12797_ _12798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24903_ _05298_ _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__25127__A2 _05905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25883_ _05120_ _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_225_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24834_ _05614_ _05615_ _05617_ _05618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_38_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23689__A2 _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24765_ _05497_ _05547_ _05548_ _05549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_107_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21977_ _03004_ _02998_ _03006_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_201_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26504_ _00414_ clknet_leaf_30_i_clk rbzero.debug_overlay.vplaneX\[-7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23716_ rbzero.wall_tracer.trackDistY\[-7\] _03043_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20928_ _12690_ _01469_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24696_ _05477_ _05478_ _05401_ _05462_ _05480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__24638__B2 _05351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23512__I _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26435_ _00345_ clknet_leaf_57_i_clk rbzero.wall_tracer.rayAddendY\[-4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23647_ _04408_ _04425_ _04423_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20859_ _12356_ _12358_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17510__I _10758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13400_ gpout0.hpos\[7\] _07210_ _07211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_25_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26366_ _00276_ clknet_leaf_5_i_clk rbzero.spi_registers.buf_texadd1\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14380_ _07980_ _08170_ _08189_ _08190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_23578_ _04364_ _04430_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_181_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25317_ _06063_ _06094_ _06100_ _06101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_187_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13331_ _07140_ _07141_ _07144_ _07145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__16879__A1 rbzero.pov.ready_buffer\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22529_ _03440_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23668__B _11134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26297_ _00207_ clknet_leaf_229_i_clk rbzero.spi_registers.buf_leak\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_16050_ _09606_ _09607_ _09603_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25248_ _05821_ _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13262_ _07046_ _07067_ _07069_ _07072_ _07075_ _07076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_84_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15001_ reg_gpout\[1\] _08802_ _07185_ _08803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20427__A2 _13023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25179_ _05912_ _05941_ _05943_ _05963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13193_ _07002_ _07006_ _07007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_103_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_248_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_209_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19740_ _12248_ _11070_ _12512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_198_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16952_ _07685_ _10364_ _10365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_194_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15903_ rbzero.spi_registers.buf_otherx\[0\] _09495_ _09496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19671_ _12439_ _12440_ _12442_ _12191_ _12443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_95_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16883_ _10295_ _10305_ _10306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_189_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19172__I _12015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16803__A1 _09462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18622_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _11629_ _11632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_216_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15834_ _08821_ _08852_ _09444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_3_1_0_i_clk_I clknet_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18553_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _11592_ _11593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_47_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15765_ _09391_ _09392_ _09384_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15205__I _08916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17504_ rbzero.tex_b0\[14\] rbzero.tex_b0\[13\] _10775_ _10777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_231_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_218_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_177_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14716_ _08517_ _08519_ _08521_ _08522_ _08285_ _08523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__20363__A1 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18484_ rbzero.tex_g1\[56\] rbzero.tex_g1\[55\] _11549_ _11553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15696_ _09339_ _09341_ _09337_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_185_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14647_ rbzero.tex_g1\[59\] _08300_ _08455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17435_ rbzero.pov.spi_buffer\[63\] _10731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14042__A1 _07589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18308__A1 _11444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20115__A1 _12471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14593__A2 _07845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14578_ _08382_ _08383_ _08385_ _07814_ _07648_ _08386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_17366_ rbzero.pov.spi_buffer\[46\] _10674_ _10671_ _10680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_231_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_231_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19105_ _08148_ rbzero.wall_tracer.rayAddendY\[10\] _11949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_16317_ rbzero.spi_registers.buf_texadd2\[21\] _09802_ _09808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13529_ _07339_ _07340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17297_ _10626_ _10619_ _10628_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16036__I _09595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_111_i_clk_I clknet_5_31__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16248_ _09755_ _09756_ _09750_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19036_ rbzero.tex_g0\[50\] rbzero.tex_g0\[49\] _11893_ _11895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24253__I _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19808__A1 rbzero.wall_tracer.size\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15542__A1 rbzero.spi_registers.buf_texadd0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24801__A1 _05388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16179_ _09703_ _09704_ _09700_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_58_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15096__B _08887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19938_ _12708_ _12709_ _12710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_227_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17047__A1 _08151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22040__A1 _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19869_ rbzero.wall_tracer.size\[8\] _12579_ _12171_ _12641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_71_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21900_ _08123_ _11064_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_22880_ _03733_ _03738_ _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_222_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_50_Left_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_36_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21831_ _11075_ _09921_ _02877_ _10071_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__21146__A3 _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23540__A1 _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24550_ _05098_ _05334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20354__A1 _12955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_21762_ _09945_ _02813_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24428__I _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23501_ _04352_ _04353_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20713_ rbzero.wall_tracer.visualWallDist\[7\] _01577_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_24481_ net80 _05264_ _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_175_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21693_ _11260_ _02729_ _02755_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26220_ _00130_ clknet_leaf_16_i_clk rbzero.spi_registers.texadd1\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23432_ _03860_ _04052_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20644_ _01687_ _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__14584__A2 _07597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26151_ _00061_ clknet_leaf_217_i_clk rbzero.map_overlay.i_mapdy\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23363_ _03862_ _04217_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20575_ _01567_ _01656_ _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_78_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25102_ _05846_ _05851_ _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_22314_ rbzero.wall_tracer.trackDistY\[2\] _03254_ _03271_ _03272_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_143_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26082_ _05022_ _06777_ _06831_ _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_171_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23294_ _04147_ _04148_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15785__I _09037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25033_ _05634_ _05812_ _05813_ _05817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__21606__A1 _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22245_ _12595_ _03210_ _03211_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__25348__A2 _06093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22176_ _03154_ _03157_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21127_ _12698_ _01981_ _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26984_ _00894_ clknet_leaf_170_i_clk rbzero.tex_g0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_109_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25935_ _06707_ _06714_ _06716_ _06695_ _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_21058_ _02146_ _12959_ _02020_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_109_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24571__A3 _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20009_ _12780_ _12693_ _12781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25866_ _06649_ _06650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13880_ rbzero.debug_overlay.playerX\[4\] _06867_ _07691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_199_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24817_ _05318_ _05323_ _05601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_193_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25797_ _05993_ _06580_ _06581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_122_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18389__I1 rbzero.tex_g1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15550_ _09208_ _09232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__20345__A1 _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24748_ _05439_ _05461_ _05472_ _05532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_139_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14501_ rbzero.tex_g0\[42\] _07600_ _08310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_194_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15481_ _09067_ _09182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24679_ _05408_ _05368_ _05462_ _05403_ _05400_ _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__18336__I _07214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25284__A1 _06051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22098__A1 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14432_ _07532_ _08241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17220_ _10543_ _10571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_42_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26418_ _00328_ clknet_leaf_18_i_clk rbzero.spi_registers.buf_texadd3\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_27398_ _01303_ clknet_leaf_80_i_clk rbzero.wall_tracer.stepDistX\[-4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14575__A2 _07807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14085__B _07808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_172_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17151_ rbzero.pov.spi_counter\[2\] rbzero.pov.spi_counter\[1\] _10517_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26349_ _00259_ clknet_leaf_2_i_clk rbzero.spi_registers.buf_texadd0\[17\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14363_ rbzero.debug_overlay.playerX\[-6\] _08040_ _08045_ _08172_ _08173_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_135_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput16 i_mode[0] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_64_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput27 i_vec_csb net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_135_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16102_ _09599_ _09646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13314_ rbzero.spi_registers.texadd2\[0\] _07036_ _07030_ rbzero.spi_registers.texadd1\[0\]
+ _07128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14327__A2 _08011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17082_ _08134_ _10466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_165_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14294_ rbzero.debug_overlay.vplaneY\[0\] _08104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16033_ _09515_ _09585_ _09594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13535__B1 _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13245_ gpout0.hpos\[2\] _07059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_123_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13176_ _06907_ _06913_ _06919_ _06926_ _06989_ _06990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_62_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_248_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_229_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24011__A2 _08813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17984_ _11102_ _11126_ _11128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_236_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22022__A1 _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19723_ _12494_ _12495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22321__I _09926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16935_ rbzero.pov.ready_buffer\[54\] _10169_ _10286_ _10350_ _10351_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_205_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13943__I rbzero.map_overlay.i_mapdy\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19654_ _12397_ _12426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16866_ _10288_ _10289_ _10290_ _10282_ _10291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18605_ rbzero.tex_r0\[44\] rbzero.tex_r0\[43\] _11618_ _11622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15817_ rbzero.spi_registers.texadd3\[21\] _09032_ _09431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_232_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19585_ rbzero.wall_tracer.visualWallDist\[-6\] _12197_ _12245_ _12357_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_177_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16797_ _10222_ _10223_ _10230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19630__I _12401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18536_ rbzero.tex_r0\[14\] rbzero.tex_r0\[13\] _11581_ _11583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15748_ rbzero.spi_registers.buf_texadd3\[3\] _09375_ _09380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_18467_ _11479_ _11543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15679_ rbzero.spi_registers.buf_texadd2\[9\] _09328_ _09329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17752__A2 rbzero.pov.ready_buffer\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17418_ rbzero.pov.spi_buffer\[59\] _10709_ _10718_ _10719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__22991__I _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14566__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18398_ _11504_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17349_ _10664_ _10666_ _10667_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_5_3__f_i_clk clknet_3_0_0_i_clk clknet_5_3__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_132_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20360_ _09901_ _01453_ _01454_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15819__B _09430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19019_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _11882_ _11885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_20291_ _12970_ _12972_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22030_ _02994_ _03031_ _03042_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_244_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_244_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15818__A2 _09118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_228_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_209_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22013__A1 _09925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22231__I _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23981_ _03158_ _04728_ _04774_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__17325__I _10542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25720_ _06484_ _06503_ _06504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_138_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22932_ _12733_ _03788_ _03789_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_78_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25651_ _06386_ _06390_ _06435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input19_I i_reg_csb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22863_ _02666_ _02671_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_168_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22316__A2 _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24602_ _05170_ net56 _05275_ _05165_ _05386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__19540__I _10289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21814_ rbzero.debug_overlay.vplaneX\[0\] _02845_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25582_ _06350_ _06356_ _06365_ _06366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__20327__A1 _12692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24158__I _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22794_ _03651_ _03652_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27321_ _01226_ clknet_leaf_115_i_clk rbzero.traced_texa\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24533_ _05297_ _05315_ _05274_ _05317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_78_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18156__I _11255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21745_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] _02799_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_241_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27252_ _01157_ clknet_leaf_99_i_clk rbzero.wall_tracer.visualWallDist\[-8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_19_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24464_ _05197_ _05173_ _05247_ _05248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_4_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21676_ _10346_ _02740_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26203_ _00113_ clknet_leaf_8_i_clk rbzero.spi_registers.texadd0\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23415_ _04154_ _04164_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27183_ _01088_ clknet_leaf_74_i_clk rbzero.wall_tracer.size_full\[-10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20627_ _01716_ _01718_ _01530_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_154_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24395_ _05159_ _05160_ _05179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19496__A2 _11076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26134_ _00044_ clknet_leaf_40_i_clk rbzero.pov.sclk_buffer\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23346_ _04199_ _03842_ _04085_ _04200_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__14309__A2 _08007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20558_ _01649_ _01650_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_85_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26065_ _02724_ _06833_ _06834_ _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_23277_ _04131_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_20489_ _01576_ _01581_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25016_ _05767_ _05799_ _05800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22228_ _11137_ _11377_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_218_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19715__I _12486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20802__A2 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22159_ _03125_ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__22004__A1 _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26967_ _00877_ clknet_leaf_109_i_clk rbzero.texV\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14981_ _06892_ _08779_ _08781_ _07153_ _08782_ _07046_ _08783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__13763__I _07507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13296__A2 _07108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14493__A1 rbzero.tex_g0\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16720_ net17 net16 _10161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25918_ _06699_ _06700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_199_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13932_ rbzero.map_overlay.i_mapdx\[4\] _07743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_199_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26898_ _00808_ clknet_leaf_136_i_clk rbzero.tex_r1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_242_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_236_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16651_ _09990_ _09928_ _10083_ _10097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_13863_ _07431_ _07667_ _07673_ _07674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25849_ _06615_ _06622_ _06624_ _06627_ _06629_ _06632_ _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_88_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15602_ _09269_ _09271_ _09267_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19370_ rbzero.tex_b1\[60\] rbzero.tex_b1\[59\] _12146_ _12150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16582_ rbzero.debug_overlay.vplaneY\[10\] _10032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_158_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13794_ _07593_ _07596_ _07598_ _07602_ _07604_ _07605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_215_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19184__A1 _11307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18321_ _11434_ _11450_ _10256_ _11455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15533_ _09208_ _09220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_151_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Left_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_139_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18252_ _11391_ _11394_ _11395_ _11396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_15464_ rbzero.spi_registers.buf_texadd0\[1\] _09165_ _09170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_211_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14415_ _08205_ _08213_ _08218_ _08223_ _08224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_93_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17203_ rbzero.pov.spi_buffer\[4\] _10558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__21818__A1 _10015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15395_ rbzero.spi_registers.buf_sky\[0\] _09119_ _09120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18183_ rbzero.map_overlay.i_otherx\[3\] _11320_ _11255_ rbzero.map_overlay.i_othery\[2\]
+ _11327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_71_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22086__A4 _07236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14346_ rbzero.debug_overlay.facingY\[-7\] _08156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17134_ rbzero.pov.ready_buffer\[7\] _10472_ _10505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17065_ _10452_ _10432_ _10453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_243_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14277_ rbzero.debug_overlay.facingX\[-5\] _08087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_90_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16016_ rbzero.spi_registers.buf_mapdy\[5\] _09572_ _09581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13228_ rbzero.spi_registers.texadd0\[23\] _07035_ _07038_ _07041_ _07042_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_228_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14720__A2 _08526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25980__A2 rbzero.wall_tracer.rcp_fsm.o_data\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_115_Left_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_237_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22794__A2 _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_226_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13159_ rbzero.texu_hot\[3\] _06949_ _06972_ _06973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17967_ rbzero.map_rom.f2 _11111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13673__I _07483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19706_ _12476_ _12477_ _12478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24687__B _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_209_i_clk_I clknet_5_7__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16918_ rbzero.debug_overlay.playerY\[-1\] _10335_ _10336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17898_ rbzero.debug_overlay.facingX\[-2\] _11001_ _11042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19637_ _12405_ _12406_ _12408_ _12409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_205_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16984__I _10373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16849_ _08175_ _10275_ _10276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_204_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_17__f_i_clk_I clknet_3_4_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_204_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17973__A2 _11099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19568_ _12339_ _12340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_149_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19175__A1 _11252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_124_Left_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18519_ _11573_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19499_ _12254_ _12271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_146_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21530_ _02609_ _02614_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14437__C _08245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14539__A2 _07894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15736__A1 rbzero.spi_registers.buf_texadd3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21461_ _12383_ _02546_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14009__I _07524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19478__A2 _11074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23200_ _04053_ _04055_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20412_ _12422_ _12519_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24180_ _04916_ _04936_ _04963_ _04849_ _04964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_161_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21392_ _02464_ _02477_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__18150__A2 _11291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23131_ _03984_ _03987_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20343_ _12303_ _01437_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Left_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_219_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23062_ _03791_ _03916_ _03917_ _03797_ _03918_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_3_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20274_ _01367_ _01368_ _13036_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22013_ _09925_ _11391_ _02981_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_179_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16464__A2 _09918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26821_ _00731_ clknet_leaf_178_i_clk rbzero.tex_g1\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23964_ rbzero.wall_tracer.rcp_fsm.operand\[-1\] _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_166_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26752_ _00662_ clknet_leaf_222_i_clk rbzero.vga_sync.vsync vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__19402__A2 _12173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25703_ _06459_ _06485_ _06486_ _06487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22915_ _03712_ _03719_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26683_ _00593_ clknet_leaf_26_i_clk rbzero.pov.ready_buffer\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23895_ _04709_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_224_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25487__A1 _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_142_Left_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25634_ _06392_ _06415_ _06417_ _06418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_22846_ _02661_ _02674_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25565_ _06271_ _06348_ _06349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22777_ _02647_ _02655_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24516_ _05299_ _05300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_27304_ _01209_ clknet_leaf_189_i_clk rbzero.row_render.texu\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21728_ _11344_ _11420_ _11119_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_25496_ _06278_ _06279_ _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16843__B _10214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27235_ _01140_ clknet_leaf_81_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24447_ _05029_ _05230_ _05231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_19_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21659_ _02726_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14200_ _07983_ _07996_ _08001_ _08009_ _08010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_0_191_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15180_ rbzero.spi_registers.spi_buffer\[9\] _08955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22473__A1 _07160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27166_ _01071_ clknet_leaf_59_i_clk rbzero.wall_tracer.rayAddendX\[-5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24378_ _05045_ _05158_ _05161_ _05056_ _05162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__22136__I _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_5_i_clk_I clknet_5_4__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18141__A2 _11282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14131_ rbzero.tex_r1\[53\] _07920_ _07941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_26117_ _00027_ clknet_leaf_3_i_clk rbzero.spi_registers.spi_buffer\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_158_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23329_ _04182_ _04183_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_27097_ _01007_ clknet_leaf_140_i_clk rbzero.tex_b1\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__24214__A2 _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26048_ _05242_ _06753_ _06820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22225__A1 _12163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21028__A2 _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14062_ _07594_ _07872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_120_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18870_ _11787_ _11788_ _11790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_167_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20787__A1 _12489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17821_ _10973_ rbzero.pov.ready_buffer\[65\] _10977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14466__A1 _08201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_210_i_clk_I clknet_5_7__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17752_ _10928_ rbzero.pov.ready_buffer\[41\] _10932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14964_ net24 _08749_ _08767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24300__B _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_221_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16703_ _10145_ _10131_ _10146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13915_ _07718_ _07723_ _07724_ _07725_ _07726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_226_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17683_ _10882_ rbzero.pov.ready_buffer\[17\] _10887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14895_ _08696_ _08697_ _08700_ _08564_ _07839_ _08701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_89_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19422_ _12169_ _12194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16634_ _10079_ _10080_ _10081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13846_ rbzero.tex_r0\[22\] _07420_ _07421_ _07657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_230_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19157__A1 _08149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19353_ _12140_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16565_ _10015_ _10016_ _10017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13777_ rbzero.tex_r0\[0\] _07579_ _07587_ _07588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_168_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18904__A1 _11779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22755__B _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22700__A2 _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18304_ _07254_ _06876_ _07251_ _11441_ _11442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_155_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15516_ rbzero.spi_registers.texadd0\[16\] _09206_ _09207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19284_ _12101_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_210_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20711__A1 _12705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16496_ _08118_ _09948_ _09951_ _09952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_45_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18235_ _11138_ _11378_ _11379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_5_21__f_i_clk clknet_3_5_0_i_clk clknet_5_21__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_183_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15447_ _09156_ _09157_ _09149_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22464__A1 _11462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18166_ rbzero.map_overlay.i_mapdy\[2\] _11308_ _11306_ _07756_ _11309_ _11310_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_15378_ rbzero.spi_registers.buf_leak\[3\] _09103_ _09106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_187_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17117_ rbzero.pov.ready_buffer\[1\] _10489_ _10494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_187_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14329_ rbzero.debug_overlay.vplaneX\[-8\] _08139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18097_ _11240_ _11213_ _11241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22216__A1 _11278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17048_ rbzero.pov.ready_buffer\[30\] _10434_ _10440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_241_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19632__A2 _11998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_206_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14499__I _07493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13617__B _07427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18999_ rbzero.tex_g0\[34\] rbzero.tex_g0\[33\] _11872_ _11874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_224_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20961_ _02048_ _02005_ _02049_ _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__14209__A1 _07713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13680__A2 _07484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14209__B2 _07698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22700_ _03560_ _01776_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23680_ _04524_ _03032_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_239_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20892_ _01981_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_198_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19148__A1 _08156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21125__I _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22631_ _03507_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25350_ _05948_ _06040_ _06134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_22562_ _11284_ _03455_ _03456_ rbzero.traced_texa\[4\] _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24301_ _05002_ _05003_ _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_63_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21513_ _02593_ _02597_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_146_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25281_ _06036_ _06065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22493_ _03411_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__24444__A2 _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27020_ _00930_ clknet_leaf_169_i_clk rbzero.tex_g0\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24232_ net78 _04997_ _04979_ _04999_ _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_133_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21258__A2 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21444_ _12647_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22455__A1 _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24163_ _04821_ _04824_ _04947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__16134__A1 _08843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21375_ _02335_ _02355_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_160_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_248_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23114_ _03967_ _03970_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_82_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22058__I1 rbzero.wall_tracer.stepDistY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20326_ _01406_ _01420_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_24094_ _04875_ _04865_ _04877_ _04878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_101_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14696__B2 _08502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23045_ _03775_ _03880_ _03901_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_12_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20257_ _13006_ _13028_ _13029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__20769__A1 _12236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16437__A2 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20188_ _12959_ _12960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_216_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26804_ _00714_ clknet_leaf_175_i_clk rbzero.tex_g1\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_32_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24996_ _05778_ _05779_ _05780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__24380__A1 _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26735_ _00645_ clknet_leaf_41_i_clk rbzero.pov.ready_buffer\[65\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_230_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23947_ rbzero.wall_tracer.rcp_fsm.i_data\[-5\] _04740_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_193_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13700_ _07418_ _07511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14680_ _08198_ _08484_ _08487_ _08488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23878_ _03000_ _04699_ _04700_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26666_ _00576_ clknet_leaf_154_i_clk rbzero.tex_b0\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_98_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_84_i_clk_I clknet_5_28__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13631_ _07321_ _07334_ _07442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_25617_ _06340_ _06341_ _06401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_22829_ _03684_ _03687_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_211_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14620__A1 _07608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26597_ _00507_ clknet_leaf_42_i_clk rbzero.pov.spi_buffer\[66\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_196_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22694__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16350_ _09830_ _09832_ _09833_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13562_ _06877_ _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_109_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25548_ _06278_ _06279_ _06332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_55_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_181_Right_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15301_ rbzero.spi_registers.buf_othery\[4\] _09038_ _09049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16281_ rbzero.spi_registers.buf_texadd2\[12\] _09780_ _09781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25479_ _06261_ _06255_ _06257_ _06259_ _06262_ _06263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_54_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16373__A1 rbzero.spi_registers.spi_buffer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13493_ _07288_ _07289_ _07304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18020_ rbzero.wall_tracer.trackDistY\[3\] _11164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_27218_ _01123_ clknet_leaf_110_i_clk rbzero.wall_tracer.stepDistY\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__14805__C _07478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15232_ rbzero.spi_registers.spi_buffer\[18\] _08997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_125_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_229_Left_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_180_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__18114__A2 _11255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15163_ _08939_ _08940_ _08941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27149_ _01054_ clknet_leaf_182_i_clk reg_rgb\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__26562__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24199__A1 _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14114_ _07526_ _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_19971_ _12712_ _12719_ _12743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15094_ rbzero.spi_registers.buf_vinf _08885_ _08886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16799__I _10231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14045_ _07599_ _07855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18922_ _11829_ _11830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_120_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_223_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18853_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] _11775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_246_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17804_ _10856_ _10966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_237_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18784_ _11713_ _11724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_238_Left_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15996_ _08983_ _09562_ _09567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_222_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17735_ _10905_ _10921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14947_ _07988_ _08750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_82_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18050__A1 _11190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_201_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17666_ _10875_ rbzero.pov.ready_buffer\[11\] _10876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14878_ _08680_ _08681_ _08682_ _08683_ _08346_ _08684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_19405_ _12176_ _12177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16617_ _10032_ _10065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13829_ rbzero.tex_r0\[31\] _07626_ _07640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17597_ rbzero.tex_b0\[54\] rbzero.tex_b0\[53\] _10828_ _10830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__25871__A1 _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19336_ rbzero.tex_b1\[45\] rbzero.tex_b1\[44\] _12130_ _12131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22685__A1 _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16548_ _09983_ _09985_ _09999_ _10000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_18_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_234_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19267_ _12091_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_247_Left_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_16479_ _09933_ _09914_ _09935_ _09936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18218_ _11338_ _11360_ _11340_ _11331_ _11361_ _11362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_171_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19198_ _11131_ _12039_ _12041_ _12042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__14914__A2 _08526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18149_ rbzero.wall_tracer.visualWallDist\[0\] _11293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16116__A1 rbzero.spi_registers.buf_texadd0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17864__A1 rbzero.debug_overlay.facingX\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21160_ _02107_ _02124_ _02247_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__21660__A2 _08741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14678__A1 _08485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20111_ _12625_ _12880_ _12881_ _12882_ _12883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xclkbuf_leaf_221_i_clk clknet_5_3__leaf_i_clk clknet_leaf_221_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_21091_ _02057_ _02126_ _02162_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13350__A1 _07147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20042_ _12812_ _12813_ _12814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13350__B2 _07150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19813__I _12584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14022__I _07831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24850_ _05632_ _05633_ _05634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_147_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_236_i_clk clknet_5_6__leaf_i_clk clknet_leaf_236_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_23801_ _11162_ _04636_ _04586_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_106_i_clk_I clknet_5_30__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24781_ _05562_ _05563_ _05564_ _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_21993_ rbzero.wall_tracer.rcp_fsm.o_data\[4\] rbzero.wall_tracer.size_full\[4\]
+ _02985_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_225_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23732_ rbzero.wall_tracer.trackDistY\[-5\] _03048_ _04571_ _04576_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26520_ _00430_ clknet_leaf_56_i_clk rbzero.debug_overlay.vplaneY\[-2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20944_ _10071_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23663_ _11141_ _04351_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26451_ _00361_ clknet_leaf_46_i_clk rbzero.debug_overlay.playerX\[-8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20875_ _01963_ _01964_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14602__B2 _07861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25402_ _06185_ _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22614_ _03481_ _03490_ _03497_ _10049_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_193_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26382_ _00292_ clknet_leaf_247_i_clk rbzero.spi_registers.buf_texadd2\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23594_ _02761_ _04355_ _04446_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13956__A3 _07697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25333_ _05869_ _05909_ _06117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_12_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22545_ _03437_ _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18164__I _11255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16355__A1 _08939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25264_ _06036_ _06047_ _06048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22476_ _07153_ _03405_ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14905__A2 _07561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24215_ _04961_ _04962_ _04998_ _04999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_32_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27003_ _00913_ clknet_leaf_200_i_clk rbzero.tex_g0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_72_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21427_ _02509_ _02512_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16107__A1 _08994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25195_ _05977_ _05978_ _05979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24146_ _04833_ _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__17855__A1 rbzero.debug_overlay.facingX\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21358_ _02308_ _02443_ _02444_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14641__B _07917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14669__A1 _07480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_248_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20309_ _13006_ _13028_ _01403_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24077_ _04761_ _04856_ _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_21289_ _02374_ _02375_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_164_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23028_ _03882_ _03885_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_217_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22600__A1 _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13892__A2 _07698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17083__A2 _10443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15850_ _08942_ _09445_ _09456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_189_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24353__A1 _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14801_ rbzero.tex_b0\[7\] _08209_ _08608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15781_ rbzero.spi_registers.texadd3\[12\] _09396_ _09404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24979_ net43 _05762_ _05763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13771__I _07481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17243__I _10564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18032__A1 _11173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17520_ _10780_ _10786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_203_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18032__B2 _11175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14732_ _07609_ _08533_ _08538_ _08539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_26718_ _00628_ clknet_leaf_29_i_clk rbzero.pov.ready_buffer\[48\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_142_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21962__I0 rbzero.wall_tracer.rcp_fsm.o_data\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17451_ _10543_ _10743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14663_ _08467_ _08468_ _08470_ _08459_ _07464_ _08471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_26649_ _00559_ clknet_leaf_146_i_clk rbzero.tex_b0\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_200_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19598__C _12369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16402_ _09870_ _09871_ _09867_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_200_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13614_ _06858_ _07424_ _06882_ _07425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_95_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17382_ _10690_ _10688_ _10691_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_223_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14594_ _07842_ _08400_ _08401_ _08402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_45_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19121_ _11962_ _11963_ _11964_ _11965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16333_ rbzero.spi_registers.spi_buffer\[0\] _09820_ _09821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13545_ rbzero.row_render.size\[6\] _07356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_125_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25605__A1 _05977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_216_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_216_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19052_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _11903_ _11904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13476_ rbzero.texV\[4\] _07285_ _07286_ _07287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16264_ _09767_ _09768_ _09762_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16897__A2 _10317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18003_ rbzero.wall_tracer.trackDistX\[8\] _11147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_35_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15215_ rbzero.spi_registers.spi_buffer\[15\] _08983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14107__I _07520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16195_ _09715_ _09716_ _09712_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17846__A1 _10845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15146_ rbzero.spi_registers.spi_buffer\[4\] _08926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_19954_ _12714_ _12717_ _12726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_15077_ _07988_ _08751_ _08869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_77_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13332__A1 _07061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14028_ _07825_ _07838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18905_ rbzero.traced_texa\[8\] rbzero.texV\[8\] _11817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19885_ _10336_ _12006_ _12169_ _12657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_18836_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] _11761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_184_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_208_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24344__A1 _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23147__A2 _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16478__B _09934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18767_ rbzero.tex_r1\[49\] rbzero.tex_r1\[48\] _11714_ _11715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15979_ rbzero.spi_registers.buf_mapdx\[1\] _09548_ _09554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_234_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_222_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17718_ _10906_ rbzero.pov.ready_buffer\[29\] _10910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_19_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22994__I _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20905__A1 _12668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18698_ _11675_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_236_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_236_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17649_ _10859_ rbzero.pov.ready_buffer\[6\] _10864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24647__A2 _05406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22658__A1 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20660_ _01746_ _01751_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_147_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14060__A2 _07829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19319_ _12121_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_190_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16337__A1 _08913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20133__A2 _12587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20591_ _12398_ _01682_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22330_ _03283_ _03275_ _03284_ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__14348__B1 _08045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14348__C2 _08035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14899__A1 rbzero.tex_b1\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22261_ _11197_ _03226_ _03227_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14017__I _07449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15560__A2 _09232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24000_ rbzero.wall_tracer.rcp_fsm.i_data\[7\] _04773_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_32_i_clk_I clknet_5_22__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21212_ _02293_ _02299_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_160_i_clk clknet_5_10__leaf_i_clk clknet_leaf_160_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__17837__A1 _10845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22192_ _03165_ _03170_ _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22234__I _11248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21143_ _12969_ _01916_ _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_247_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13323__A1 _07045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25951_ _06668_ _06732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_21074_ _02127_ _02161_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19543__I _12314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_175_i_clk clknet_5_8__leaf_i_clk clknet_leaf_175_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_20025_ _12703_ _12712_ _12718_ _12797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_24902_ _05650_ _05680_ _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__17065__A2 _10432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25882_ _06663_ _06664_ _06665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24335__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24833_ _05616_ _05606_ _05608_ _05617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_21976_ rbzero.wall_tracer.size\[5\] _03005_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24764_ _05499_ _05541_ _05548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_107_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26503_ _00413_ clknet_leaf_30_i_clk rbzero.debug_overlay.vplaneX\[-8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23715_ _11198_ _04554_ _04561_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20927_ _02016_ _12958_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24695_ _05477_ _05478_ _05479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15379__A2 _09106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26434_ _00344_ clknet_leaf_51_i_clk rbzero.wall_tracer.rayAddendY\[-5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20858_ _01947_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23646_ _04475_ _04491_ _04497_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_138_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_113_i_clk clknet_5_31__leaf_i_clk clknet_leaf_113_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23577_ _04394_ _04429_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26365_ _00275_ clknet_leaf_17_i_clk rbzero.spi_registers.buf_texadd1\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20789_ _01874_ _01879_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_135_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13330_ _07142_ _07143_ _07144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22528_ _12595_ _03436_ _03438_ rbzero.traced_texa\[-10\] _03440_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_25316_ _06074_ _06098_ _06099_ _06100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__16879__A2 _10252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26296_ _00206_ clknet_leaf_229_i_clk rbzero.spi_registers.buf_leak\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15000__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13261_ _07053_ _06996_ _07073_ _07074_ _07075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_25247_ _06030_ _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22459_ _03361_ _03398_ _03399_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15551__A2 _09232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_128_i_clk clknet_5_13__leaf_i_clk clknet_leaf_128_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15000_ net86 _08793_ _08801_ _08802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25178_ _05912_ _05941_ _05962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13192_ rbzero.spi_registers.texadd0\[18\] _07003_ _07005_ _07006_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13766__I _07576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24129_ _04724_ _04912_ _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16142__I _09660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_248_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16951_ _10266_ _10360_ _10314_ _10364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__21388__A1 _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19453__I _12194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18253__A1 _09925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17056__A2 _10445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15902_ _09494_ _09495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19670_ rbzero.debug_overlay.playerX\[-3\] _11095_ _12441_ _12157_ _12442_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_144_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16882_ _10303_ _10304_ _10305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__24326__A1 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18621_ _11631_ _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15833_ _08827_ _09443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24877__A2 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18552_ _11586_ _11592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_231_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15764_ rbzero.spi_registers.buf_texadd3\[7\] _09387_ _09392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17503_ _10776_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__18800__I0 _07171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14715_ _07613_ _08522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18483_ _11552_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_218_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21560__A1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15695_ rbzero.spi_registers.buf_texadd2\[13\] _09340_ _09341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_5_0_i_clk_I clknet_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17434_ _10728_ _10724_ _10730_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14646_ _07889_ _08441_ _08453_ _08454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18308__A2 _08788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17365_ rbzero.pov.spi_buffer\[45\] _10679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_126_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20115__A2 _12885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14577_ rbzero.tex_g1\[20\] _07810_ _08384_ _08385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_231_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19104_ _11916_ _11947_ _11914_ _11948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_16316_ _09803_ _09805_ _09807_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13528_ _07321_ _07338_ _07339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17296_ rbzero.pov.spi_buffer\[28\] _10627_ _10624_ _10628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19035_ _11894_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16247_ _08922_ _09748_ _09756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13459_ _07269_ _07270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__19808__A2 _12514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16178_ _08959_ _09698_ _09704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13676__I _07486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15129_ _08911_ _08912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_92_i_clk clknet_5_24__leaf_i_clk clknet_leaf_92_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_229_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19937_ _12356_ _12358_ _12361_ _12192_ _12709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__17047__A2 _10432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19868_ rbzero.wall_tracer.size\[8\] _12579_ _12640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_71_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18819_ _11738_ _11747_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19799_ _12276_ _12570_ _12497_ _12502_ _12571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_223_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21830_ _02875_ _02876_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21761_ _10455_ _08140_ _08144_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_148_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_i_clk clknet_5_22__leaf_i_clk clknet_leaf_30_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_20712_ _01682_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_23500_ _04245_ _04246_ _04249_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24480_ _05033_ _05260_ _05262_ _05263_ _05264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_176_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21692_ _12046_ _02754_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25968__C _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23431_ _04219_ _04050_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20643_ _01709_ _01734_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_190_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer41_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26150_ _00060_ clknet_leaf_217_i_clk rbzero.map_overlay.i_mapdx\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23362_ _02079_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20574_ _01562_ _01566_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_45_i_clk clknet_5_16__leaf_i_clk clknet_leaf_45_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25101_ _05854_ _05855_ _05885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22313_ _11165_ _03270_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19538__I _12255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26081_ _06811_ _06803_ _06804_ _06662_ _06847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_61_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23293_ _04031_ _04045_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25032_ _05808_ _05814_ _05815_ _05816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_104_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22244_ _11209_ _03204_ _03213_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21606__A2 _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17058__I _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22175_ rbzero.wall_tracer.rcp_fsm.i_data\[1\] _03144_ _03156_ _03157_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_5_6__f_i_clk_I clknet_3_1_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21126_ _12685_ _02213_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__24556__A1 _05292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26983_ _00893_ clknet_leaf_171_i_clk rbzero.tex_g0\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13847__A2 _07576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25934_ _06696_ _06715_ _06716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21057_ _02016_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_109_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24308__A1 _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20008_ _12779_ _12780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25865_ _05091_ _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_202_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24816_ _05323_ _05600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25796_ _05976_ _05989_ _05992_ _06580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_186_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_122_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19735__A1 _12384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24747_ _05526_ _05530_ _05531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21959_ rbzero.wall_tracer.rcp_fsm.o_data\[-8\] _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_159_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14500_ rbzero.tex_g0\[43\] _07898_ _08309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15480_ rbzero.spi_registers.buf_texadd0\[6\] _09137_ _09181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24678_ _05439_ _05461_ _05393_ _05462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__25878__C _10992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14431_ rbzero.tex_g0\[6\] _08227_ _08240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26417_ _00327_ clknet_leaf_18_i_clk rbzero.spi_registers.buf_texadd3\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23629_ _04384_ _04389_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27397_ _01302_ clknet_leaf_76_i_clk rbzero.wall_tracer.stepDistX\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_42_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_213_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17150_ _10512_ _10516_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20882__I _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_172_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26348_ _00258_ clknet_leaf_2_i_clk rbzero.spi_registers.buf_texadd0\[16\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14362_ rbzero.debug_overlay.playerX\[-7\] _08172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 i_mode[1] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput28 i_vec_mosi net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16101_ rbzero.spi_registers.buf_texadd0\[16\] _09644_ _09645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_137_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13313_ _06981_ _07127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14293_ _08102_ _08103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17081_ _10447_ _10464_ _10465_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_220_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26279_ _00189_ clknet_leaf_244_i_clk rbzero.spi_registers.texadd3\[22\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16721__A1 _08875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24795__A1 _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16032_ rbzero.spi_registers.buf_mapdyw\[1\] _09583_ _09593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13244_ _07048_ _07051_ _07055_ _07019_ _07057_ _07058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_122_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13175_ _06929_ _06988_ _06989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_150_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17521__I0 rbzero.tex_b0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15288__A1 _07721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15827__A3 _08843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17983_ _11102_ _11126_ _11127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_229_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19722_ _12355_ _12357_ _12360_ _12494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_179_Left_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__18226__A1 _11107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16934_ _10238_ _10348_ _10349_ _10350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_236_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16600__I _10048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25913__I _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19653_ _12398_ _12403_ _12414_ _12424_ _12425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_217_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16865_ rbzero.pov.ready_buffer\[45\] _10274_ _10290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__26010__S _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19911__I _12489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15216__I _08951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18604_ _11621_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14120__I _07498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15816_ _09426_ _09427_ _09430_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19026__I0 rbzero.tex_g0\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19584_ _12355_ _12356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_88_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16796_ _10164_ _10229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_172_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18535_ _11582_ _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15747_ rbzero.spi_registers.texadd3\[3\] _09373_ _09379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18466_ _11542_ _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15678_ _09305_ _09328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15212__A1 _08980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_188_Left_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17417_ _10705_ _10718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22089__A2 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14629_ rbzero.tex_g1\[38\] _07898_ _07819_ _08437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18397_ rbzero.tex_g1\[18\] rbzero.tex_g1\[17\] _11502_ _11504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16960__A1 _08066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17348_ rbzero.pov.spi_buffer\[41\] _10662_ _10659_ _10667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_205_i_clk_I clknet_5_18__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17279_ _10602_ _10615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19018_ _11884_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_20290_ _12970_ _12972_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19662__B1 _12430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_197_Left_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_244_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_244_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22512__I _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13829__A2 _07626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_209_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_209_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22013__A2 _11391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23980_ _04772_ _04773_ _09113_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__23210__B2 _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19965__A1 _12305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23761__A2 _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22931_ _02600_ _03788_ _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19821__I _12592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25650_ _06395_ _06432_ _06433_ _06434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_22862_ _03710_ _03720_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_88_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15451__A1 rbzero.spi_registers.vshift\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24601_ _05347_ _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_88_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21813_ rbzero.debug_overlay.vplaneX\[0\] _02845_ _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25581_ _06357_ _06364_ _06365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22793_ _02349_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_189_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27320_ _01225_ clknet_leaf_115_i_clk rbzero.traced_texa\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24532_ _05297_ _05274_ _05315_ _05316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_21744_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] _02798_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_164_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15203__A1 _08973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27251_ _01156_ clknet_leaf_99_i_clk rbzero.wall_tracer.visualWallDist\[-9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24463_ _05214_ _05174_ _05176_ _05099_ _05247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_21675_ _02739_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_188_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26202_ _00112_ clknet_leaf_8_i_clk rbzero.spi_registers.texadd0\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20626_ _01528_ _01717_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23414_ _04266_ _04188_ _04267_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_184_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27182_ _01087_ clknet_leaf_74_i_clk rbzero.wall_tracer.size_full\[-11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24394_ _05173_ _05177_ _05075_ _05178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_154_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23345_ _04084_ _04087_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26133_ _00043_ clknet_leaf_213_i_clk rbzero.pov.sclk_buffer\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16703__A1 _10145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20557_ _12209_ _01478_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_119_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26064_ _04799_ rbzero.wall_tracer.rcp_fsm.o_data\[3\] _06834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_23276_ _04115_ _04118_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20488_ _12675_ _01580_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22227_ _11392_ _03196_ _03198_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25015_ _05770_ _05798_ _05799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14190__A1 _06888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22158_ _03140_ _03143_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_160_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21109_ _12731_ _01967_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__18208__B2 _11112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26966_ _00876_ clknet_leaf_110_i_clk rbzero.texV\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_22089_ _03081_ _03082_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_14980_ net9 _08780_ _08782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_22_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14493__A2 _08298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25917_ _05214_ _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_199_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13931_ rbzero.map_overlay.i_mapdx\[3\] rbzero.map_overlay.i_mapdx\[2\] _07741_ _07737_
+ _07742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_26897_ _00807_ clknet_leaf_136_i_clk rbzero.tex_r1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_214_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_1_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16650_ _10090_ _10095_ _10096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25848_ _06631_ _06632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__20877__I _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13862_ rbzero.color_floor\[0\] _07669_ _07670_ _07672_ _07673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_199_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_154_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15601_ rbzero.spi_registers.buf_texadd1\[13\] _09270_ _09271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16581_ _10030_ _10031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25779_ _06480_ _06523_ _06563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21515__A1 _12789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13793_ _07603_ _07604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_85_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17251__I _10571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18320_ _11434_ _11449_ _08871_ _11445_ _11454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_186_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15532_ rbzero.spi_registers.texadd0\[20\] _09218_ _09219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_139_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18251_ _11137_ _11390_ _11395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_139_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27449_ _01354_ clknet_leaf_71_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__23268__A1 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15463_ rbzero.spi_registers.texadd0\[1\] _09163_ _09169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15745__A2 _09375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17202_ _10554_ _10545_ _10557_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14414_ _08219_ _08221_ _08222_ _08223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_210_Left_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18182_ rbzero.map_overlay.i_otherx\[1\] _11315_ _11106_ _09027_ _11326_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_15394_ _09118_ _09119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17133_ _10503_ _10504_ _10492_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_14345_ rbzero.debug_overlay.facingY\[-6\] _08155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__25908__I _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17064_ _08140_ _10452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14276_ _08084_ _08035_ _08040_ _08085_ _08086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_90_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16015_ _09579_ _09580_ _09576_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_79_i_clk_I clknet_5_30__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13227_ _07040_ _07041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_55_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13158_ _06951_ _06971_ _06972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_237_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_226_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13089_ rbzero.wall_tracer.rcp_fsm.i_start _06895_ _06900_ _06903_ _00004_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_17966_ _11109_ _11101_ _11110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_237_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20006__A1 _12777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14484__A2 _08288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19705_ _12412_ _12477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16917_ _07704_ _10330_ _10335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17897_ _11040_ _11032_ _11041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__20557__A2 _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19636_ rbzero.debug_overlay.playerX\[-4\] _11096_ _12407_ _12158_ _12408_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_16848_ _10181_ _10275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_189_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_195_Right_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_205_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_204_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19567_ rbzero.wall_tracer.visualWallDist\[-7\] _12197_ _12245_ _12339_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_177_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20309__A2 _13028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16779_ _10211_ _10213_ _10214_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18518_ rbzero.tex_r0\[6\] rbzero.tex_r0\[5\] _11571_ _11573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__19175__A2 _12007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19498_ rbzero.wall_tracer.size\[2\] _12247_ _12269_ _12166_ _12270_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_76_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18449_ _11522_ _11533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_34_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16933__A1 _10346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_248_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_21460_ _01469_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_209_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20411_ _12884_ _12379_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21391_ _02471_ _02476_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23130_ _03985_ _03986_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__18150__A3 _11292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20342_ _01436_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23061_ _03790_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20273_ _01366_ _13034_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_102_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25039__B _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22012_ _03028_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17110__A1 _09915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26820_ _00730_ clknet_leaf_180_i_clk rbzero.tex_g1\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_209_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26751_ _00661_ clknet_leaf_121_i_clk rbzero.wall_tracer.mapX\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23963_ _04759_ _04760_ _04752_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_243_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25702_ _06448_ _06458_ _06486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22914_ _01905_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_242_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26682_ _00592_ clknet_leaf_26_i_clk rbzero.pov.ready_buffer\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23894_ rbzero.wall_tracer.rcp_fsm.o_data\[3\] _01699_ _04693_ _04709_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_211_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_162_Right_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25633_ _06416_ _06365_ _06417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_168_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22845_ _02661_ _02674_ _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14695__I _07808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25564_ _06143_ _06346_ _06347_ _06348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_182_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22776_ _02649_ _02654_ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27303_ _01208_ clknet_leaf_190_i_clk rbzero.row_render.texu\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24515_ _05268_ net69 _05299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_164_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21727_ _11134_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25495_ _06035_ _06006_ _06156_ _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__16924__A1 _08018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27234_ _01139_ clknet_leaf_84_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24446_ net69 _05207_ _05219_ _05229_ _05230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_137_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21658_ _02724_ _08628_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20609_ _01699_ _12445_ _01700_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_27165_ _01070_ clknet_leaf_205_i_clk rbzero.wall_tracer.mapX\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24377_ _05105_ _05106_ _05159_ _05160_ _05161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_21589_ _02662_ _02673_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__23670__A1 _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22473__A2 _08750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18141__A3 _11283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14130_ _07515_ _07940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26116_ _00026_ clknet_leaf_3_i_clk rbzero.spi_registers.spi_buffer\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23328_ _04062_ _04059_ _04064_ _01744_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_27096_ _01006_ clknet_leaf_141_i_clk rbzero.tex_b1\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_50_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_80_i_clk_I clknet_5_30__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14163__A1 _07775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26047_ _06739_ _06633_ _06818_ _06819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__22225__A2 _11394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14061_ rbzero.tex_r1\[5\] _07832_ _07587_ _07871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23259_ _04016_ _04114_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17820_ _10972_ _10734_ _10975_ _10976_ _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_219_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19929__A1 _12334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19929__B2 _12700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23725__A2 _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17751_ _10927_ _10664_ _10930_ _10931_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_26949_ _00859_ clknet_leaf_181_i_clk rbzero.tex_r1\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14963_ net41 _08760_ _08766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_180_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16702_ _09990_ _10145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_221_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13914_ _07226_ rbzero.map_overlay.i_othery\[3\] _07725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_180_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17682_ _10881_ _10593_ _10885_ _10886_ _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_187_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14894_ rbzero.tex_b1\[42\] _08698_ _08699_ _08700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_199_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19421_ _12192_ _12193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16633_ _10059_ _10058_ _10056_ _10080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_230_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13845_ rbzero.tex_r0\[23\] _07591_ _07656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19352_ rbzero.tex_b1\[52\] rbzero.tex_b1\[51\] _12136_ _12140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16564_ _10009_ _10010_ _10013_ _10016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_230_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13776_ _07586_ _07587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22161__A1 _11986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18303_ _07139_ _07160_ _06859_ _07149_ _11441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_242_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15515_ _09205_ _09206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19283_ rbzero.tex_b1\[22\] rbzero.tex_b1\[21\] _12099_ _12101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16495_ _08111_ rbzero.wall_tracer.rayAddendY\[-4\] _09950_ _09951_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_57_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16915__A1 _07704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18234_ _11248_ _11377_ _11378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13729__A1 rbzero.tex_r0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15446_ rbzero.spi_registers.buf_vshift\[2\] _09154_ _09157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18165_ rbzero.map_overlay.i_mapdy\[1\] _11252_ _11309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_167_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15377_ rbzero.floor_leak\[3\] _09101_ _09105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17116_ _09933_ _10487_ _10493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_187_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14328_ rbzero.debug_overlay.vplaneX\[-1\] _08138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18096_ rbzero.wall_tracer.trackDistY\[-11\] _11240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_208_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17047_ _08151_ _10432_ _10439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14259_ _08057_ _08058_ _08060_ _08061_ _08068_ _08069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_241_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13684__I _07444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25166__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_206_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18998_ _11873_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_224_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14457__A2 _07584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23716__A2 _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17949_ _08076_ _11092_ _11093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_206_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20960_ _01905_ _01994_ _02006_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__16928__C _10221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14209__A2 _08007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19619_ _12373_ _12390_ _12391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_221_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20891_ rbzero.wall_tracer.stepDistX\[8\] _12445_ _01980_ _01981_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_177_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_239_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15404__I _09067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22630_ rbzero.wall_tracer.texu\[5\] rbzero.texu_hot\[5\] _03503_ _03507_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_221_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22561_ _03459_ _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16906__A1 _07706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24300_ _05076_ _05081_ _05083_ _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_21512_ _02594_ _02596_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_63_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25280_ _06053_ _06056_ _06064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22492_ _03409_ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_161_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24231_ _05014_ _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_21443_ _02409_ _02403_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_151_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16235__I _09746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_102_i_clk_I clknet_5_27__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24162_ _04874_ _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24452__I _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21374_ _02370_ _02395_ _02368_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16134__A2 _09669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20325_ _01414_ _01419_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_23113_ _03968_ _03969_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_24093_ _04746_ _04876_ _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_31_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23044_ _03776_ _03879_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_112_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_231_Right_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20256_ _13009_ _13011_ _13027_ _13028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__23955__A2 _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21966__A1 rbzero.wall_tracer.size\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20187_ _12958_ _12959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14448__A2 _08202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26803_ _00713_ clknet_leaf_168_i_clk rbzero.tex_g1\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24995_ _05304_ net91 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__21718__A1 _11338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26734_ _00644_ clknet_leaf_41_i_clk rbzero.pov.ready_buffer\[64\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23946_ _04746_ _04743_ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_162_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22391__A1 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26665_ _00575_ clknet_leaf_154_i_clk rbzero.tex_b0\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA_clkbuf_leaf_27_i_clk_I clknet_5_20__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23877_ rbzero.wall_tracer.stepDistX\[-5\] _04694_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_212_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25616_ _06339_ _06400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13959__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13630_ _07434_ _07440_ _07441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_22828_ _03685_ _03686_ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__21760__B _10455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24627__I _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22143__A1 rbzero.wall_tracer.visualWallDist\[-5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26596_ _00506_ clknet_leaf_42_i_clk rbzero.pov.spi_buffer\[65\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22143__B2 _11074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14620__A2 _08427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25547_ _06297_ _06305_ _06331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13561_ rbzero.row_render.size\[3\] _07372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__18898__A1 rbzero.traced_texa\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22759_ _11165_ rbzero.wall_tracer.stepDistX\[2\] _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_137_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15300_ _09047_ _09048_ _09042_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16280_ _09742_ _09780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25478_ _06203_ _06209_ _06249_ _06254_ _06262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_13492_ _07301_ _07302_ _07303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_81_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27217_ _01122_ clknet_leaf_75_i_clk rbzero.wall_tracer.stepDistY\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__14384__A1 _07222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15231_ rbzero.spi_registers.spi_buffer\[19\] _08992_ _08996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24429_ _05209_ _05211_ _05124_ _05053_ _05126_ _05212_ _05213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_180_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14093__C _07638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15162_ _08917_ _08940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_27148_ _01053_ clknet_leaf_182_i_clk reg_rgb\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14113_ _07546_ _07923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19970_ _12741_ _12742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15093_ _08884_ _08885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_27079_ _00989_ clknet_leaf_153_i_clk rbzero.tex_b1\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__23946__A2 _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18921_ _11828_ _11829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14044_ _07803_ _07815_ _07828_ _07840_ _07853_ _07854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_197_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_223_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_182_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_18852_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] _11774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25193__I _05948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17803_ _10848_ _10965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18783_ _11723_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15995_ rbzero.spi_registers.buf_mapdx\[5\] _09560_ _09566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_222_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17734_ _10903_ _10920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_222_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24371__A2 _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14946_ net5 _08748_ _08749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_238_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_17665_ _10874_ _10875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_201_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14877_ rbzero.tex_b1\[33\] _08541_ _08497_ _08683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_214_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25320__A1 _05977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19404_ _12175_ _12176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16616_ _10032_ _10063_ _10064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13828_ _07627_ _07631_ _07634_ _07637_ _07638_ _07639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_203_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17596_ _10829_ _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14611__A2 _07832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16547_ _08110_ rbzero.debug_overlay.vplaneY\[-9\] _09999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19335_ _12114_ _12130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__18889__A1 _11769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13759_ _07348_ _07570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_63_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19266_ rbzero.tex_b1\[15\] rbzero.tex_b1\[14\] _12088_ _12091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16478_ _09933_ _09914_ _09934_ _09935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18217_ _11263_ _11354_ _11361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_170_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15429_ rbzero.spi_registers.buf_floor\[4\] _09131_ _09144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14375__A1 _07677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19197_ _09895_ _12040_ _12041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18148_ rbzero.wall_tracer.visualWallDist\[1\] _11292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18079_ _11200_ _11219_ _11222_ _11223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20110_ _12620_ _12624_ _12882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15875__A1 _08942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21090_ _02051_ _02176_ _02177_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_102_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20041_ _12781_ _12783_ _12778_ _12813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_237_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23800_ _02751_ _04635_ _03889_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_217_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24780_ _05241_ _05232_ _05564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21992_ _03015_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_240_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14850__A2 _08496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23731_ _11193_ _03048_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20943_ _01895_ _02032_ _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_240_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16052__A1 _09522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26450_ _00360_ clknet_leaf_47_i_clk rbzero.debug_overlay.playerX\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23662_ _04459_ _04512_ _04513_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_20874_ _12789_ _01957_ _01826_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__22125__A1 rbzero.wall_tracer.visualWallDist\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25401_ _06184_ _06182_ _06185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22613_ _12163_ _03486_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26381_ _00291_ clknet_leaf_247_i_clk rbzero.spi_registers.buf_texadd2\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14973__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23873__A1 _12499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22676__A2 _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23593_ _03560_ _04445_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25332_ _06053_ _06056_ _06070_ _06116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_22544_ _03435_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13810__C _07604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25263_ _06046_ _06047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_161_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22475_ _03404_ _03406_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_27002_ _00912_ clknet_leaf_193_i_clk rbzero.tex_g0\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24214_ _04946_ _04923_ _04915_ _04934_ _04998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_17_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21426_ _02510_ _02511_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_162_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25194_ _05968_ _05978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24145_ _04915_ _04917_ _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_21357_ rbzero.traced_texVinit\[8\] _01551_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20308_ _12986_ _13005_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21288_ _02205_ _02219_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24076_ _04858_ _04859_ _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_31_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21939__A1 _10048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15309__I _09054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18804__A1 _11449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20239_ _12894_ _12897_ _13010_ _13011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_164_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14213__I _08022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23027_ _03632_ _03883_ _03884_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_164_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15094__A2 _08885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14800_ rbzero.tex_b0\[6\] _08247_ _08607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24353__A2 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15780_ _09402_ _09403_ _09395_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_204_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24978_ _05761_ _05576_ _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22364__A1 _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14841__A2 _07633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14731_ _08534_ _08535_ _08537_ _07463_ _08262_ _08538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_26717_ _00627_ clknet_leaf_29_i_clk rbzero.pov.ready_buffer\[47\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23929_ rbzero.wall_tracer.rcp_fsm.operand\[-8\] _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21962__I1 rbzero.wall_tracer.size\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__26058__B _08909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17450_ rbzero.pov.spi_buffer\[67\] _10742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14662_ rbzero.tex_g1\[52\] _07940_ _08469_ _08470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26648_ _00558_ clknet_leaf_132_i_clk rbzero.tex_b0\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_16401_ rbzero.spi_registers.spi_buffer\[18\] _09865_ _09871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13613_ _06890_ _07423_ _07424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_17381_ rbzero.pov.spi_buffer\[50\] _10685_ _10682_ _10691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__23864__A1 _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18355__I _11478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14593_ rbzero.tex_g1\[31\] _07845_ _08401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26579_ _00489_ clknet_leaf_28_i_clk rbzero.pov.spi_buffer\[48\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_19120_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] _11964_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16332_ _09819_ _09820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13544_ rbzero.row_render.size\[7\] _07355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_94_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_216_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_216_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19051_ _11892_ _11903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_180_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16263_ _08944_ _09759_ _09768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13475_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] _07286_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_153_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18002_ _11145_ rbzero.wall_tracer.trackDistY\[9\] _11146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_152_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15214_ rbzero.spi_registers.spi_buffer\[16\] _08975_ _08982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22605__I _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16194_ _08980_ _09709_ _09716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25369__A1 _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15145_ _08923_ _08925_ _08887_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17846__A2 _10992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19953_ _12723_ _12724_ _12725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__24041__A1 _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15076_ _08868_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13868__B1 _07677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_160_Left_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__19914__I _12685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15219__I _08986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14027_ rbzero.tex_r1\[18\] _07834_ _07836_ _07837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_18904_ _11779_ _11816_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_207_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19884_ _10231_ _12160_ _11097_ _12656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_207_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18835_ _11752_ _11760_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_175_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_223_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18766_ _11713_ _11714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15978_ _09549_ _09552_ _09553_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22355__A1 _11296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14832__A2 _08291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17717_ _10904_ _10629_ _10908_ _10909_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14929_ rbzero.color_sky\[5\] _08735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_19_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20905__A2 _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18697_ rbzero.tex_r1\[19\] rbzero.tex_r1\[18\] _11672_ _11675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_188_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_236_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_236_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17648_ _10858_ _10561_ _10861_ _10863_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_33_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14596__A1 _07507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22658__A2 _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17579_ _10819_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19318_ rbzero.tex_b1\[37\] rbzero.tex_b1\[36\] _12120_ _12121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_20590_ rbzero.wall_tracer.visualWallDist\[6\] _01577_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_18_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14348__A1 _08155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14348__B2 _08156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19249_ _12081_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14899__A2 _07577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22260_ _11238_ _03221_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21211_ _02295_ _02298_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__24407__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22191_ _11284_ _03166_ _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22830__A2 _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21142_ _02226_ _02229_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_76_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_247_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25950_ _06721_ _06730_ _06696_ _06731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__25780__A1 _06051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14033__I _07486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21073_ _02127_ _02161_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_10_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22594__A1 _12231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20024_ _12794_ _12795_ _12796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24901_ _05638_ _05683_ _05685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__16669__B _10113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25881_ _06625_ _06638_ _06643_ _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24335__A2 _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24832_ _05329_ _05492_ _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_214_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24763_ _05499_ _05541_ _05547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21975_ _02991_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer40 _05000_ net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_26502_ _00412_ clknet_leaf_31_i_clk rbzero.debug_overlay.vplaneX\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23714_ _03553_ _04559_ _04560_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_124_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20926_ _12713_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24694_ _05365_ _05470_ _05347_ _05478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_166_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26433_ _00343_ clknet_leaf_213_i_clk rbzero.pov.ss_buffer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23645_ _04403_ _04492_ _04496_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_138_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20857_ _12492_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_194_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26364_ _00274_ clknet_leaf_18_i_clk rbzero.spi_registers.buf_texadd1\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23576_ _04396_ _04428_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20788_ _01877_ _01878_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_25_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25315_ _06097_ _06092_ _06099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22527_ _03439_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26295_ _00205_ clknet_leaf_229_i_clk rbzero.spi_registers.buf_leak\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25246_ _05720_ _06030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_135_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13260_ _07044_ _07074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_22458_ rbzero.wall_tracer.texu\[5\] _03323_ _03299_ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19817__A3 _12282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21409_ _02462_ _02494_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25177_ _05940_ _05960_ _05961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13191_ _07003_ _07004_ _07005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22389_ _12907_ _08049_ _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__20832__A1 _12780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24128_ _04812_ _04718_ _04912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24023__A1 _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14511__A1 _08316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24059_ _04842_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_21_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16950_ _10358_ _10283_ _10363_ _09441_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_124_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15901_ _08822_ _08858_ _09494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19450__A1 _12214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16881_ rbzero.debug_overlay.playerY\[-7\] _08028_ _08048_ rbzero.debug_overlay.playerY\[-6\]
+ _10304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_144_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24326__A2 _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15832_ rbzero.spi_registers.buf_sky\[1\] _09438_ _09442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18620_ rbzero.tex_r0\[50\] rbzero.tex_r0\[49\] _11629_ _11631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_217_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22337__A1 _11282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18551_ _11591_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15763_ rbzero.spi_registers.texadd3\[7\] _09385_ _09391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__26079__A2 _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17502_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _10775_ _10776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14714_ rbzero.tex_b0\[63\] _08288_ _08520_ _08521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_47_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18482_ rbzero.tex_g1\[55\] rbzero.tex_g1\[54\] _11549_ _11552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_234_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18800__I1 rbzero.tex_r1\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15694_ _09305_ _09340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_218_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_177_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17433_ rbzero.pov.spi_buffer\[63\] _10721_ _10729_ _10730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_200_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14645_ _07841_ _08446_ _08452_ _08453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_86_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14578__B2 _07814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17364_ _10676_ _10677_ _10678_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_60_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14576_ rbzero.tex_g1\[21\] _07811_ _08384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_172_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_231_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19103_ _11917_ _11944_ _11946_ _11947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16315_ _09806_ _09807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13527_ _07299_ _07300_ _07338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_17295_ _10602_ _10627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14118__I _07349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24036__B _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19034_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _11893_ _11894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_141_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16246_ rbzero.spi_registers.buf_texadd2\[3\] _09743_ _09755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_235_i_clk clknet_5_1__leaf_i_clk clknet_leaf_235_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_207_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13458_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] _07269_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_149_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16177_ rbzero.spi_registers.buf_texadd1\[10\] _09696_ _09703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17819__A2 rbzero.pov.ready_buffer\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13389_ gpout0.vpos\[4\] _07200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_93_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20823__A1 _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15128_ rbzero.spi_registers.spi_buffer\[0\] _08911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__24550__I _05098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_229_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14502__A1 _08308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19936_ _12338_ _12340_ _12343_ _12223_ _12708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_15059_ _08840_ _08852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22576__A1 _11296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19867_ _11067_ _11983_ _12345_ _12639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14788__I _07603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_201_i_clk_I clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18818_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] _11746_ _11747_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_223_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19798_ _12569_ _12570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_222_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18749_ _11704_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16007__A1 _08946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21760_ _10452_ _02697_ _10455_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20711_ _12705_ _01579_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21691_ _02751_ _02752_ _02753_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23430_ _04171_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20642_ _01711_ _01733_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_19_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13241__A1 _07053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__22500__A1 rbzero.wall_tracer.size\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20573_ _01556_ _01660_ _01664_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_23361_ _04213_ _04215_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_74_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer34_I _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25100_ _05878_ _05883_ _05884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22312_ _03205_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26080_ _06902_ _06846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23292_ _04037_ _04044_ _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14472__B _08280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13867__I _07101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25031_ _05758_ _05805_ _05801_ _05815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_30_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22243_ _11212_ _03206_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22174_ _11981_ _03134_ _03155_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_21125_ _02212_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26982_ _00892_ clknet_leaf_224_i_clk gpout2.clk_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25933_ _06625_ _06638_ _06641_ _06640_ _06710_ _06702_ _06715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_21056_ _02143_ _02144_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20007_ _12688_ _12779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25864_ _06646_ _06647_ _06630_ _06648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_226_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22319__A1 _11163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24815_ _05345_ _05488_ _05599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_241_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25795_ _06559_ _06567_ _06579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_2_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24746_ _05367_ _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_167_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21958_ _02990_ _02984_ _02993_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13480__A1 rbzero.traced_texVinit\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20909_ _12211_ _01859_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24677_ _05239_ _05363_ _05282_ _05461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_90_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21889_ _10113_ _02931_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_210_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15322__I _08877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14430_ _07574_ _08224_ _08238_ _08239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26416_ _00326_ clknet_leaf_18_i_clk rbzero.spi_registers.buf_texadd3\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23628_ _04292_ _02293_ _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_27396_ _01301_ clknet_leaf_76_i_clk rbzero.wall_tracer.stepDistX\[-6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19729__I _12500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_213_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14980__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26347_ _00257_ clknet_leaf_238_i_clk rbzero.spi_registers.buf_texadd0\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14361_ rbzero.debug_overlay.playerX\[0\] _08171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_213_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23559_ _04329_ _04330_ _04411_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 i_mode[2] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16100_ _09595_ _09644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13312_ _07123_ _07035_ _07124_ _07125_ _07052_ _07126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_220_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput29 i_vec_sclk net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17080_ rbzero.pov.ready_buffer\[15\] _10445_ _10465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14292_ rbzero.debug_overlay.vplaneY\[-2\] _08102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_137_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26278_ _00188_ clknet_leaf_245_i_clk rbzero.spi_registers.texadd3\[21\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16031_ _09590_ _09592_ _09587_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_150_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25229_ _06012_ _06013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13535__A2 _07329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14732__A1 _07609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13243_ _07056_ _07057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_123_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24795__A2 _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16153__I _09671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19671__A1 _12439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13174_ _06987_ _06988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_150_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17521__I1 rbzero.tex_b0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15992__I _09428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__19464__I _12235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20281__A2 _12199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_176_Right_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17982_ _11103_ _11104_ _11125_ _11126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_237_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22558__A1 _11291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19721_ _12489_ _12492_ _12493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18226__A2 _11369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16933_ _10346_ _10341_ _10349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16237__A1 _09591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19652_ _12423_ _12424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16864_ _08028_ _08048_ _10289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_244_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18603_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _11618_ _11621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15815_ _09429_ _09430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14799__A1 _08603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19583_ _08041_ _12014_ _12310_ _12354_ _12355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xclkbuf_5_15__f_i_clk clknet_3_3_0_i_clk clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16795_ _10170_ _10228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19026__I1 rbzero.tex_g0\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17712__I _10905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15746_ _09377_ _09378_ _09372_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18534_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _11581_ _11582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_198_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_75_i_clk_I clknet_5_31__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18465_ rbzero.tex_g1\[48\] rbzero.tex_g1\[47\] _11538_ _11542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16328__I _09815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15677_ rbzero.spi_registers.texadd2\[9\] _09326_ _09327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14628_ rbzero.tex_g1\[39\] _07834_ _08436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17416_ rbzero.pov.spi_buffer\[58\] _10717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13223__A1 rbzero.spi_registers.texadd3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18396_ _11503_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__24545__I _05328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17347_ _10665_ _10666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_174_i_clk clknet_5_9__leaf_i_clk clknet_leaf_174_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14559_ _08275_ _08359_ _08367_ _08368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13774__A2 _07584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24235__A1 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23038__A2 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17278_ rbzero.pov.spi_buffer\[23\] _10614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_126_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21049__A1 _12661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13687__I _07482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_16229_ _09457_ _09443_ _09669_ _09741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_19017_ rbzero.tex_g0\[42\] rbzero.tex_g0\[41\] _11882_ _11884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_189_i_clk clknet_5_9__leaf_i_clk clknet_leaf_189_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__19662__A1 _12427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19662__B2 _12433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_228_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_244_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24538__A2 _05321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_244_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_209_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19919_ _12690_ _12691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_112_i_clk clknet_5_31__leaf_i_clk clknet_leaf_112_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_209_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22930_ _03669_ _03786_ _03787_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_208_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22861_ _03712_ _03719_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_24600_ _05360_ _05382_ _05383_ _05384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__15451__A2 _09151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17622__I _10843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21812_ rbzero.debug_overlay.vplaneX\[10\] _11077_ _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_25580_ _06362_ _06363_ _06364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_127_i_clk clknet_5_13__leaf_i_clk clknet_leaf_127_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_104_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22792_ _02071_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22721__A1 _11173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24531_ _05313_ _05314_ _05315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_94_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21743_ _02789_ _02796_ _02797_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16238__I _09711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27250_ _01155_ clknet_leaf_103_i_clk rbzero.wall_tracer.visualWallDist\[-10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24462_ _05086_ _05119_ _05169_ _05246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_171_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21674_ _11132_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26201_ _00111_ clknet_leaf_7_i_clk rbzero.spi_registers.texadd0\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23413_ _04149_ _04166_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20625_ rbzero.wall_tracer.size_full\[6\] _01614_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_27181_ _01086_ clknet_leaf_47_i_clk rbzero.wall_tracer.rayAddendX\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14962__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24393_ _05059_ _05174_ _05176_ _05177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_46_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26132_ _00042_ clknet_leaf_226_i_clk rbzero.pov.sclk_buffer\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23344_ _03845_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20556_ _01647_ _01648_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_172_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26063_ _05007_ _06832_ _06660_ _06833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__25974__A1 _05261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13517__A2 _07327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23275_ _04119_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_20487_ _01579_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25014_ _05792_ _05797_ _05798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22226_ _03196_ _03197_ _03111_ _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19653__A1 _12398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22157_ rbzero.wall_tracer.rcp_fsm.i_data\[-3\] _03126_ _03142_ _03143_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_7_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21108_ _02194_ _02195_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_234_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26965_ _00875_ clknet_leaf_111_i_clk rbzero.texV\[-5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_245_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22088_ _11135_ _07235_ _11136_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_234_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13930_ rbzero.map_overlay.i_mapdx\[1\] _07741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25916_ _06697_ _06623_ _06698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_21039_ _02007_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_35_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26896_ _00806_ clknet_leaf_136_i_clk rbzero.tex_r1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_199_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22960__A1 _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25847_ _06630_ _06631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13861_ _07671_ _07668_ _07672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19169__B1 _12011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15600_ _09258_ _09270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_187_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16580_ rbzero.wall_tracer.rayAddendY\[2\] _10030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_215_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25778_ _06530_ _06562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13792_ _07331_ _07603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15531_ _09205_ _09218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24729_ _05361_ _05265_ _05513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18250_ _11393_ _11394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_91_i_clk clknet_5_26__leaf_i_clk clknet_leaf_91_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_155_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27448_ _01353_ clknet_leaf_72_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_15462_ _09167_ _09168_ _09162_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17201_ rbzero.pov.spi_buffer\[4\] _10556_ _10552_ _10557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19459__I _12202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14413_ _07935_ _08222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13756__A2 _07566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18181_ rbzero.map_overlay.i_othery\[1\] _11302_ _11325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_27379_ _01284_ clknet_leaf_105_i_clk rbzero.wall_tracer.trackDistY\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15393_ _09117_ _09118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_245_Right_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17132_ rbzero.pov.ready_buffer\[6\] _10489_ _10504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14344_ _08151_ _08006_ _08010_ _08152_ _08022_ _08153_ _08154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_108_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19892__A1 _12211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17063_ _10447_ _10450_ _10451_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14275_ rbzero.debug_overlay.facingX\[-6\] _08085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21938__B _09934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25196__I _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16014_ _08957_ _09574_ _09580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13226_ _07039_ _07040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23440__A2 _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13157_ rbzero.texu_hot\[2\] _06955_ _06970_ _06971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_226_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_185_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13088_ _06902_ _06903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17965_ rbzero.map_rom.f1 _11109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_29_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19704_ _12475_ _12476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21203__A1 _11296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16916_ _07713_ _10328_ _10334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17896_ rbzero.debug_overlay.facingX\[10\] _11033_ _11040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_44_i_clk clknet_5_16__leaf_i_clk clknet_leaf_44_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_192_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19635_ _12320_ _12322_ _10208_ _12324_ _12407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_16847_ _10181_ _10274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_204_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_204_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19566_ _12337_ _12338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_189_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13444__A1 _07139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16778_ _09855_ _10214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_177_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18517_ _11572_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_158_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15729_ rbzero.spi_registers.texadd2\[22\] _09362_ _09366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16058__I _09428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19497_ _12176_ _11991_ _12246_ _12268_ _12269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xclkbuf_leaf_59_i_clk clknet_5_23__leaf_i_clk clknet_leaf_59_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_201_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24275__I _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20190__A1 _12841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18448_ _11532_ _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_1_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13747__A2 _07537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18379_ _11493_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_248_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20410_ _12561_ _12297_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_212_Right_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__24208__A1 _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21390_ _02472_ _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_161_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24208__B2 _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20341_ _01435_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18150__A4 _11293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21690__A1 _10359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23060_ _03793_ _03796_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20272_ _01366_ _13034_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22523__I _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22011_ rbzero.wall_tracer.rcp_fsm.o_data\[10\] rbzero.wall_tracer.size_full\[10\]
+ _02985_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__20245__A2 _12011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25708__A1 _06037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Left_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_228_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24392__B1 _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26750_ _00660_ clknet_leaf_121_i_clk rbzero.wall_tracer.mapX\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23962_ rbzero.wall_tracer.rcp_fsm.i_data\[-2\] _04755_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_243_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17949__A1 _08076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25701_ _06448_ _06458_ _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input24_I i_tex_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22913_ _03708_ _03742_ _03770_ _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14976__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26681_ _00591_ clknet_leaf_26_i_clk rbzero.pov.ready_buffer\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23893_ _04708_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_155_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25632_ _06350_ _06356_ _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_169_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22844_ _03701_ _03702_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25563_ _05521_ _06024_ _05967_ _06347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_151_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22775_ _02644_ _02678_ _02676_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_156_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27302_ _01207_ clknet_leaf_201_i_clk rbzero.row_render.texu\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24514_ _05297_ _05298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_137_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21726_ _02768_ _02781_ _02783_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25494_ _06153_ _06155_ _06278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24447__A1 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27233_ _01138_ clknet_leaf_86_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24445_ _05228_ _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21657_ _02692_ _08491_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15600__I _09258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14644__C _07924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20608_ _12206_ _01433_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_163_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27164_ _01069_ clknet_leaf_209_i_clk rbzero.map_rom.i_col\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24376_ _04978_ _05107_ _05108_ _05109_ _05160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_21588_ _02672_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26115_ _00025_ clknet_leaf_241_i_clk rbzero.spi_registers.spi_buffer\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18141__A4 _11284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23327_ _01744_ _04062_ _04058_ _04064_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_160_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20539_ _12431_ _12968_ _01377_ _01631_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_27095_ _01005_ clknet_leaf_141_i_clk rbzero.tex_b1\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_34_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_23_i_clk_I clknet_5_20__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26046_ _06634_ _06644_ _06818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14060_ rbzero.tex_r1\[4\] _07829_ _07870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23258_ _04019_ _04113_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_162_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14163__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14660__B _07946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22209_ _03177_ _03184_ _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23189_ _04037_ _04044_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_167_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_233_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14962_ net6 _08759_ _08764_ _08765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_17750_ _10928_ rbzero.pov.ready_buffer\[40\] _10931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26948_ _00858_ clknet_leaf_180_i_clk rbzero.tex_r1\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_50_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21736__A2 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16701_ _10067_ _10140_ _10143_ _10144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_221_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_248_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13913_ rbzero.map_overlay.i_otherx\[0\] _07078_ _07724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_221_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14893_ rbzero.tex_b1\[43\] _07484_ _08699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_17681_ _10882_ rbzero.pov.ready_buffer\[16\] _10886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26879_ _00789_ clknet_leaf_161_i_clk rbzero.tex_r0\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13790__I _07448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17262__I _10542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19420_ _12191_ _12192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16632_ _10057_ _10060_ _10079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_18_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13844_ _07651_ _07652_ _07653_ _07654_ _07541_ _07655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_186_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19351_ _12139_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16563_ _09917_ _10015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13775_ _07442_ _07586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18302_ rbzero.hsync _11440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_168_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15514_ _09204_ _09205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16494_ _09949_ _09950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_19282_ _12100_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_210_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15445_ rbzero.spi_registers.vshift\[2\] _09151_ _09156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14926__A1 _08360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18233_ _11330_ _11368_ _11376_ _11377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_66_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18117__A1 rbzero.debug_overlay.playerX\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23110__A1 _12212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15376_ _09102_ _09104_ _09100_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18164_ _11255_ _11308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__19865__A1 _12283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17115_ _10488_ _10490_ _10492_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14327_ _08125_ _08011_ _08017_ _08126_ _08136_ _08137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_18095_ _11197_ _11238_ _11204_ _11202_ _11222_ _11239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_187_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17046_ _10427_ _10437_ _10438_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__19617__A1 _12384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14258_ _07720_ _07202_ _08067_ _08068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__24461__I1 _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21424__A1 _12666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13209_ rbzero.spi_registers.texadd0\[21\] _07020_ _07022_ _07023_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14189_ _06872_ _07189_ _07999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_241_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25166__A2 _05948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_30__f_i_clk clknet_3_7_0_i_clk clknet_5_30__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_18997_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _11872_ _11873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_225_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_206_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15654__A2 _09303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24913__A2 _05696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17948_ rbzero.wall_tracer.rayAddendX\[10\] _11092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_240_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14796__I _07337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17879_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] _11023_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_19618_ _12389_ _12390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_178_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20890_ _11388_ _01979_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_85_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19549_ _11041_ _11067_ _11068_ _11085_ _12321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_88_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_215_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_165_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16717__S _10125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22560_ _11290_ _03455_ _03456_ rbzero.traced_texa\[3\] _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21511_ _02595_ _02078_ _01969_ _12414_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22491_ _03416_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15420__I _09029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24230_ _05012_ _05013_ _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_151_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21442_ _02526_ _02527_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_151_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24161_ _04888_ _04944_ _04945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_116_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21373_ _02397_ _02434_ _02458_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_226_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23112_ _03844_ _01945_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20324_ _01415_ _01418_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24092_ _04869_ _04863_ _04831_ _04876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA_clkbuf_leaf_197_i_clk_I clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Left_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17347__I _10665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23043_ _03771_ _03774_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20255_ _13015_ _13026_ _13027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__16251__I _09747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20186_ _12957_ _12958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26802_ _00712_ clknet_leaf_168_i_clk rbzero.tex_g1\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24994_ _05420_ _05332_ _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_99_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23945_ rbzero.wall_tracer.rcp_fsm.operand\[-5\] _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_99_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26733_ _00643_ clknet_leaf_42_i_clk rbzero.pov.ready_buffer\[63\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26664_ _00574_ clknet_leaf_153_i_clk rbzero.tex_b0\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_233_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23876_ _04689_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_169_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25615_ _06344_ _06397_ _06398_ _06399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_169_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22827_ _02277_ _02120_ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13959__A2 _07212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26595_ _00505_ clknet_leaf_42_i_clk rbzero.pov.spi_buffer\[64\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_25546_ _06327_ _06329_ _06330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13560_ _07365_ _07059_ _07056_ _07367_ _07369_ _07370_ _07371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XANTENNA__20154__A1 _12668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22758_ _11409_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14908__A1 _08304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21709_ _11331_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25477_ _06250_ _06254_ _06261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_26_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13491_ _07293_ _07294_ _07302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_82_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22689_ _11199_ rbzero.wall_tracer.stepDistX\[-7\] _03551_ _03557_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_180_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15230_ _08993_ _08995_ _08988_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_27216_ _01121_ clknet_leaf_75_i_clk rbzero.wall_tracer.stepDistY\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24428_ _05118_ _05212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__19847__A1 _12476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27147_ _00003_ clknet_leaf_73_i_clk rbzero.wall_tracer.rcp_fsm.state\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15161_ rbzero.spi_registers.spi_buffer\[6\] _08939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24359_ _05141_ _05142_ _05085_ _05143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14112_ rbzero.tex_r1\[44\] _07919_ _07921_ _07922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_73_Left_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15092_ _08883_ _08884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_27078_ _00988_ clknet_leaf_153_i_clk rbzero.tex_b1\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_132_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26029_ _06626_ _06621_ _06732_ _06733_ _06710_ _06645_ _06803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_18920_ _10757_ _11828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14043_ _07841_ _07852_ _07853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_197_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17086__A1 _08143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_223_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18851_ _11769_ _11773_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23159__A1 _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19472__I _11382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17802_ _10958_ _10717_ _10961_ _10964_ _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_100_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18782_ rbzero.tex_r1\[56\] rbzero.tex_r1\[55\] _11719_ _11723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15994_ _09561_ _09563_ _09565_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_235_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17733_ _10912_ _10645_ _10916_ _10919_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14945_ net4 _08748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_82_Left_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14549__C _08357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17664_ _10843_ _10874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_201_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14876_ rbzero.tex_b1\[32\] _08496_ _08682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19403_ rbzero.wall_tracer.side _12175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16615_ _10062_ _10063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13827_ _07449_ _07638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_134_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17595_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _10828_ _10829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_197_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19334_ _12129_ _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16546_ _09923_ _09998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13758_ _07560_ _07568_ _07569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19265_ _12090_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16477_ _09916_ _09934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13689_ rbzero.tex_r0\[55\] _07499_ _07500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_234_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18216_ _11301_ _11360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15428_ rbzero.color_floor\[4\] _09129_ _09143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19196_ _11130_ _11378_ _12040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Left_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_208_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21645__A1 _09942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18147_ rbzero.wall_tracer.visualWallDist\[2\] _11291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15359_ _09077_ _09092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14127__A2 _07641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18078_ _11220_ _11221_ _11195_ _11196_ _11222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_145_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17029_ rbzero.pov.ready_buffer\[25\] _10425_ _10426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20040_ _12667_ _12807_ _12808_ _12809_ _12811_ _12812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21991_ rbzero.wall_tracer.rcp_fsm.o_data\[3\] rbzero.wall_tracer.size_full\[3\]
+ _02985_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_23730_ _11221_ _04554_ _04574_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20942_ _02030_ _02031_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16955__B _10214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23661_ _04459_ _04512_ _02732_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_20873_ _01824_ _01825_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_89_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18329__A1 _10988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25400_ _06025_ _06184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22125__A2 _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22612_ _03490_ _03495_ _03496_ _03193_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_159_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26380_ _00290_ clknet_leaf_1_i_clk rbzero.spi_registers.buf_texadd2\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23592_ _04358_ _04441_ _04444_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__23873__A2 _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__17001__A1 _08079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25331_ _06108_ _06114_ _06115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_193_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22543_ _03448_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__23788__B _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25262_ _06045_ _06046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22474_ _10256_ _11449_ _03405_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_173_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_27001_ _00911_ clknet_leaf_193_i_clk rbzero.tex_g0\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24213_ _04852_ _04872_ _04880_ _04891_ _04997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_16_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21425_ _12689_ _02112_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25193_ _05948_ _05977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24144_ _04919_ _04927_ _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__15315__A1 _07736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21356_ _02309_ _02442_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_32_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20307_ _13009_ _01400_ _01401_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_24075_ _04764_ _04856_ _04857_ _04859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_21287_ _02206_ _02218_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13877__A1 _07687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_229_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23026_ _03633_ _03749_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_20238_ _12895_ _12896_ _13010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_164_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20611__A2 _12496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20169_ _12608_ _12671_ _12941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_216_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_129_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__24353__A3 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24977_ _05561_ _05565_ _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_231_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15325__I _09034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22364__A2 _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14730_ rbzero.tex_b0\[44\] _08298_ _08536_ _08537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26716_ _00626_ clknet_leaf_29_i_clk rbzero.pov.ready_buffer\[46\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_203_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23928_ _04731_ _04732_ _10508_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14661_ rbzero.tex_g1\[53\] _07625_ _08469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_23859_ _12395_ _04687_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26647_ _00557_ clknet_leaf_132_i_clk rbzero.tex_b0\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_200_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14054__A1 rbzero.tex_r1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24361__I0 _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16400_ rbzero.spi_registers.buf_texadd3\[18\] _09863_ _09870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13612_ gpout0.hpos\[7\] _07423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_14592_ rbzero.tex_g1\[30\] _07843_ _08400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17380_ rbzero.pov.spi_buffer\[49\] _10690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_26578_ _00488_ clknet_leaf_27_i_clk rbzero.pov.spi_buffer\[47\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16331_ _09818_ _09819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13543_ rbzero.row_render.size\[8\] _07354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25529_ _06270_ _06306_ _06312_ _06313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_45_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_216_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_216_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16262_ rbzero.spi_registers.buf_texadd2\[7\] _09757_ _09767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19050_ _11902_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13474_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] _07285_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_125_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_18001_ rbzero.wall_tracer.trackDistX\[9\] _11145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15213_ _08979_ _08981_ _08971_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16193_ rbzero.spi_registers.buf_texadd1\[14\] _09707_ _09715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15144_ _08924_ _08907_ _08925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25369__A2 _06012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_26__f_i_clk_I clknet_3_6_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19952_ _12674_ _12430_ _12681_ _12724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_26_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15075_ _08822_ _08863_ _08865_ _08867_ _08868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__24041__A2 _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13868__A1 _07244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13868__B2 _07678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14026_ rbzero.tex_r1\[19\] _07835_ _07836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_18903_ rbzero.traced_texa\[8\] _07262_ _11815_ _11816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_19883_ _12615_ _12651_ _12654_ _12655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__17715__I _10884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18834_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] _11759_ _11760_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_101_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_223_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18765_ _11649_ _11713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15977_ _09504_ _09553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17716_ _10906_ rbzero.pov.ready_buffer\[28\] _10909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_171_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14928_ _07801_ _08728_ _08731_ _08733_ _08734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_18696_ _11674_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_145_i_clk_I clknet_5_14__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17647_ _10859_ rbzero.pov.ready_buffer\[5\] _10863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_236_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_202_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_195_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14859_ rbzero.tex_b1\[0\] _08248_ _08665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23304__A1 _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17578_ rbzero.tex_b0\[46\] rbzero.tex_b0\[45\] _10817_ _10819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_147_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19317_ _12114_ _12120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_128_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16529_ _09934_ _09982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14348__A2 _08040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15545__A1 rbzero.spi_registers.buf_texadd1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19248_ rbzero.tex_b1\[7\] rbzero.tex_b1\[6\] _12078_ _12081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24804__A1 _05388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19179_ _12019_ _12021_ _12022_ _12023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_182_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21210_ _02296_ _02297_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22190_ _03154_ _03169_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__24407__I1 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21141_ _02227_ _02228_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_223_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_247_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14520__A2 _08317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21072_ _02131_ _02160_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_238_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22594__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20023_ _12707_ _12710_ _12795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24900_ _05637_ _05638_ _05683_ _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_25880_ _06645_ _06663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_225_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24831_ _05419_ _05252_ _05303_ _05286_ _05615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_225_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24762_ _05491_ _05496_ _05546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_21974_ rbzero.wall_tracer.rcp_fsm.o_data\[-3\] _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xrebuffer30 _05138_ net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_179_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer41 net92 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__23362__I _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23713_ _04527_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26501_ _00411_ clknet_leaf_56_i_clk rbzero.debug_overlay.facingY\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_124_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20925_ _01806_ _02014_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_124_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24693_ _05476_ _05372_ _05477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_139_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23644_ _04493_ _04494_ _04495_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_26432_ _00342_ clknet_leaf_229_i_clk rbzero.pov.ss_buffer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20856_ _12733_ _01945_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14587__A2 _08317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24394__S _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23846__A2 _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26363_ _00273_ clknet_leaf_7_i_clk rbzero.spi_registers.buf_texadd1\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23575_ _04399_ _04427_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20787_ _12489_ _12956_ _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25314_ _06097_ _06092_ _06098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__25289__I _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22526_ _12834_ _03436_ _03438_ rbzero.traced_texa\[-11\] _03439_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_187_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25599__A2 _06382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26294_ _00204_ clknet_leaf_229_i_clk rbzero.spi_registers.buf_leak\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21609__A1 _11456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25245_ _06002_ _06019_ _06028_ _06029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_150_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22457_ _03396_ _03397_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_157_Right_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__24271__A2 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14652__C _07935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_21408_ _02478_ _02493_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25176_ _05933_ _05934_ _05947_ _05959_ _05960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13190_ rbzero.spi_registers.texadd3\[18\] _06997_ _06992_ rbzero.spi_registers.texadd2\[18\]
+ _06998_ rbzero.spi_registers.texadd1\[18\] _07004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_22388_ _12947_ _01363_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_115_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24127_ _04905_ _04907_ _04910_ _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_21339_ _12382_ _01466_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20832__A2 _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25220__A1 _06003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24058_ _04841_ rbzero.wall_tracer.rcp_fsm.operand\[8\] _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23009_ _03865_ _03866_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15900_ _09492_ _09493_ _09491_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_159_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16880_ rbzero.debug_overlay.playerY\[-6\] rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerY\[-8\]
+ rbzero.debug_overlay.playerY\[-9\] _10303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__23909__I0 rbzero.wall_tracer.rcp_fsm.o_data\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15831_ _08911_ _09439_ _09440_ _09441_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_217_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13078__A2 _06888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22597__B _12229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18550_ rbzero.tex_r0\[20\] rbzero.tex_r0\[19\] _11587_ _11591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20348__A1 _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15762_ _09389_ _09390_ _09384_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_231_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17501_ _10759_ _10775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_231_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14713_ rbzero.tex_b0\[62\] _08291_ _08520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_47_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18481_ _11551_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__18366__I _11480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15693_ rbzero.spi_registers.texadd2\[13\] _09338_ _09339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_218_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_177_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_218_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17432_ _10705_ _10729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14644_ _08447_ _08449_ _08451_ _07923_ _07924_ _08452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__13731__C _07541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23837__A2 _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21848__B2 _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14575_ rbzero.tex_g1\[23\] _07807_ _07808_ _08383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17363_ rbzero.pov.spi_buffer\[45\] _10674_ _10671_ _10678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20115__A4 _12501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19102_ _11945_ _11946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16314_ _09659_ _09806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_231_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13526_ _07336_ _07337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_125_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17294_ rbzero.pov.spi_buffer\[27\] _10626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_137_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19033_ _11892_ _11893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_179_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16245_ _09753_ _09754_ _09750_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13457_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] _07268_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_125_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_179_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22273__A1 rbzero.wall_tracer.visualWallDist\[-5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13388_ gpout0.vpos\[5\] _07199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16176_ _09701_ _09702_ _09700_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_93_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_71_i_clk_I clknet_5_29__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15127_ _08903_ _08907_ _08910_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20823__A2 _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19935_ _12705_ _12706_ _12707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_15058_ _08832_ _08851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_229_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_208_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14009_ _07524_ _07819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22576__A2 _09974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19866_ _12636_ _12637_ _12638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__19441__A2 _12212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18817_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] _11745_ _11746_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__25514__A2 _06102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19797_ _12568_ _12569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_223_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18748_ rbzero.tex_r1\[41\] rbzero.tex_r1\[40\] _11703_ _11704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__24278__I _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18679_ _11664_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14018__B2 _07826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20710_ _01799_ _01800_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_21690_ _10359_ _02740_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20641_ _01714_ _01732_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13213__I _06927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23360_ _03861_ _04214_ _04056_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_191_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20572_ _01557_ _01659_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18180__A2 rbzero.map_rom.f2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22311_ _03268_ _03269_ _03252_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23291_ _04144_ _04071_ _04145_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16191__A1 _08977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25030_ _05634_ _05812_ _05813_ _05814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_5_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22242_ _03202_ _03208_ _03212_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14741__A2 _08206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22173_ _11292_ _03135_ _03083_ _12908_ _03114_ _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_169_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21124_ _12231_ _02210_ _02211_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_26981_ _00891_ clknet_leaf_224_i_clk gpout2.clk_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_25932_ _06700_ _06709_ _06713_ _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_21055_ _02013_ _02022_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20006_ _12777_ _12686_ _12778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25863_ _06373_ _06422_ _06647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__14257__A1 _08062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14257__B2 _08066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24814_ _05545_ _05597_ _05598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_25794_ _06560_ _06566_ _06577_ _06578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_2_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13832__B _07642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21957_ rbzero.wall_tracer.size_full\[-9\] _02992_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24745_ _05473_ _05474_ _05527_ _05528_ _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_29_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13480__A2 rbzero.spi_registers.vshift\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_226_Right_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20908_ _01865_ _01866_ _01997_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24676_ _05397_ _05458_ _05459_ _05460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_21888_ _02925_ _02926_ _02929_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_194_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26415_ _00325_ clknet_leaf_19_i_clk rbzero.spi_registers.buf_texadd3\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23627_ _03979_ _04180_ _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20839_ _01921_ _01928_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_27395_ _01300_ clknet_leaf_106_i_clk rbzero.wall_tracer.stepDistX\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_42_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14360_ _08019_ _08070_ _08169_ _08170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_213_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23558_ _04321_ _04327_ _04331_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_26346_ _00256_ clknet_leaf_11_i_clk rbzero.spi_registers.buf_texadd0\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15759__B _09384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_213_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13311_ rbzero.spi_registers.texadd3\[2\] _07027_ _07028_ _07125_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 i_reg_csb net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_22509_ _03427_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14291_ _08099_ _08036_ _08047_ _08100_ _08101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_26277_ _00187_ clknet_leaf_1_i_clk rbzero.spi_registers.texadd3\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23489_ _04234_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_165_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16030_ _09591_ _09585_ _09592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13242_ gpout0.hpos\[1\] _07056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_162_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25228_ _05824_ _05865_ _06011_ _06012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_33_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__27175__CLK clknet_5_17__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25159_ _05872_ _05907_ _05943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_32_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13173_ _06930_ _06984_ _06986_ _06987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_150_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22007__A1 _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25744__A2 _06440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17981_ _11105_ _11124_ _11125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14496__A1 rbzero.tex_g0\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13793__I _07603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19720_ _12491_ _12492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23755__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16932_ _10346_ _10341_ _10348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_229_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19651_ _12422_ _12423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_53_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16863_ _10182_ _10288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_205_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19480__I _12165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18602_ _11620_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15814_ _09428_ _09429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19582_ _11953_ _11999_ _10305_ _12004_ _12354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__15996__A1 _08983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16794_ _07709_ _10215_ _10227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22120__B _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18533_ _11565_ _11581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15745_ rbzero.spi_registers.buf_texadd3\[2\] _09375_ _09378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_18_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15513__I _08876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18464_ _11541_ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15676_ _09302_ _09326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17415_ _10715_ _10713_ _10716_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_201_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14627_ _08431_ _08432_ _08433_ _08434_ _07924_ _08435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_185_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18395_ rbzero.tex_g1\[17\] rbzero.tex_g1\[16\] _11502_ _11503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22494__A1 rbzero.wall_tracer.size\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17346_ _10546_ _10665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14558_ _08363_ _08366_ _07670_ _08367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13509_ _07260_ _07319_ gpout0.vinf _07320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_17277_ _10610_ _10606_ _10613_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_181_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14489_ _08276_ _08298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19016_ _11883_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21049__A2 _12594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16228_ _09739_ _09740_ _09734_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14723__A2 _08529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19111__A1 _08159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19655__I _12426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16159_ rbzero.spi_registers.buf_texadd1\[5\] _09685_ _09690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19662__A2 _12428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_244_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14487__B2 _08294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19918_ _12501_ _12690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_209_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19414__A2 _12185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_209_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17108__C _10357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19849_ _12409_ _12500_ _12621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25499__A1 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19390__I _12159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22860_ _03715_ _03718_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14748__B _08459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24171__A1 _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21811_ rbzero.debug_overlay.vplaneX\[10\] _11077_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_88_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22791_ _02593_ _02597_ _02594_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__16519__I _09972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15423__I _06898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24530_ _05218_ net63 _05314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_21742_ _11103_ _02782_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24736__I _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24461_ _05152_ _05220_ _05082_ _05245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21673_ _02737_ _12021_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23412_ _04167_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_26200_ _00110_ clknet_leaf_239_i_clk rbzero.spi_registers.texadd0\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20624_ rbzero.wall_tracer.size_full\[6\] _01614_ _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27180_ _01085_ clknet_leaf_47_i_clk rbzero.wall_tracer.rayAddendX\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24392_ _05042_ _05062_ _05063_ _05064_ _05175_ _05176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_190_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26131_ _00041_ clknet_leaf_250_i_clk rbzero.spi_registers.spi_buffer\[23\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23343_ _12950_ _03792_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20555_ _12659_ _12448_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16254__I _09761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23796__B _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26062_ _06780_ _06806_ _06831_ _06803_ _06771_ _06691_ _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_119_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23274_ _04124_ _04125_ _04128_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__14714__A2 _08288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20486_ _01578_ _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_225_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25013_ _05793_ _05796_ _05797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__24404__C _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22225_ _12163_ _11394_ _03080_ _03091_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_104_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19653__A2 _12403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22156_ _11988_ _03134_ _03141_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14478__A1 rbzero.tex_g0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21107_ _02188_ _02193_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26964_ _00874_ clknet_leaf_111_i_clk rbzero.texV\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_22087_ _11129_ _12163_ _07239_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__21748__B1 _09921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25915_ _06650_ _06697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_21038_ _02057_ _02126_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_227_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26895_ _00805_ clknet_leaf_136_i_clk rbzero.tex_r1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_199_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25846_ _05047_ _06630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13860_ rbzero.color_sky\[0\] _07671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_234_i_clk clknet_5_3__leaf_i_clk clknet_leaf_234_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25777_ _06519_ _06525_ _06561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22989_ _03845_ _02524_ _03716_ _03718_ _02336_ _03846_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_4
X_13791_ rbzero.tex_r0\[4\] _07600_ _07601_ _07602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15333__I _09054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13453__A2 rbzero.spi_registers.vshift\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18767__I1 rbzero.tex_r1\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15530_ _09215_ _09216_ _09217_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24728_ _05292_ _05410_ _05512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_195_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27447_ _01352_ clknet_leaf_71_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_139_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15461_ rbzero.spi_registers.buf_texadd0\[0\] _09165_ _09168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24659_ _05240_ _05258_ _05265_ _05273_ _05443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_155_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_249_i_clk clknet_5_0__leaf_i_clk clknet_leaf_249_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_231_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17200_ _10555_ _10556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_166_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14412_ rbzero.tex_g0\[25\] _08210_ _08220_ _08221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18180_ rbzero.map_overlay.i_otherx\[2\] rbzero.map_rom.f2 _11324_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__22476__A1 _07153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27378_ _01283_ clknet_leaf_104_i_clk rbzero.wall_tracer.trackDistY\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15392_ _08882_ _09117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_93_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17131_ _08118_ _10487_ _10503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14343_ rbzero.debug_overlay.facingY\[-3\] _08153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_26329_ _00239_ clknet_leaf_234_i_clk rbzero.spi_registers.buf_mapdxw\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19892__A2 _12224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26565__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_244_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14274_ rbzero.debug_overlay.facingX\[-8\] _08084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17062_ rbzero.pov.ready_buffer\[11\] _10445_ _10451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14705__A2 _08252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16013_ rbzero.spi_registers.buf_mapdy\[4\] _09572_ _09579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13225_ gpout0.hpos\[0\] _07039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_90_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19644__A2 _11998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13156_ _06957_ _06969_ _06970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_226_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23728__A1 _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13087_ _06901_ _06902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17964_ _11106_ _11100_ _11108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19703_ _11385_ _12366_ _12474_ _12475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__21203__A2 _12229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16915_ _07704_ _10328_ _10333_ _10221_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_224_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17895_ _11035_ _11038_ _11039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__17723__I _10905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19634_ rbzero.wall_tracer.visualWallDist\[-4\] _11381_ _11383_ _12406_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_205_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16846_ _10166_ _10269_ _10264_ _10273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24153__A1 _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_204_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19565_ _08042_ _12014_ _12310_ _12336_ _12337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_137_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16777_ _08176_ _10212_ _10213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_220_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13989_ _07764_ _07789_ _07798_ _07799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_232_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23900__A1 _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18516_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _11571_ _11572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15728_ _09363_ _09365_ _09361_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19496_ _12175_ _11076_ _12268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18447_ rbzero.tex_g1\[40\] rbzero.tex_g1\[39\] _11528_ _11532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15659_ _09289_ _09314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_200_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18378_ rbzero.tex_g1\[10\] rbzero.tex_g1\[9\] _11491_ _11493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_145_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17329_ rbzero.pov.spi_buffer\[36\] _10652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__16074__I _09614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24208__A2 _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_20340_ _12399_ _01433_ _01434_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13904__B1 _07052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20271_ _12952_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22010_ _03026_ _02986_ _03027_ _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_102_Left_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_209_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__24392__B2 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23961_ _04757_ _04758_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18729__I _11692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25700_ _06477_ _06483_ _06484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__18997__I1 rbzero.tex_g0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22912_ _03706_ _03743_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23892_ rbzero.wall_tracer.rcp_fsm.o_data\[2\] rbzero.wall_tracer.stepDistX\[2\]
+ _04685_ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_26680_ _00590_ clknet_leaf_23_i_clk rbzero.pov.ready_buffer\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24144__A1 _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25850__I _05212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I i_mode[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25631_ _06395_ _06396_ _06414_ _06415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_22843_ _03643_ _03700_ _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16249__I _09742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15153__I _08932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_193_i_clk_I clknet_5_12__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25562_ _05237_ _05605_ _05967_ _06346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_177_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22774_ _02580_ _02683_ _02681_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27301_ _01206_ clknet_leaf_201_i_clk rbzero.row_render.size\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24513_ _05296_ _05297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21725_ _11343_ _02782_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25493_ _06271_ _06276_ _06277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_23_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_111_Left_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27232_ _01137_ clknet_leaf_86_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22458__A1 rbzero.wall_tracer.texu\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24444_ _05083_ _05220_ _05221_ _05222_ _05227_ _05005_ _05228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
X_21656_ _02725_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_192_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18126__A2 _11269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20607_ rbzero.wall_tracer.stepDistX\[3\] _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_24375_ _05065_ _05067_ _05069_ _04959_ _05159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__16137__A1 rbzero.spi_registers.buf_texadd1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27163_ _01068_ clknet_leaf_202_i_clk rbzero.map_rom.f1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_21587_ _02666_ _02671_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_151_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26114_ _00024_ clknet_leaf_241_i_clk rbzero.spi_registers.spi_buffer\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23326_ _04179_ _04180_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20538_ _01468_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27094_ _01004_ clknet_leaf_141_i_clk rbzero.tex_b1\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_26045_ _06802_ _03010_ _06814_ _06817_ _06810_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_23257_ _04025_ _04112_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20469_ _01465_ _01490_ _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22208_ _11281_ _03096_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21433__A2 _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23188_ _03918_ _04043_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_37_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22139_ _11991_ _03121_ _03094_ _03127_ _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_167_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13123__B2 rbzero.spi_registers.texadd2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14961_ net6 _08763_ _08764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26947_ _00857_ clknet_leaf_181_i_clk rbzero.tex_r1\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__13674__A2 _07484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14871__A1 _08315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16700_ _10122_ _10141_ _10142_ _10115_ _10143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xclkbuf_leaf_173_i_clk clknet_5_9__leaf_i_clk clknet_leaf_173_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_50_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13912_ _07720_ _07721_ _07722_ _07678_ _07723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_221_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17680_ _10884_ _10885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_180_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14892_ _07535_ _08698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26878_ _00788_ clknet_leaf_161_i_clk rbzero.tex_r0\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_57_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16631_ _10074_ _10077_ _10078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13292__B _07045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25829_ _06611_ _06601_ _06606_ _06612_ _06613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_13843_ rbzero.tex_r0\[16\] _07420_ _07586_ _07654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_214_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19350_ rbzero.tex_b1\[51\] rbzero.tex_b1\[50\] _12136_ _12139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16562_ _10009_ _10010_ _10013_ _10014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_58_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13774_ rbzero.tex_r0\[1\] _07584_ _07585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_188_i_clk clknet_5_3__leaf_i_clk clknet_leaf_188_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__19562__A1 rbzero.wall_tracer.stepDistX\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18301_ _11431_ _11439_ _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15513_ _08876_ _09204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19281_ rbzero.tex_b1\[21\] rbzero.tex_b1\[20\] _12099_ _12100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_167_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16493_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] _09931_
+ _09949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24438__A2 _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18232_ _11299_ _11370_ _11371_ _11375_ _11376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_128_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15444_ _09152_ _09155_ _09149_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18117__A2 rbzero.map_rom.f4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_i_clk clknet_5_31__leaf_i_clk clknet_leaf_111_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18163_ _11250_ _11307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__21121__A1 _12194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15375_ rbzero.spi_registers.buf_leak\[2\] _09103_ _09104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17114_ _10491_ _10492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14326_ _08130_ _08135_ _08136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25938__A2 _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18094_ rbzero.wall_tracer.trackDistX\[-7\] _11238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_123_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_187_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17045_ rbzero.pov.ready_buffer\[29\] _10425_ _10438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14257_ _08062_ _08064_ _08065_ _08066_ _08067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_126_i_clk clknet_5_13__leaf_i_clk clknet_leaf_126_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13362__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13362__B2 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13208_ _07020_ _07021_ _07022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__18676__I0 rbzero.tex_r1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14188_ _07997_ _07998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_241_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13139_ _06909_ _06953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18996_ _11871_ _11872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_206_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13114__A1 _06927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_206_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I i_gpout1_sel[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18428__I0 rbzero.tex_g1\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17947_ _11040_ _11089_ _11090_ _11091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_206_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17878_ _11007_ _11019_ _11021_ _11022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_19617_ _12384_ _12388_ _12389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_16829_ _07687_ _10258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_68_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19548_ _12319_ _12320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__14090__A2 _07857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19479_ _12248_ _11990_ _12180_ _12250_ _12251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__16367__A1 _08955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21510_ _02068_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14378__B1 _08036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14917__A2 _08554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22490_ rbzero.wall_tracer.size\[3\] _03410_ _03412_ _07372_ _03416_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_185_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21441_ _02410_ _02413_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24160_ _04737_ _04906_ _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_116_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22534__I _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21372_ _02331_ _02396_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__25929__A2 _06652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23111_ _03851_ _01957_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20323_ _01416_ _01417_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_24091_ _04768_ _04805_ _04875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_142_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_229_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25845__I _06628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23042_ _03882_ _03885_ _03888_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_20254_ _12303_ _13025_ _13026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20989__I _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20185_ _12956_ _12957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_228_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_90_i_clk clknet_5_24__leaf_i_clk clknet_leaf_90_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24365__A1 _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26801_ _00711_ clknet_leaf_175_i_clk rbzero.tex_g1\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_244_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_24993_ _05505_ _05506_ _05775_ _05776_ _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_243_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14853__B2 _08502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26732_ _00642_ clknet_leaf_42_i_clk rbzero.pov.ready_buffer\[62\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23944_ _04744_ _04745_ _04736_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_162_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26663_ _00573_ clknet_leaf_153_i_clk rbzero.tex_b0\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_223_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23875_ _02997_ _04690_ _04698_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_212_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25614_ _06338_ _06342_ _06398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22826_ _02001_ _02502_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26594_ _00504_ clknet_leaf_33_i_clk rbzero.pov.spi_buffer\[63\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14081__A2 _07890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25545_ _06274_ _06275_ _06276_ _06328_ _06329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__16358__A1 _08944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20154__A2 _12728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22757_ _03547_ _03616_ _03617_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14369__B1 _08017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13490_ _07299_ _07300_ _07301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21708_ _02767_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25476_ _06257_ _06259_ _06260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_165_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22688_ _02760_ _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_212_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27215_ _01120_ clknet_leaf_109_i_clk rbzero.wall_tracer.stepDistY\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_165_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24427_ _05035_ _05091_ _05210_ _05211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21639_ _09944_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27146_ _00002_ clknet_leaf_72_i_clk rbzero.wall_tracer.rcp_fsm.state\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__17858__A1 rbzero.debug_overlay.facingX\[-2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15160_ _08936_ _08938_ _08934_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24358_ _05133_ net62 _05054_ _05142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__22851__A1 _12760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_43_i_clk clknet_5_16__leaf_i_clk clknet_leaf_43_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_117_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_16__f_i_clk_I clknet_3_4_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14111_ rbzero.tex_r1\[45\] _07920_ _07921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23309_ _04155_ _04163_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15091_ _08882_ _08883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_239_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24289_ _05059_ _05061_ _05072_ _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_27077_ _00987_ clknet_leaf_153_i_clk rbzero.tex_b1\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__16442__I _09899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13344__A1 _07153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26028_ _06902_ _06802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14042_ _07589_ _07847_ _07851_ _07852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_120_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_i_clk clknet_5_23__leaf_i_clk clknet_leaf_58_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_18850_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] _11772_ _11773_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_120_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_223_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24356__A1 _05133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17801_ _10959_ rbzero.pov.ready_buffer\[58\] _10964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_206_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18781_ _11722_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_206_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15993_ _09564_ _09565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17732_ _10913_ rbzero.pov.ready_buffer\[34\] _10919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_206_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14944_ net82 _08747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__24371__A4 _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19783__A1 _12402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17663_ _10872_ _10873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_187_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14875_ rbzero.tex_b1\[34\] _08250_ _08308_ _08681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_201_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19402_ rbzero.wall_tracer.size_full\[-11\] _12173_ _12174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_201_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16614_ rbzero.wall_tracer.rayAddendY\[4\] _10062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_187_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13826_ rbzero.tex_r0\[24\] _07635_ _07636_ _07637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_207_Left_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17594_ _10822_ _10828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_203_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_197_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19535__A1 _12305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14072__A2 _07876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_197_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19333_ rbzero.tex_b1\[44\] rbzero.tex_b1\[43\] _12125_ _12129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_202_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16545_ _09924_ _09996_ _09997_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13757_ _07562_ _07564_ _07565_ _07567_ _07551_ _07568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__20145__A2 _12915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19264_ rbzero.tex_b1\[14\] rbzero.tex_b1\[13\] _12088_ _12090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16476_ _08099_ _09933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_183_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13688_ _07498_ _07499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_14_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15021__A1 _08807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_234_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18215_ _11342_ _11346_ _11351_ _11358_ _11359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__19928__I _12352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23095__A1 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15427_ _09140_ _09141_ _09142_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_19195_ _11329_ _11368_ _11376_ _12038_ _12039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_183_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24831__A2 _05252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18146_ rbzero.wall_tracer.visualWallDist\[3\] _11290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_171_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15358_ rbzero.mapdyw\[0\] _09090_ _09091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23890__I0 rbzero.wall_tracer.rcp_fsm.o_data\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14309_ _08116_ _08007_ _08023_ _08118_ _08119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_clkbuf_leaf_141_i_clk_I clknet_5_14__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_216_Left_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18077_ _11193_ _11221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_41_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15289_ rbzero.map_overlay.i_othery\[1\] _09019_ _09040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17028_ _10396_ _10425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15088__A1 _07164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16824__A2 _10183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18979_ _11862_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__17183__I _10541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21990_ _03014_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__19774__A1 _12504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23913__I _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20941_ _01897_ _01898_ _02029_ _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_225_Left_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__16588__A1 _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20872_ _01837_ _01846_ _01835_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_23660_ _04463_ _04467_ _04511_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_152_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18329__A2 _07202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14063__A2 _07835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_66_i_clk_I clknet_5_21__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22611_ _11135_ _03489_ _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23591_ _04253_ _04442_ _04443_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22542_ rbzero.wall_tracer.visualWallDist\[-4\] _03443_ _03444_ rbzero.traced_texa\[-4\]
+ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_25330_ _06109_ _06113_ _06114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_48_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21884__A2 _08143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25075__A2 _05856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25261_ _05822_ _05756_ _06044_ _06045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__14047__I _07518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22473_ _07160_ _08750_ _11443_ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_146_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24822__A2 _05605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27000_ _00910_ clknet_leaf_193_i_clk rbzero.tex_g0\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24212_ _04914_ _04928_ _04938_ _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_21424_ _12666_ _02233_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25192_ _05333_ _05975_ _05976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__22833__A1 _12691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21636__A2 _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_234_Left_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_161_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24143_ _04920_ _04921_ _04901_ _04926_ _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_86_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21355_ _02312_ _02441_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20306_ _01399_ _13027_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24074_ _04856_ _04857_ _04764_ _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21286_ _02371_ _02372_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19573__I rbzero.wall_tracer.side vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23025_ _03633_ _03749_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_20237_ _13007_ _12920_ _13008_ _13009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_164_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15079__A1 _07719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_164_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20168_ _12870_ _12939_ _12940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_157_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19065__I0 rbzero.tex_g0\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_243_Left_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20099_ _12615_ _12651_ _12871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24976_ _05554_ _05594_ _05759_ _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_98_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26715_ _00625_ clknet_leaf_29_i_clk rbzero.pov.ready_buffer\[45\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_243_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23927_ rbzero.wall_tracer.rcp_fsm.i_data\[-9\] _04728_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14660_ rbzero.tex_g1\[55\] _07938_ _07946_ _08468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26646_ _00556_ clknet_leaf_132_i_clk rbzero.tex_b0\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23858_ _04683_ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14054__A2 _07818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24510__A1 _05292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13611_ _07420_ _07421_ _07332_ _07422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_22809_ _02491_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_184_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14591_ _07848_ _08397_ _08398_ _08399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_26577_ _00487_ clknet_leaf_27_i_clk rbzero.pov.spi_buffer\[46\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23789_ _11184_ _04619_ _04626_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13801__A2 _07584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16330_ _08829_ _09745_ _09818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_55_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25528_ _06307_ _06311_ _06312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_223_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13542_ rbzero.row_render.size\[9\] _07353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_165_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21875__A2 _11069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15003__A1 _06900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_216_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16261_ _09765_ _09766_ _09762_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25459_ _06234_ _06228_ _06243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_216_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15554__A2 _09232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14357__A3 _08166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13473_ _07282_ _07283_ _07284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18000_ _11139_ rbzero.wall_tracer.trackDistX\[10\] _11141_ _11143_ _11144_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_164_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15212_ _08980_ _08969_ _08981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16192_ _09713_ _09714_ _09712_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15143_ rbzero.spi_registers.spi_buffer\[2\] _08924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16172__I _09660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27129_ _01039_ clknet_leaf_120_i_clk rbzero.traced_texVinit\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19951_ _12721_ _12722_ _12435_ _12723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_15074_ rbzero.spi_registers.sclk_buffer\[1\] _08866_ _08867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13868__A2 _07676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14025_ _07531_ _07835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18902_ _11811_ _11813_ _11814_ _11815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_19882_ _12567_ _12600_ _12653_ _12654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__20063__A1 _12834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18833_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] _11758_ _11759_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18764_ _11712_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15976_ _08965_ _09551_ _09552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_207_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_199_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19756__A1 _12527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17715_ _10884_ _10908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14927_ _07475_ _08732_ _07665_ _08733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18695_ rbzero.tex_r1\[18\] rbzero.tex_r1\[17\] _11672_ _11674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_216_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17646_ _10858_ _10558_ _10861_ _10862_ _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_26_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14858_ _08660_ _08661_ _08663_ _08294_ _08509_ _08664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_236_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13809_ rbzero.tex_r0\[12\] _07600_ _07587_ _07620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20118__A2 _12500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16347__I _09819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17577_ _10818_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_175_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14789_ rbzero.tex_b0\[3\] _07930_ _08596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19316_ _12119_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16528_ _09970_ _09976_ _09981_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19247_ _12080_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16459_ _09916_ _09917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_155_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19178_ rbzero.map_rom.b6 _12015_ _12022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_170_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_6__f_i_clk clknet_3_1_0_i_clk clknet_5_6__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_18129_ _11270_ _11271_ _11272_ _11273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_131_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_21140_ _01484_ _01924_ _01925_ _12779_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25860__S0 _06628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21071_ _02132_ _02159_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_67_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19995__A1 _12761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20022_ _12786_ _12792_ _12793_ _12794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23791__A2 rbzero.wall_tracer.stepDistY\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_207_Right_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24830_ _05337_ _05613_ _05607_ _05614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__17470__A2 _10547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24739__I _05522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24761_ _05343_ _05543_ _05544_ _05545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_21973_ _03003_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_213_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer20 _05508_ net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer31 _04846_ net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_26500_ _00410_ clknet_leaf_55_i_clk rbzero.debug_overlay.facingY\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__17641__I _10844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23712_ _04530_ _04558_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xrebuffer42 _05269_ net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_20924_ _01802_ _01808_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_124_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24692_ _05356_ _05476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_124_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15233__A1 _08997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14036__A2 _07845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26431_ _00341_ clknet_leaf_243_i_clk rbzero.spi_registers.spi_cmd\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20855_ _01944_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23643_ _04219_ _04052_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16981__A1 _08085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26362_ _00272_ clknet_leaf_7_i_clk rbzero.spi_registers.buf_texadd1\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24474__I _05257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20786_ _01875_ _01876_ _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_23574_ _04426_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18183__B1 _11255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19568__I _12339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25313_ _06026_ _06095_ _06096_ _06097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_22525_ _03437_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_148_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26293_ _00203_ clknet_leaf_233_i_clk rbzero.spi_registers.buf_leak\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25244_ _06021_ _06023_ _06027_ _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_22456_ _07713_ _07709_ _03342_ _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21407_ _02480_ _02492_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_40_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25175_ _05888_ _05957_ _05958_ _05959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22387_ _01453_ _03332_ _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24126_ _04909_ _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_21338_ _12299_ _01631_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22722__I _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24057_ rbzero.wall_tracer.rcp_fsm.operand\[7\] _04830_ _04834_ _04831_ _04841_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_21269_ _02335_ _02355_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23782__A2 rbzero.wall_tracer.stepDistY\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23008_ _03684_ _03687_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_159_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_217_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15336__I _09074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23909__I1 rbzero.wall_tracer.stepDistX\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15830_ _09113_ _09441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__24326__A4 _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13284__C _07074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15761_ rbzero.spi_registers.buf_texadd3\[6\] _09387_ _09390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24959_ _05737_ _05740_ _05741_ _05742_ _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_17500_ _10774_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14712_ rbzero.tex_b0\[60\] _08518_ _08289_ _08519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18480_ rbzero.tex_g1\[54\] rbzero.tex_g1\[53\] _11549_ _11551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_47_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15692_ _09302_ _09338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15224__A1 _08990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14027__A2 _07834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_218_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_177_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_218_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17431_ rbzero.pov.spi_buffer\[62\] _10728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_197_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14643_ rbzero.tex_g1\[44\] _08291_ _08450_ _08451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26629_ _00539_ clknet_leaf_160_i_clk rbzero.tex_b0\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_185_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16972__A1 _08084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14822__I1 _08628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17362_ _10665_ _10677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_185_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21848__A2 _10040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14574_ rbzero.tex_g1\[22\] _07805_ _08382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_200_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19101_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] _11945_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16313_ _09005_ _09804_ _09805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13525_ _07335_ _07336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_231_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17293_ _10623_ _10619_ _10625_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_165_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19032_ _11828_ _11892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16244_ _08915_ _09748_ _09754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13456_ rbzero.texV\[7\] _07267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22273__A2 _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16175_ _08955_ _09698_ _09702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19674__B1 _12419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13387_ _07196_ _07197_ _07198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__20284__A1 _12427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_149_Left_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_14_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15126_ rbzero.spi_registers.spi_buffer\[0\] _08906_ _08909_ _08910_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17726__I _09034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19934_ _12487_ _12706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23222__A1 _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15057_ _08847_ _08848_ _08849_ _08850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_229_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20036__A1 _12433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14008_ _07518_ _07818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19865_ _12283_ _12521_ _12637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19941__I _12261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18816_ _11744_ _11745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_128_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19796_ _12490_ _12568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_208_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_235_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19162__B _12005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18747_ _11692_ _11703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15959_ _09537_ _09538_ _09536_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_239_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18678_ rbzero.tex_r1\[11\] rbzero.tex_r1\[10\] _11661_ _11664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_106_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17629_ _08809_ _10850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20640_ _01724_ _01731_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19388__I _12159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18292__I _10271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20571_ _01663_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_184_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16715__A1 _10145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22310_ _11292_ _03250_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23290_ _04033_ _04046_ _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22241_ _12834_ _03210_ _03211_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22172_ _10151_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__17140__A1 _10145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21123_ rbzero.wall_tracer.stepDistX\[10\] _12231_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_140_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26980_ _00890_ clknet_leaf_124_i_clk rbzero.texV\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_245_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25931_ _06711_ _06712_ _06699_ _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20062__I rbzero.wall_tracer.visualWallDist\[-11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21054_ _02015_ _02021_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_245_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21775__A1 _10121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20005_ _12691_ _12777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_126_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25862_ _06424_ _06467_ _06646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_226_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14257__A2 _08064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24813_ _05596_ _05546_ _05597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_119_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25793_ _06561_ _06565_ _06577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18467__I _11479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24744_ _05365_ _05470_ _05476_ _05528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_21956_ _02991_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_201_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_190_Right_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_179_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15206__A1 rbzero.spi_registers.spi_buffer\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20907_ _01996_ _01642_ _01863_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_96_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24675_ _05328_ _05399_ _05459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_166_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16954__A1 rbzero.pov.ready_buffer\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21887_ _02925_ _02926_ _02929_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_26414_ _00324_ clknet_leaf_19_i_clk rbzero.spi_registers.buf_texadd3\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23626_ _04385_ _04388_ _04477_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_27394_ _01299_ clknet_leaf_79_i_clk rbzero.wall_tracer.stepDistX\[-8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_193_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20838_ _01922_ _01927_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_166_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19298__I _12093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26345_ _00255_ clknet_leaf_11_i_clk rbzero.spi_registers.buf_texadd0\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23557_ _04323_ _04333_ _04409_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_213_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20769_ _12236_ _01859_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_213_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13310_ rbzero.spi_registers.texadd2\[2\] _07108_ _07109_ rbzero.spi_registers.texadd1\[2\]
+ _07124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14663__C _07464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22508_ rbzero.wall_tracer.size\[10\] _03423_ _03424_ rbzero.row_render.size\[10\]
+ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_190_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14290_ rbzero.debug_overlay.vplaneY\[-9\] _08100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26276_ _00186_ clknet_leaf_0_i_clk rbzero.spi_registers.texadd3\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_220_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23488_ _04253_ _04255_ _04341_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_80_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25227_ _05867_ _05807_ _06011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13241_ _07053_ _07054_ _07055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22439_ _03380_ _03381_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_220_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13279__C _07057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25158_ _05912_ _05941_ _05942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13172_ rbzero.spi_registers.texadd1\[14\] _06985_ _06981_ rbzero.spi_registers.texadd0\[14\]
+ _06929_ _06986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_20_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_188_i_clk_I clknet_5_3__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17131__A1 _08118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_229_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24109_ _04862_ _04873_ _04892_ _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_TAPCELL_ROW_150_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23204__A1 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17980_ _11107_ _11104_ _11123_ _11124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25089_ _05773_ _05832_ _05791_ _05835_ _05873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_130_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15693__A1 rbzero.spi_registers.texadd2\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14496__A2 _07600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16931_ _10346_ _10329_ _10347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19423__A3 _12015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21766__A1 _08143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19650_ _12421_ _12422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16862_ _10283_ _10285_ _10287_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_53_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15445__A1 rbzero.spi_registers.vshift\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18601_ rbzero.tex_r0\[42\] rbzero.tex_r0\[41\] _11618_ _11620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15813_ _08931_ _09428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19581_ _12338_ _12340_ _12343_ _12352_ _12353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_clkbuf_leaf_240_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16793_ _10222_ _10215_ _10226_ _10221_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_18532_ _11580_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15744_ rbzero.spi_registers.texadd3\[2\] _09373_ _09377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22191__A1 _11284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18463_ rbzero.tex_g1\[47\] rbzero.tex_g1\[46\] _11538_ _11541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15675_ _09323_ _09324_ _09325_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_185_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15748__A2 _09375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17414_ rbzero.pov.spi_buffer\[58\] _10709_ _10706_ _10716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14626_ rbzero.tex_g1\[32\] _07894_ _07630_ _08434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18394_ _11501_ _11502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_114_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14420__A2 _07832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17345_ rbzero.pov.spi_buffer\[40\] _10664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14557_ _07665_ _08365_ _08366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13508_ rbzero.traced_texVinit\[10\] rbzero.texV\[10\] _07318_ _07319_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_17276_ rbzero.pov.spi_buffer\[23\] _10603_ _10612_ _10613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14488_ rbzero.tex_g0\[45\] _08210_ _08297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_24__f_i_clk clknet_3_6_0_i_clk clknet_5_24__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_157_Left_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19015_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _11882_ _11883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16227_ _09667_ _09732_ _09740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13439_ _07249_ _06859_ net1 _07250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_180_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_248_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16158_ _09686_ _09688_ _09689_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__17122__A1 _08106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19872__S _12159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15109_ rbzero.spi_registers.spi_counter\[3\] _08857_ _08892_ _08897_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__16360__I _09815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16089_ _09614_ _09637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__20009__A1 _12780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_244_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15684__A1 rbzero.spi_registers.texadd2\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19917_ _12688_ _12689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_48_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_209_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_209_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19848_ _12558_ _12618_ _12619_ _12620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_108_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_166_Left_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__25499__A2 _06012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21706__I _11397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13933__B _07743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19779_ _12549_ _12550_ _12551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__19178__A2 _12015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21810_ _10121_ _02857_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_22790_ _03647_ _03648_ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_121_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21741_ _08175_ _02784_ _02795_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16936__A1 _10345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24460_ _05005_ _05141_ _05243_ _05133_ _05244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_21672_ _12035_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_176_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23411_ _04190_ _04231_ _04264_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20623_ _01524_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_149_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24391_ _04865_ _05066_ _05068_ _05070_ _05175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_190_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_175_Left_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26130_ _00040_ clknet_leaf_249_i_clk rbzero.spi_registers.spi_buffer\[22\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23342_ _04196_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_20554_ _12930_ _12690_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26061_ _06830_ _06698_ _06629_ _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23273_ _04126_ _04127_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20485_ rbzero.wall_tracer.visualWallDist\[5\] _01577_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_15_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25012_ _05794_ _05795_ _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22224_ _11391_ _02091_ _03084_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_42_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19653__A3 _12414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_22155_ _11288_ _03135_ _03130_ _11071_ _03136_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_100_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14478__A2 _08258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21106_ _02188_ _02193_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26963_ _00873_ clknet_leaf_111_i_clk rbzero.texV\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_22086_ _08379_ _08374_ _07775_ _07236_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_7_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_184_Left_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_227_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25914_ _05076_ _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21037_ _02106_ _02125_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_201_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26894_ _00804_ clknet_leaf_176_i_clk rbzero.tex_r0\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_35_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22221__B _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25845_ _06628_ _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_226_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13843__B _07586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25776_ _06531_ _06534_ _06560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13790_ _07448_ _07601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22988_ _12212_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22173__A1 _11292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22173__B2 _12908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14650__A2 _07906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24727_ _05445_ _05448_ _05510_ _05511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_195_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21939_ _10048_ _02976_ _02977_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16927__A1 rbzero.pov.ready_buffer\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27446_ _01351_ clknet_leaf_71_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15460_ rbzero.spi_registers.texadd0\[0\] _09163_ _09167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24658_ _05240_ _05266_ _05273_ _05258_ _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_193_Left_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14411_ _07825_ _08220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23609_ _04330_ _04460_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27377_ _01282_ clknet_leaf_105_i_clk rbzero.wall_tracer.trackDistY\[-3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15391_ rbzero.color_sky\[0\] _09115_ _09116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24589_ _05352_ _05372_ _05373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_25_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17130_ _06900_ _10501_ _10502_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14342_ rbzero.debug_overlay.facingY\[-2\] _08152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_26328_ _00238_ clknet_leaf_233_i_clk rbzero.spi_registers.buf_mapdxw\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17061_ _10449_ _10443_ _10450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22228__A2 _11377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14273_ _08081_ _08045_ _08047_ _08082_ _08083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_26259_ _00169_ clknet_leaf_241_i_clk rbzero.spi_registers.texadd3\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16012_ _09577_ _09578_ _09576_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13224_ _07026_ _07037_ _07038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13913__A1 rbzero.map_overlay.i_otherx\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25178__A1 _05912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13155_ rbzero.texu_hot\[1\] _06961_ _06968_ _06969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_55_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_226_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13086_ rbzero.wall_tracer.rcp_fsm.state\[1\] _06901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17963_ _11106_ _11107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19702_ rbzero.wall_tracer.stepDistX\[-9\] _12288_ _12474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13141__A2 _06952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16914_ rbzero.pov.ready_buffer\[51\] _10201_ _10329_ _10332_ _10333_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_205_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17894_ _11036_ _11037_ _11038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19633_ rbzero.debug_overlay.playerY\[-4\] _12013_ _12254_ _12404_ _12405_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_192_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16845_ _10271_ _10272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_205_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25350__A1 _05948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_204_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19564_ _11954_ _11999_ _10297_ _12004_ _12336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_16776_ _10178_ _10212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_204_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22164__A1 _11286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13988_ _07686_ _07791_ _07792_ _07797_ _07798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_125_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14641__A2 _08448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15727_ rbzero.spi_registers.buf_texadd2\[21\] _09364_ _09365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18515_ _11565_ _11571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_19495_ _11383_ _12267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_5_5__f_i_clk_I clknet_3_1_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19580__A2 _12202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18446_ _11531_ _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15658_ rbzero.spi_registers.buf_texadd2\[4\] _09306_ _09313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14609_ rbzero.tex_g1\[6\] _07579_ _07580_ _08417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_83_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18377_ _11492_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15589_ rbzero.spi_registers.buf_texadd1\[10\] _09259_ _09262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17328_ _10648_ _10641_ _10651_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18391__I0 rbzero.tex_g1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17259_ rbzero.pov.spi_buffer\[19\] _10591_ _10599_ _10600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13904__A1 _07709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20270_ _12947_ _01363_ _01364_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__13904__B2 _07699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17186__I _10544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15657__A1 rbzero.spi_registers.texadd2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23719__A2 _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24392__A2 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23960_ _04721_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__20402__A1 _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14880__A2 _08494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22911_ _03638_ _03748_ _03746_ _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__23852__S _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23891_ _04707_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_223_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25630_ _06399_ _06411_ _06413_ _06414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__24144__A2 _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22842_ _03643_ _03700_ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__22155__A1 _11288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_136_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22155__B2 _11071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25561_ _06338_ _06342_ _06344_ _06345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_196_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22773_ _02577_ _02579_ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_151_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27300_ _01205_ clknet_leaf_209_i_clk rbzero.row_render.size\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24512_ _05295_ _05296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_156_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21724_ _11399_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25492_ _06143_ _06272_ _06273_ _06274_ _06275_ _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_176_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13889__I _07699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27231_ _01136_ clknet_leaf_86_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14396__A1 _07463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24443_ _04719_ _05223_ _05224_ _05226_ _05227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_21655_ _02724_ _08377_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__16265__I _09742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20606_ _01692_ _01697_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_152_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27162_ _01067_ clknet_leaf_208_i_clk rbzero.map_rom.f2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24374_ _05040_ _05043_ _04967_ _05158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21586_ _02667_ _02670_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_105_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26113_ _00023_ clknet_leaf_241_i_clk rbzero.spi_registers.spi_buffer\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14148__A1 _07928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23325_ _01920_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23407__A1 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16688__A3 _10024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20537_ _01473_ _01475_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_144_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27093_ _01003_ clknet_leaf_140_i_clk rbzero.tex_b1\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_144_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26044_ _06768_ _06815_ _06741_ _06816_ _06742_ _06817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_23256_ _04110_ _04111_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20468_ _01462_ _01559_ _01560_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__21969__A1 rbzero.wall_tracer.size\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22207_ _03163_ _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_247_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_23187_ _03922_ _04038_ _04042_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20399_ _01402_ _01442_ _01492_ _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_218_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22138_ rbzero.wall_tracer.visualWallDist\[-6\] _03100_ _03117_ _11076_ _03127_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_167_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14320__A1 _08128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14960_ _08761_ _08762_ _08763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26946_ _00856_ clknet_leaf_178_i_clk rbzero.tex_r1\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_22069_ _03017_ _03060_ _03068_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_199_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14871__A2 _08676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13911_ rbzero.map_overlay.i_otherx\[1\] _07722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26877_ _00787_ clknet_leaf_164_i_clk rbzero.tex_r0\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14891_ rbzero.tex_b1\[41\] _07592_ _08214_ _08697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_221_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_221_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16073__A1 _08957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16630_ _10075_ _10076_ _10077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25828_ _06602_ _06605_ _06612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13842_ rbzero.tex_r0\[17\] _07583_ _07653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15820__A1 rbzero.spi_registers.texadd3\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14623__A2 _07890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16561_ _09993_ _10011_ _10012_ _10013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_25759_ _06538_ _06539_ _06542_ _06543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_13773_ _07583_ _07584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18655__I _11650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22697__A2 rbzero.wall_tracer.stepDistX\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18300_ _11432_ _07228_ _11436_ _11438_ rbzero.vga_sync.vsync _11439_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_15512_ _06907_ _09180_ _09203_ _09182_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_57_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19280_ _12093_ _12099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16492_ rbzero.wall_tracer.rayAddendY\[-3\] _09948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18231_ _11372_ _11374_ _11375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27429_ _01334_ clknet_leaf_69_i_clk rbzero.wall_tracer.rcp_fsm.operand\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15443_ rbzero.spi_registers.buf_vshift\[1\] _09154_ _09155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_210_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18162_ _11256_ _11306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_15374_ _09077_ _09103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_17113_ _08932_ _10491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14325_ _08132_ _08063_ _08059_ _08134_ gpout0.vpos\[3\] _08135_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_18093_ _11144_ _11236_ _11237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17044_ _08152_ _10423_ _10437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14256_ rbzero.debug_overlay.playerY\[5\] _08066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_187_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13207_ rbzero.spi_registers.texadd3\[21\] _07014_ _07009_ rbzero.spi_registers.texadd2\[21\]
+ _07015_ rbzero.spi_registers.texadd1\[21\] _07021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_111_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14187_ _07983_ _07996_ _07997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__18676__I1 rbzero.tex_r1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13138_ rbzero.spi_registers.texadd3\[8\] _06920_ _06923_ rbzero.spi_registers.texadd2\[8\]
+ _06915_ rbzero.spi_registers.texadd1\[8\] _06952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_241_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18995_ _11828_ _11871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_209_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_206_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17946_ rbzero.debug_overlay.facingX\[10\] _11033_ _11090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13069_ gpout0.hpos\[3\] _06885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_224_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22385__A1 _12907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14862__A2 _08528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_206_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17877_ _08087_ _11020_ _11021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19616_ _12385_ _12387_ _12388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16828_ _10254_ _10257_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_233_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14614__A2 _07843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19547_ _11091_ _11038_ _12319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_76_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16759_ _10195_ _10196_ _10197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_75_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19478_ _12249_ _11074_ _12250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_186_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14378__A1 _07699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18429_ _11521_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14378__B2 _08180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23637__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25398__I _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21440_ _02411_ _02412_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_134_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18364__I0 rbzero.tex_g1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19856__A3 _12496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21371_ _02453_ _02456_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_116_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20322_ _12490_ _12584_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23110_ _12212_ _03842_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_233_i_clk clknet_5_3__leaf_i_clk clknet_leaf_233_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24090_ _04772_ _04808_ _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20253_ _13024_ _13025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23041_ _12035_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_62_i_clk_I clknet_5_21__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20184_ rbzero.wall_tracer.visualWallDist\[2\] _12200_ _12956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_86_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_248_i_clk clknet_5_0__leaf_i_clk clknet_leaf_248_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_26800_ _00710_ clknet_leaf_170_i_clk rbzero.tex_g1\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__24365__A2 _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13105__A2 _06918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24992_ _05563_ _05564_ _05776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__22376__A1 _11394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25861__I _06628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26731_ _00641_ clknet_leaf_32_i_clk rbzero.pov.ready_buffer\[61\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23943_ rbzero.wall_tracer.rcp_fsm.i_data\[-6\] _04740_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15164__I _08935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_162_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26662_ _00572_ clknet_leaf_154_i_clk rbzero.tex_b0\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__24477__I _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23874_ rbzero.wall_tracer.stepDistX\[-6\] _04694_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14605__A2 _07811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25613_ _06338_ _06342_ _06397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_169_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22825_ _02540_ _01580_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26593_ _00503_ clknet_leaf_33_i_clk rbzero.pov.spi_buffer\[62\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25544_ _06271_ _06328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22756_ _11168_ _03605_ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14369__A1 _07701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21707_ _02766_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_165_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25475_ _06136_ _06258_ _06139_ _06259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__14508__I _07831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22687_ _03547_ _03554_ _03555_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_27214_ _01119_ clknet_leaf_108_i_clk rbzero.wall_tracer.stepDistY\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24426_ _05136_ _05090_ _05210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21638_ _09915_ _02703_ rbzero.wall_tracer.rayAddendY\[-9\] _02714_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22300__A1 _11286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27145_ _00001_ clknet_leaf_73_i_clk rbzero.wall_tracer.rcp_fsm.state\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24357_ net92 _05132_ _05134_ net71 _05140_ _05141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_151_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21569_ _02650_ _02653_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_151_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14110_ _07582_ _07920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15869__A1 _09462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23308_ _04156_ _04161_ _04162_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_169_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24053__A1 _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27076_ _00986_ clknet_leaf_152_i_clk rbzero.tex_b1\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_15090_ _08881_ _08882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24288_ _05040_ _05062_ _05063_ _05064_ _05071_ _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__24940__I _05640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26027_ _06800_ _06801_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_132_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14041_ _07848_ _07849_ _07850_ _07851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_23239_ _03984_ _03987_ _04094_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_132_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23800__A1 _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__27175__D _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_223_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17800_ _10958_ _10715_ _10961_ _10963_ _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_235_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18780_ rbzero.tex_r1\[55\] rbzero.tex_r1\[54\] _11719_ _11722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15992_ _09428_ _09564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_147_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22367__A1 rbzero.mapdyw\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14844__A2 _07595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17731_ _10912_ _10643_ _10916_ _10918_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_14943_ rbzero.hsync _08744_ _08746_ net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_26929_ _00839_ clknet_leaf_172_i_clk rbzero.tex_r1\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__16046__A1 _09515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__26088__B _06842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19783__A2 _12553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14874_ rbzero.tex_b1\[35\] _08298_ _08680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17662_ _10847_ _10872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__26519__D _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19401_ _12172_ _12173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_201_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16613_ _10056_ _10058_ _10060_ _10061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_13825_ _07524_ _07636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_230_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17593_ _10827_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_197_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15802__I _09117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16544_ _09992_ _09940_ _09997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19332_ _12128_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13756_ rbzero.tex_r0\[44\] _07566_ _07549_ _07567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_156_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__23619__A1 _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16475_ _09928_ rbzero.wall_tracer.rayAddendY\[-4\] _09931_ _09932_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_39_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19263_ _12089_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_63_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13687_ _07482_ _07498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14418__I _08226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_234_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15426_ rbzero.spi_registers.buf_floor\[3\] _08885_ _09142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18214_ _11305_ _11356_ _11357_ _11358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_234_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19194_ _11299_ _11314_ _12038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_170_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18145_ _11286_ _11287_ _11288_ _11289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_15357_ _09074_ _09090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_171_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23890__I1 rbzero.wall_tracer.stepDistX\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_130_Left_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_170_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14308_ _08117_ _08118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18076_ rbzero.wall_tracer.trackDistX\[-5\] _11220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_145_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15288_ _07721_ _09031_ _09039_ _09036_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_180_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17027_ _08155_ _10423_ _10424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_229_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24595__A2 _05264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14239_ _08048_ _08049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13992__I _07326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15088__A2 _08879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18978_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _11861_ _11862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14835__A2 _08248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17929_ _08088_ _11072_ _11022_ _11073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_206_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21030__A1 _12705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20940_ _01897_ _01898_ _02029_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20871_ _01935_ _01943_ _01960_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__18295__I _07979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15260__A2 _08885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22610_ _03493_ _03471_ _03480_ _03482_ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_23590_ _04255_ _04341_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_220_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22530__A1 rbzero.wall_tracer.visualWallDist\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22541_ _03447_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14328__I rbzero.debug_overlay.vplaneX\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13232__I _07045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25260_ _05635_ _05755_ _06044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22545__I _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22472_ _08750_ _11443_ _07160_ _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24211_ _04977_ _04987_ _04993_ _04994_ _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_0_106_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21423_ _12777_ _01917_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25191_ _05974_ _05975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_172_i_clk clknet_5_9__leaf_i_clk clknet_leaf_172_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__22833__A2 _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24142_ _04922_ _04886_ _04923_ _04925_ _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__20065__I _12836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21354_ _02314_ _02440_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_20_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19854__I _12486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20305_ _01399_ _13027_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14523__A1 _08245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24073_ _04811_ _04761_ _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21285_ _02230_ _02238_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23024_ _03768_ _03769_ _03881_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xclkbuf_leaf_187_i_clk clknet_5_9__leaf_i_clk clknet_leaf_187_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_20236_ _12904_ _12905_ _13008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__19462__A1 _10224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20167_ _12873_ _12925_ _12938_ _12939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_129_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14826__A2 _08631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_110_i_clk clknet_5_31__leaf_i_clk clknet_leaf_110_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_20098_ _12670_ _12868_ _12869_ _12870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24975_ _05557_ _05593_ _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_232_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23926_ _04730_ _04725_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26714_ _00624_ clknet_leaf_29_i_clk rbzero.pov.ready_buffer\[44\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13851__B _07570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26645_ _00555_ clknet_leaf_146_i_clk rbzero.tex_b0\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23857_ _04685_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__23849__A1 rbzero.wall_tracer.stepDistY\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13610_ _07336_ _07421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22808_ _02608_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_125_i_clk clknet_5_13__leaf_i_clk clknet_leaf_125_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13262__A1 _07046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14590_ rbzero.tex_g1\[28\] _08226_ _08398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26576_ _00486_ clknet_leaf_27_i_clk rbzero.pov.spi_buffer\[45\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23788_ _03624_ _04624_ _04625_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__24935__I _05308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21324__A2 _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25527_ _05996_ _05975_ _06308_ _06310_ _06144_ _06311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_13541_ _07346_ _07350_ _07351_ _07352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22739_ _03600_ _03594_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16200__A1 rbzero.spi_registers.buf_texadd1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16260_ _08939_ _09759_ _09766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_216_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25458_ _06240_ _06241_ _06242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13472_ rbzero.texV\[6\] _07274_ _07283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_192_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_192_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15211_ rbzero.spi_registers.spi_buffer\[14\] _08980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18154__B _11295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24409_ _05075_ _05138_ _05139_ _05193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_63_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14762__A1 rbzero.tex_b0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16191_ _08977_ _09709_ _09714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25389_ _06072_ _06093_ _06173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15142_ _08922_ _08918_ _08923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27128_ _01038_ clknet_leaf_120_i_clk rbzero.traced_texVinit\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16503__A2 rbzero.wall_tracer.rayAddendY\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19950_ _12432_ _12429_ _12722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_22_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15073_ rbzero.spi_registers.sclk_buffer\[2\] _08866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_27059_ _00969_ clknet_leaf_133_i_clk rbzero.tex_b1\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__22588__A1 rbzero.wall_tracer.wall\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14024_ _07594_ _07834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_18901_ rbzero.traced_texa\[7\] _07267_ _11814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19881_ _12652_ _12599_ _12653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_120_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20063__A2 _12301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18832_ _11755_ _11757_ _11758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_18763_ rbzero.tex_r1\[48\] rbzero.tex_r1\[47\] _11708_ _11712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_234_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15975_ _09550_ _09551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_223_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22060__I0 rbzero.wall_tracer.rcp_fsm.o_data\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17714_ _10904_ _10626_ _10899_ _10907_ _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_89_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14926_ _08360_ _07461_ _08732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_234_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18694_ _11673_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_10_i_clk_I clknet_5_4__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17645_ _10859_ rbzero.pov.ready_buffer\[4\] _10862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14857_ rbzero.tex_b1\[10\] _08541_ _08662_ _08663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_236_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13808_ rbzero.tex_r0\[13\] _07577_ _07619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14788_ _07603_ _08595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17576_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _10817_ _10818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19315_ rbzero.tex_b1\[36\] rbzero.tex_b1\[35\] _12115_ _12119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16527_ _09965_ _09977_ _09980_ _09918_ _09981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13739_ rbzero.tex_r0\[36\] _07545_ _07549_ _07550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18192__A1 _11301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19246_ rbzero.tex_b1\[6\] rbzero.tex_b1\[5\] _12078_ _12080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_16458_ _09895_ _09916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_128_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21079__A1 rbzero.traced_texVinit\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15409_ _09074_ _09129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16389_ rbzero.spi_registers.spi_buffer\[15\] _09853_ _09862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19177_ _11269_ _12020_ _12021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_235_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18128_ rbzero.debug_overlay.playerX\[5\] rbzero.wall_tracer.mapX\[5\] _11272_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13308__A2 _07035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14505__A1 _08264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18059_ _11202_ _11203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__21709__I _11331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21070_ _02142_ _02158_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23240__A2 _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20021_ _12687_ _12702_ _12793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__21251__A1 _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_171_Right_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_214_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13227__I _07040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24760_ _05490_ _05542_ _05544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21972_ rbzero.wall_tracer.rcp_fsm.o_data\[-4\] rbzero.wall_tracer.size\[4\] _03002_
+ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer10 _05032_ net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_1
Xrebuffer21 _05299_ net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21444__I _12647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_42_i_clk clknet_5_22__leaf_i_clk clknet_leaf_42_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_240_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer32 _05268_ net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_23711_ _11197_ _03043_ _04557_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20923_ _02011_ _02012_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24691_ _05469_ _05471_ _05473_ _05474_ _05475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_124_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26430_ _00340_ clknet_leaf_231_i_clk rbzero.spi_registers.spi_cmd\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23642_ rbzero.wall_tracer.visualWallDist\[2\] _12229_ _01980_ _04494_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_20854_ _01620_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26361_ _00271_ clknet_leaf_10_i_clk rbzero.spi_registers.buf_texadd1\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23573_ _04408_ _04425_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14992__A1 _06894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14058__I _07526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20785_ _12501_ _01376_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18183__A1 rbzero.map_overlay.i_otherx\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_i_clk clknet_5_23__leaf_i_clk clknet_leaf_57_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25312_ _06021_ _06023_ _06096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18183__B2 rbzero.map_overlay.i_othery\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22524_ _09938_ _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_135_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26292_ _00202_ clknet_leaf_228_i_clk rbzero.spi_registers.buf_floor\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25243_ _06026_ _06027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14744__A1 _08264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22455_ _02306_ _03344_ _03395_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_161_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21406_ _02484_ _02491_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_40_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25174_ _05929_ _05956_ _05958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22386_ _03327_ _08029_ _03331_ _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19584__I _12355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24125_ _04730_ _04908_ _04909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_21337_ _12522_ _01474_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24056_ _04839_ _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__18238__A2 _11381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21268_ _02348_ _02354_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23007_ _03685_ _03686_ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__21242__A1 _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_20219_ _12987_ _12989_ _12988_ _12557_ _12991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_60_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21199_ _02248_ _02286_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_217_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15760_ rbzero.spi_registers.texadd3\[6\] _09385_ _09389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24958_ _05727_ _05732_ _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_188_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13483__A1 rbzero.texV\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22742__A1 _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14711_ _07566_ _08518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23909_ rbzero.wall_tracer.rcp_fsm.o_data\[10\] rbzero.wall_tracer.stepDistX\[10\]
+ _04693_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15691_ _09334_ _09335_ _09337_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24889_ _05612_ _05618_ _05611_ _05673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_87_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_184_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_218_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_177_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14642_ rbzero.tex_g1\[45\] _07920_ _08450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_17430_ _10726_ _10724_ _10727_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_218_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_177_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26628_ _00538_ clknet_leaf_160_i_clk rbzero.tex_b0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_194_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14983__A1 _07979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14573_ _07764_ _07776_ _07789_ _08380_ _08381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_17361_ rbzero.pov.spi_buffer\[44\] _10676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_26559_ _00469_ clknet_leaf_67_i_clk rbzero.pov.spi_buffer\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18174__A1 rbzero.map_overlay.i_otherx\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19100_ _11918_ _11942_ _11943_ _11944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_60_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16312_ _09746_ _09804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13524_ _07322_ _07334_ _07335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17292_ rbzero.pov.spi_buffer\[27\] _10615_ _10624_ _10625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_231_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17921__A1 _08071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17279__I _10602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16243_ rbzero.spi_registers.buf_texadd2\[2\] _09743_ _09753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_97_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19031_ _11891_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16183__I _09671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13455_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] _07262_ _07266_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_82_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16174_ rbzero.spi_registers.buf_texadd1\[9\] _09696_ _09701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19674__A1 _12417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13386_ gpout0.vpos\[3\] _07197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19494__I rbzero.wall_tracer.stepDistX\[-6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15125_ _08908_ _08909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__20284__A2 _12788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19933_ _12704_ _12705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15056_ rbzero.spi_registers.spi_counter\[6\] rbzero.spi_registers.spi_counter\[5\]
+ _08849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_75_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13756__B _07549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_229_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14007_ rbzero.tex_r1\[24\] _07816_ _07817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_246_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19864_ _12263_ _12586_ _12636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18815_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] _11742_ _11744_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_235_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19795_ _12526_ _12528_ _12530_ _12567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_235_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18746_ _11702_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15958_ _09522_ _09528_ _09538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13474__A1 rbzero.traced_texVinit\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22733__A1 _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14909_ rbzero.tex_b1\[63\] _08568_ _08715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18677_ _11663_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15889_ _08924_ _09477_ _09486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17628_ _10848_ _10849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_187_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14974__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13777__A2 _07579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17559_ _10808_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__18165__A1 rbzero.map_overlay.i_mapdy\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22309__B _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20570_ rbzero.traced_texVinit\[2\] _01553_ _01661_ _01662_ _01663_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_156_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19229_ _12061_ _12051_ _12068_ _12069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14726__B2 _08522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_240_Right_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__23919__I _08813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22240_ _03110_ _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19665__A1 _12405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16479__A1 _09933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22171_ _03140_ _03153_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17140__A2 _10485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21122_ rbzero.wall_tracer.stepDistY\[10\] _12194_ _02209_ _02210_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_246_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_169_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24410__A1 _05186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25930_ _06710_ _06647_ _06712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14341__I rbzero.debug_overlay.facingY\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21053_ _02133_ _02141_ _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13701__A2 _07511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20004_ _12768_ _12772_ _12776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_25861_ _06628_ _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_126_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17652__I _10844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24812_ _05549_ _05595_ _05596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_158_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25792_ _06556_ _06574_ _06575_ _06576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_193_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22724__A1 _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21174__I _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24743_ _05526_ _05367_ _05527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_21955_ _02982_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15206__A2 _08975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20906_ _12662_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24674_ _05398_ _05458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_179_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21886_ _02927_ _02928_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26413_ _00323_ clknet_leaf_20_i_clk rbzero.spi_registers.buf_texadd3\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23625_ _04292_ _04382_ _04386_ _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_27393_ _01298_ clknet_leaf_108_i_clk rbzero.wall_tracer.stepDistX\[-9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20837_ _01923_ _01926_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14965__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26344_ _00254_ clknet_leaf_11_i_clk rbzero.spi_registers.buf_texadd0\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23556_ _04326_ _04332_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20768_ _12594_ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16706__A2 _10087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_213_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_213_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14717__A1 _07609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22507_ _03426_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_119_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26275_ _00185_ clknet_leaf_0_i_clk rbzero.spi_registers.texadd3\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23487_ _04262_ _04340_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20699_ _01741_ _01766_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_137_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25226_ _06009_ _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_137_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13240_ _07013_ _07018_ _07054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_150_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22438_ rbzero.wall_tracer.texu\[3\] _03361_ _03111_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25157_ _05936_ _05938_ _05940_ _05941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13171_ _06918_ _06985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22369_ _03307_ _03315_ _03316_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_131_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24108_ _04880_ _04891_ _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15142__A1 _08922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24401__A1 _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25088_ _05828_ _05861_ _05872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15693__A2 _09338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24039_ _04795_ rbzero.wall_tracer.rcp_fsm.operand\[3\] _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16930_ rbzero.debug_overlay.playerY\[1\] _10346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14251__I rbzero.debug_overlay.playerY\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21766__A2 _12185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16861_ _08049_ _10286_ _10174_ _10287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_53_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16642__A1 _10072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18600_ _11619_ _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15445__A2 _09151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16642__B2 _10049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15812_ rbzero.spi_registers.buf_texadd3\[20\] _09420_ _09427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19580_ rbzero.wall_tracer.stepDistX\[-8\] _12202_ _12351_ _12352_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_16792_ rbzero.pov.ready_buffer\[66\] _10201_ _10202_ _10225_ _10226_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_205_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22715__A1 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18531_ rbzero.tex_r0\[12\] rbzero.tex_r0\[11\] _11576_ _11580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_204_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15743_ _09374_ _09376_ _09372_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_18462_ _11540_ _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_158_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15674_ _09289_ _09325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_185_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19489__I _12260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17413_ rbzero.pov.spi_buffer\[57\] _10715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14625_ rbzero.tex_g1\[33\] _07635_ _08433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__18393__I _11479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18393_ _11479_ _11501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14556_ _07433_ _08364_ _07447_ _08365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17344_ _10661_ _10653_ _10663_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_101_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13507_ _07316_ _07317_ _07318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_181_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17275_ _10611_ _10612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14487_ _08287_ _08290_ _08293_ _08294_ _08295_ _08296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_71_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19014_ _11871_ _11882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16226_ rbzero.spi_registers.buf_texadd1\[23\] _09730_ _09739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13438_ gpout0.vpos\[9\] _07249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_77_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer1 _05560_ net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20257__A2 _13028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_248_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16157_ _09660_ _09689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13369_ gpout0.vpos\[0\] _07181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15108_ _08857_ _08892_ rbzero.spi_registers.spi_counter\[3\] _08896_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16088_ _08973_ _09635_ _09636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_244_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19916_ _12472_ _12688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15039_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\] _08832_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_209_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21757__A2 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_209_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19847_ _12476_ _12470_ _12411_ _12561_ _12619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_242_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_236_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17472__I _10757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19778_ _12275_ _12495_ _12550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21509__A2 _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18729_ _11692_ _11693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__24171__A3 _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17189__A2 _10547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21740_ _02779_ _02794_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_121_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24459__A1 _05242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21671_ _11360_ _12020_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23410_ _04146_ _04263_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20622_ _01597_ _01598_ _01713_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_188_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24390_ _04866_ _04889_ _05060_ _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_190_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23341_ _04047_ _04194_ _04195_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_11_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21693__A1 _11260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20553_ _01644_ _01486_ _01645_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_34_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26060_ _06632_ _06615_ _06830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_190_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23272_ _04008_ _04009_ _04012_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14175__A2 _07189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20484_ _12301_ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25011_ _05520_ _05580_ _05582_ _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_22223_ _03193_ _03195_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_132_i_clk_I clknet_5_15__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22154_ _10151_ _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_132_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21105_ _02189_ _02192_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_160_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26962_ _00872_ clknet_leaf_111_i_clk rbzero.texV\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_22085_ _10048_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21748__A2 _09982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25913_ _05171_ _06695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21036_ _02107_ _02124_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_22_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19810__A1 _12576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26893_ _00803_ clknet_leaf_176_i_clk rbzero.tex_r0\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_195_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25844_ _05126_ _06628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_214_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25775_ _06557_ _06558_ _06559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__19811__B _12267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22987_ _03844_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_201_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24726_ _05240_ _05272_ _05446_ _05510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_139_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21938_ _10478_ _02959_ _09934_ _10484_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_57_i_clk_I clknet_5_23__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27445_ _01350_ clknet_leaf_69_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24657_ _05411_ _05440_ _05441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_26_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21869_ _08126_ _10466_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_139_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14410_ rbzero.tex_g0\[24\] _08207_ _08219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23608_ _04321_ _01972_ _04419_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_155_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15390_ _09064_ _09115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_27376_ _01281_ clknet_leaf_81_i_clk rbzero.wall_tracer.trackDistY\[-4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24588_ _05371_ _05350_ _05372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_93_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14341_ rbzero.debug_overlay.facingY\[-1\] _08151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_26327_ _00237_ clknet_leaf_234_i_clk rbzero.spi_registers.buf_mapdy\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__21684__A1 _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23539_ _04284_ _04376_ _04391_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17060_ _10448_ _10449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14272_ rbzero.debug_overlay.facingX\[-9\] _08082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26258_ _00168_ clknet_leaf_240_i_clk rbzero.spi_registers.texadd3\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16011_ _08950_ _09574_ _09578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25209_ _05976_ _05989_ _05992_ _05993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_TAPCELL_ROW_189_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13223_ rbzero.spi_registers.texadd3\[23\] _07014_ _07036_ rbzero.spi_registers.texadd2\[23\]
+ _07030_ rbzero.spi_registers.texadd1\[23\] _07037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26189_ _00099_ clknet_leaf_236_i_clk rbzero.spi_registers.texadd0\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold48_I i_gpout1_sel[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13154_ _06966_ _06967_ _06968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_103_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13085_ _06899_ _06900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_17962_ rbzero.map_rom.i_col\[4\] _11106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_236_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21739__A2 _11420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19701_ _12472_ _12423_ _12473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_16913_ _10209_ _10331_ _10332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_109_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17893_ _08075_ rbzero.wall_tracer.rayAddendX\[10\] _11037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_205_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20411__A2 _12379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19632_ _11953_ _11998_ _10317_ _12003_ _12404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_16844_ _07167_ _10271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_233_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19563_ _12315_ _12318_ _12328_ _12334_ _12335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_16775_ _10165_ _10210_ _10211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_204_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13987_ _07793_ _07794_ _07795_ _07796_ _07797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18514_ _11570_ _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15726_ _09352_ _09364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19494_ rbzero.wall_tracer.stepDistX\[-6\] _12266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_158_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18337__B _10751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18445_ rbzero.tex_g1\[39\] rbzero.tex_g1\[38\] _11528_ _11531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15657_ rbzero.spi_registers.texadd2\[4\] _09303_ _09312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_200_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14608_ rbzero.tex_g1\[7\] _07597_ _08416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__19868__A1 rbzero.wall_tracer.size\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18376_ rbzero.tex_g1\[9\] rbzero.tex_g1\[8\] _11491_ _11492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_145_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15588_ rbzero.spi_registers.texadd1\[10\] _09255_ _09261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17327_ rbzero.pov.spi_buffer\[36\] _10650_ _10646_ _10651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14156__I _07425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14539_ rbzero.tex_g0\[57\] _07894_ _08348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18391__I1 rbzero.tex_g1\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22373__I _12577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17258_ _10564_ _10599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24613__A1 _05098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13995__I _07804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16209_ _08997_ _09721_ _09727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13904__A2 _07060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17189_ rbzero.pov.spi_buffer\[1\] _10547_ _10174_ _10548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_183_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15657__A2 _09303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13944__B _07754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22910_ _03634_ _03637_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14759__C _08565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23890_ rbzero.wall_tracer.rcp_fsm.o_data\[1\] rbzero.wall_tracer.stepDistX\[1\]
+ _04685_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__17135__C _09441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__23932__I _10491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22841_ _03676_ _03699_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_169_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13235__I _07040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25560_ _06343_ _06333_ _06344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_182_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22772_ _02744_ _03630_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_195_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24511_ _05165_ _05295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__21902__A2 _11069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21723_ _10249_ _02773_ _02778_ _02780_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_231_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25491_ _06272_ _06082_ _06123_ _06143_ _06275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_38_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25859__I _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24442_ _05008_ _05018_ _05025_ _05225_ _05226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_27230_ _01135_ clknet_leaf_86_i_clk rbzero.wall_tracer.rcp_fsm.i_data\[-7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21654_ _10255_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20605_ _01695_ _01696_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_47_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27161_ _01066_ clknet_leaf_204_i_clk rbzero.map_rom.f3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24373_ _05059_ _05153_ _05156_ _05157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_145_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14066__I _07511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21585_ _02668_ _02669_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_26112_ _00022_ clknet_leaf_242_i_clk rbzero.spi_registers.spi_buffer\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23324_ _03811_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_201_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20536_ _01379_ _01476_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_61_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27092_ _01002_ clknet_leaf_140_i_clk rbzero.tex_b1\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_201_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17377__I _10665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26043_ _05006_ _06691_ _06816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23255_ _04027_ _04109_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20467_ _01464_ _01543_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13838__C _07648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22206_ _03161_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_162_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23186_ _04040_ _04041_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20398_ _01404_ _01441_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22137_ _03125_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__20641__A2 _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22068_ _03067_ _03054_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26945_ _00855_ clknet_leaf_178_i_clk rbzero.tex_r1\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_234_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21019_ _01963_ _01964_ _01984_ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_50_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13910_ rbzero.map_overlay.i_othery\[0\] _07721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_233_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26876_ _00786_ clknet_leaf_165_i_clk rbzero.tex_r0\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14890_ rbzero.tex_b1\[40\] _08518_ _08696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_221_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_221_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25827_ _06608_ _06609_ _06610_ _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13841_ rbzero.tex_r0\[18\] _07459_ _07343_ _07652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_202_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23343__A1 _12950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15820__A2 _09032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16560_ rbzero.debug_overlay.vplaneY\[0\] _09992_ _10012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13772_ _07582_ _07583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25758_ _06488_ _06502_ _06541_ _06542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15511_ rbzero.spi_registers.buf_texadd0\[15\] _09030_ _09203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24709_ _05440_ _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_168_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16491_ _09945_ _09946_ _09947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25689_ _06461_ _06473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_195_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18230_ _09056_ _11343_ _11320_ rbzero.map_overlay.i_mapdx\[3\] _11373_ _11374_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_27428_ _01333_ clknet_leaf_83_i_clk rbzero.wall_tracer.rcp_fsm.operand\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__14387__A2 _08194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15442_ _09153_ _09154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_65_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_43_Left_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18161_ _11300_ _11260_ _11251_ _11304_ _11305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_27359_ _01264_ clknet_leaf_106_i_clk rbzero.wall_tracer.trackDistX\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15373_ rbzero.floor_leak\[2\] _09101_ _09102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17112_ rbzero.pov.ready_buffer\[0\] _10489_ _10490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14139__A2 _07940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14324_ _08133_ _08134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18092_ _11146_ _11235_ _11236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17043_ _10433_ _10435_ _10436_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14255_ _08021_ _08033_ _08065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13206_ _07008_ _07020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22082__A1 _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14186_ _07991_ _07995_ _07996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13137_ _06950_ _06951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_18994_ _11870_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_209_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19435__C _12206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_206_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20441__I _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17945_ _11087_ _11066_ _11088_ _11089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13068_ gpout0.hpos\[5\] _06884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_206_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17876_ rbzero.wall_tracer.rayAddendX\[3\] _11020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23752__I _12035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19615_ _12260_ _12386_ _12387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16827_ _10249_ _10165_ _10256_ _10257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18846__I _11737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14075__A1 _07841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19546_ _12317_ _12318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_239_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16758_ _08172_ _08180_ rbzero.debug_overlay.playerX\[-9\] rbzero.debug_overlay.playerX\[-6\]
+ _10196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_49_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_215_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15709_ rbzero.spi_registers.texadd2\[17\] _09350_ _09351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19477_ rbzero.wall_tracer.side _12249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16689_ _10066_ _10131_ _10133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18428_ rbzero.tex_g1\[32\] rbzero.tex_g1\[31\] _11517_ _11521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14378__A2 _08023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21648__A1 _08106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18359_ _11482_ _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_173_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20320__A1 _12486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21370_ _02454_ _02455_ _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13338__B1 _07149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20321_ _12495_ _12519_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22073__A1 _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23040_ _03892_ _03893_ _03896_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_20252_ _13023_ _13024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_247_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14550__A2 _08358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20183_ _12953_ _12938_ _12954_ _12955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__25011__A1 _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_216_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25562__A2 _05605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24991_ _05563_ _05564_ _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_243_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22376__A2 _12173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26730_ _00640_ clknet_leaf_32_i_clk rbzero.pov.ready_buffer\[60\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23942_ _04742_ _04743_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input22_I i_reg_sclk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23873_ _12499_ _04686_ _04697_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_162_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26661_ _00571_ clknet_leaf_158_i_clk rbzero.tex_b0\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__18756__I _11692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25612_ _06357_ _06364_ _06396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22824_ _03681_ _03682_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__20139__A1 rbzero.wall_tracer.size\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26592_ _00502_ clknet_leaf_33_i_clk rbzero.pov.spi_buffer\[61\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25543_ _06326_ _06296_ _06327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_22755_ _03611_ _03614_ _03615_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_183_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21706_ _11397_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25474_ _06104_ _06105_ _06258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_192_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14369__A2 _08011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22686_ _11199_ _03522_ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24425_ _04896_ _05091_ _05111_ _05209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_27213_ _01118_ clknet_leaf_79_i_clk rbzero.wall_tracer.stepDistY\[-2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_191_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21637_ _02708_ _02712_ _02713_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22300__A2 _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27144_ _00000_ clknet_leaf_74_i_clk rbzero.wall_tracer.rcp_fsm.state\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24356_ _05133_ net74 _05139_ _05114_ _05140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_23_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21568_ _02651_ _02652_ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_133_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23307_ _03651_ _04157_ _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_185_Right_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20519_ _12263_ _01534_ _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_169_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27075_ _00985_ clknet_leaf_138_i_clk rbzero.tex_b1\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24287_ net49 _05066_ _05068_ _05070_ _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_133_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21499_ _02495_ _02517_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_169_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14040_ rbzero.tex_r1\[20\] _07843_ _07850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26026_ _06758_ rbzero.wall_tracer.rcp_fsm.o_data\[-2\] _06759_ _06801_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23238_ _03985_ _03986_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_63_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23169_ _04023_ _04024_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_182_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_223_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24356__A3 _05139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15991_ _08980_ _09562_ _09563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_147_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15355__I _09054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17730_ _10913_ rbzero.pov.ready_buffer\[33\] _10918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14942_ _08743_ reg_hsync _08746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26928_ _00838_ clknet_leaf_172_i_clk rbzero.tex_r1\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_17661_ _10865_ _10576_ _10868_ _10871_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_243_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_26859_ _00769_ clknet_leaf_187_i_clk rbzero.tex_r0\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14873_ _08654_ _08678_ _08355_ _08679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_215_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19400_ _12171_ _12172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__17794__A2 rbzero.pov.ready_buffer\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16612_ _10041_ _10042_ _10059_ _10060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_201_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13824_ _07628_ _07635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17592_ rbzero.tex_b0\[52\] rbzero.tex_b0\[51\] _10823_ _10827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_67_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19331_ rbzero.tex_b1\[43\] rbzero.tex_b1\[42\] _12125_ _12128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_197_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16543_ _09982_ _09987_ _09995_ _09996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13755_ _07486_ _07566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15090__I _08881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19262_ rbzero.tex_b1\[13\] rbzero.tex_b1\[12\] _12088_ _12089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__20550__A1 _12235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16474_ _09929_ _09930_ _09931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13686_ _07485_ _07490_ _07491_ _07494_ _07496_ _07497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_26_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18213_ _11347_ _11263_ _11334_ _11308_ _11357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_234_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15425_ rbzero.color_floor\[3\] _08879_ _09141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_234_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19193_ _11396_ _12037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_171_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18144_ rbzero.wall_tracer.visualWallDist\[-3\] _11288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20436__I _12311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20302__A1 _12984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15356_ _09087_ _09088_ _09089_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14780__A2 _07629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14307_ rbzero.debug_overlay.vplaneY\[-3\] _08117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_152_Right_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18075_ _11198_ _11199_ _11201_ _11203_ _11208_ _11218_ _11219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_180_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15287_ rbzero.spi_registers.buf_othery\[0\] _09038_ _09039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_123_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17026_ _10392_ _10423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14238_ rbzero.debug_overlay.playerY\[-9\] _08048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_123_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19446__B _12182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_179_i_clk_I clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14169_ _07686_ _07979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_111_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18977_ _11850_ _11861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_226_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19960__I _12731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17928_ _11004_ _11072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__24578__I _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17859_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] _11003_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_231_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14048__A1 rbzero.tex_r1\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20870_ _01946_ _01959_ _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15796__A1 rbzero.spi_registers.texadd3\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14599__A2 _07857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19529_ _12198_ _12301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_147_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22540_ rbzero.wall_tracer.visualWallDist\[-5\] _03443_ _03444_ rbzero.traced_texa\[-5\]
+ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_220_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22471_ _08033_ _03402_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24210_ _04930_ _04952_ _04957_ _04965_ _04994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_8_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21422_ _12788_ _02292_ _02387_ _02507_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_25190_ _05973_ _05974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24141_ _04904_ _04907_ _04909_ _04924_ _04925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_31_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21353_ _02317_ _02439_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20304_ _13011_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_142_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24072_ _04801_ _04803_ _04855_ _04810_ _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_31_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21284_ _02113_ _02237_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23023_ _03775_ _03880_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20235_ _12904_ _12905_ _13007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_228_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19462__A2 _11099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20166_ _12937_ _12938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_228_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14287__A1 _08096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20097_ _12611_ _12655_ _12869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_24974_ _05502_ _05518_ _05553_ _05758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_157_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26713_ _00623_ clknet_leaf_29_i_clk rbzero.pov.ready_buffer\[43\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_243_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_23925_ rbzero.wall_tracer.rcp_fsm.operand\[-9\] _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_157_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26644_ _00554_ clknet_leaf_146_i_clk rbzero.tex_b0\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23856_ _04684_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_142_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22807_ _03649_ _03665_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26575_ _00485_ clknet_leaf_27_i_clk rbzero.pov.spi_buffer\[44\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20999_ _12696_ _01982_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23787_ _04527_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_179_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24437__B _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25526_ _06309_ _06124_ _06310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_196_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15539__A1 rbzero.spi_registers.buf_texadd0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13540_ rbzero.floor_leak\[5\] _07325_ _07349_ rbzero.floor_leak\[4\] _07351_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_22738_ rbzero.wall_tracer.trackDistX\[-1\] _01993_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13471_ _07278_ _07281_ _07282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22669_ rbzero.wall_tracer.stepDistX\[-8\] _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25457_ _06222_ _06224_ _06229_ _06231_ _06241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_164_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_216_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15210_ rbzero.spi_registers.spi_buffer\[15\] _08975_ _08979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24408_ _05186_ _05081_ _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_192_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18154__C _11297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14762__A2 _08568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16190_ rbzero.spi_registers.buf_texadd1\[13\] _09707_ _09713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25388_ _06171_ _06135_ _06172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__19150__A1 _08160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15141_ rbzero.spi_registers.spi_buffer\[3\] _08922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27127_ _01037_ clknet_leaf_121_i_clk rbzero.traced_texVinit\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24339_ _05121_ _05122_ _05123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22037__A1 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15072_ _08864_ _08865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_27058_ _00968_ clknet_leaf_133_i_clk rbzero.tex_b1\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_95_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14514__A2 _08317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_180_i_clk_I clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14023_ rbzero.tex_r1\[17\] _07832_ _07587_ _07833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18900_ rbzero.traced_texa\[7\] _07267_ _11813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26009_ _06678_ _06786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_120_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19880_ _12573_ _12652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_247_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_18831_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] _11757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_235_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15085__I _08876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18762_ _11711_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15974_ _09437_ _08831_ _09550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_199_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_199_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17713_ _10906_ rbzero.pov.ready_buffer\[27\] _10907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22060__I1 rbzero.wall_tracer.stepDistY\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14925_ _08364_ _08729_ _08730_ _07963_ _07440_ _08731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_18693_ rbzero.tex_r1\[17\] rbzero.tex_r1\[16\] _11672_ _11673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_231_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15813__I _08931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17767__A2 rbzero.pov.ready_buffer\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22760__A2 rbzero.wall_tracer.stepDistX\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17644_ _10850_ _10861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14856_ rbzero.tex_b1\[11\] _08448_ _08662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_232_i_clk clknet_5_0__leaf_i_clk clknet_leaf_232_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_5_18__f_i_clk clknet_3_4_0_i_clk clknet_5_18__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_236_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13807_ rbzero.tex_r0\[14\] _07617_ _07462_ _07618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_203_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17575_ _10801_ _10817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_221_Right_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14787_ _08304_ _08593_ _08594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13333__I _07046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19314_ _12118_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16526_ _09902_ _09979_ _09980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13738_ _07443_ _07549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19245_ _12079_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16457_ _09914_ _09915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_247_i_clk clknet_5_1__leaf_i_clk clknet_leaf_247_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13669_ _07479_ _07480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14202__A1 _07373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24265__A2 _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25957__I _06737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22276__A1 _11190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15408_ _09114_ _09127_ _09128_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_19176_ rbzero.map_rom.c6 _12007_ _12020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14753__A2 _08494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16388_ rbzero.spi_registers.buf_texadd3\[15\] _09851_ _09861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18127_ rbzero.debug_overlay.playerX\[1\] rbzero.map_rom.f3 _11271_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15339_ _09077_ _09078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18058_ rbzero.wall_tracer.trackDistY\[-8\] _11202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22381__I _12907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17009_ _08073_ _10410_ _10411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20020_ _12674_ _12788_ _12789_ _12791_ _12792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_10_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21251__A2 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21971_ _02991_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_179_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16819__I _07694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer11 _05032_ net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_222_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer22 _04849_ net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23710_ _04555_ _04556_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_20922_ _01877_ _01878_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xrebuffer33 _05190_ net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_24690_ _05306_ _05461_ _05407_ _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_124_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20853_ _01937_ _01942_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_166_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23641_ _04222_ _01972_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23572_ _04423_ _04424_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26360_ _00270_ clknet_leaf_10_i_clk rbzero.spi_registers.buf_texadd1\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20784_ _12472_ _01468_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22523_ _03435_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25311_ _06021_ _06023_ _06095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26291_ _00201_ clknet_leaf_230_i_clk rbzero.spi_registers.buf_floor\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16194__A1 _08980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25242_ _06025_ _06015_ _06026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22454_ _02167_ _03393_ _03394_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__19132__A1 _08152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21405_ _12837_ _02489_ _02490_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_17_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25173_ _05929_ _05956_ _05957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_199_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22385_ _12907_ _10176_ _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22019__A1 _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24124_ _04724_ _04718_ _04812_ _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18730__I1 rbzero.tex_r1\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21336_ _02227_ _02422_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22291__I _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24055_ _04833_ _04836_ _04838_ _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__24964__B1 _05746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21267_ _02350_ _02353_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23006_ _03859_ _03863_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_20218_ _12987_ _12988_ _12557_ _12989_ _12990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_21_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21198_ _02266_ _02285_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__23519__A1 _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14023__B _07587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20149_ _12904_ _12905_ _12920_ _12921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_144_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19199__A1 _11131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13862__B _07670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24957_ _05696_ _05739_ _05722_ _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14680__A1 _08198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24319__I0 _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14710_ rbzero.tex_b0\[61\] _08233_ _08517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23908_ _03026_ _04687_ _04716_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_213_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15690_ _09336_ _09337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24888_ _05671_ _05672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22667__S _11400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_127_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14641_ rbzero.tex_g1\[47\] _08448_ _07917_ _08449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26627_ _00537_ clknet_leaf_160_i_clk rbzero.tex_b0\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XTAP_TAPCELL_ROW_177_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23839_ _04668_ _04669_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_194_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17360_ _10673_ _10666_ _10675_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_170_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26558_ _00468_ clknet_leaf_67_i_clk rbzero.pov.spi_buffer\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14572_ _07767_ _07798_ _08380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14983__A2 _07707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18174__A2 rbzero.map_rom.f4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16311_ rbzero.spi_registers.buf_texadd2\[20\] _09802_ _09803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25509_ _06151_ _06158_ _06293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_60_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13523_ _07301_ _07302_ _07334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17291_ _10611_ _10624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_153_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26489_ _00399_ clknet_leaf_57_i_clk rbzero.debug_overlay.facingX\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_231_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19030_ rbzero.tex_g0\[48\] rbzero.tex_g0\[47\] _11887_ _11891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_97_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16242_ _09751_ _09752_ _09750_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13454_ _07262_ _07263_ _07264_ _07265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13385_ gpout0.vpos\[4\] _07196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16173_ _09697_ _09699_ _09700_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15124_ _08805_ _08908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_51_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20714__I _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17295__I _10602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19932_ _12553_ _12704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15055_ rbzero.spi_registers.spi_counter\[4\] rbzero.spi_registers.spi_counter\[3\]
+ rbzero.spi_registers.spi_counter\[2\] _08848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_75_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_229_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_246_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14006_ _07804_ _07816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19863_ _12547_ _12551_ _12634_ _12635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_208_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22430__A1 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18814_ _11738_ _11743_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19794_ _12552_ _12565_ _12566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__15999__A1 _09525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16660__A2 _10020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18745_ rbzero.tex_r1\[40\] rbzero.tex_r1\[39\] _11698_ _11702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15957_ rbzero.spi_registers.buf_vshift\[3\] _09531_ _09537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_222_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14671__A1 _07888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_171_i_clk clknet_5_11__leaf_i_clk clknet_leaf_171_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13474__A2 rbzero.spi_registers.vshift\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14908_ _08304_ _08708_ _08713_ _08714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_78_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18676_ rbzero.tex_r1\[10\] rbzero.tex_r1\[9\] _11661_ _11663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15888_ rbzero.spi_registers.buf_leak\[2\] _09482_ _09485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17627_ _10847_ _10848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_106_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14839_ _08641_ _08642_ _08644_ _08255_ _08532_ _08645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_77_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17558_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _10807_ _10808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_186_i_clk clknet_5_8__leaf_i_clk clknet_leaf_186_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__14974__A2 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13998__I _07520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18165__A2 _11252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16509_ _09956_ _09940_ _09964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17489_ _10768_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19228_ rbzero.wall_tracer.mapY\[9\] _12062_ _12065_ _12068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15923__A1 _08965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19114__A1 _08153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14108__B _07917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19159_ _12000_ _12002_ _11949_ _12003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_5_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__22325__B _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22170_ rbzero.wall_tracer.rcp_fsm.i_data\[0\] _03144_ _03152_ _03153_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21121_ _12194_ _02208_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19417__A2 _12169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_124_i_clk clknet_5_18__leaf_i_clk clknet_leaf_124_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21052_ _02135_ _02140_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_10_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22421__A1 _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13238__I _06905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20003_ _12673_ _12774_ _12775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_10_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22972__A2 _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25860_ _06638_ _06640_ _06641_ _06642_ _06628_ _06643_ _06644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__20983__A1 _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24811_ _05554_ _05594_ _05595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__16651__A2 _09928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25791_ _06553_ _06568_ _06575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_139_i_clk clknet_5_15__leaf_i_clk clknet_leaf_139_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23921__A1 _11392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15453__I _09111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24742_ _05334_ _05526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21954_ rbzero.wall_tracer.rcp_fsm.o_data\[-9\] _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_179_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_25__f_i_clk_I clknet_3_6_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20905_ _12668_ _01994_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24673_ _05392_ _05455_ _05456_ _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21885_ _08121_ _08125_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26412_ _00322_ clknet_leaf_21_i_clk rbzero.spi_registers.buf_texadd3\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20836_ _12969_ _01924_ _01925_ _12787_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_23624_ _04372_ _04392_ _04368_ _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__22488__A1 rbzero.wall_tracer.size\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27392_ _01297_ clknet_leaf_107_i_clk rbzero.wall_tracer.stepDistX\[-10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26343_ _00253_ clknet_leaf_11_i_clk rbzero.spi_registers.buf_texadd0\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__16284__I _09761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23555_ _04400_ _04407_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_20767_ _01681_ _01685_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_42_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_213_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_213_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22506_ rbzero.wall_tracer.size\[9\] _03423_ _03424_ _07353_ _03426_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_108_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23486_ _04265_ _04339_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_135_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_26274_ _00184_ clknet_leaf_0_i_clk rbzero.spi_registers.texadd3\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20698_ _01742_ _01765_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25225_ _05521_ _06009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_190_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22437_ _03351_ _03378_ _03379_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_134_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13170_ _06979_ _06983_ _06984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25156_ _05936_ _05938_ _05939_ _05940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_22368_ rbzero.mapdxw\[1\] _03307_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24107_ _04882_ _04885_ _04888_ _04890_ _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_21319_ _02259_ _02263_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25087_ _05825_ _05826_ _05870_ _05863_ _05871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_22299_ _11178_ _03254_ _03259_ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_150_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24401__A2 _05183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24038_ _04813_ _04814_ _04815_ _04816_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_102_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__16890__A2 _10310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22963__A2 _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16860_ _10281_ _10286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15811_ rbzero.spi_registers.texadd3\[20\] _09418_ _09426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16791_ _10194_ _10224_ _10225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_244_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25989_ _05171_ _05030_ _06768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_244_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18919__A1 _11456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18530_ _11579_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22715__A2 _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15742_ rbzero.spi_registers.buf_texadd3\[1\] _09375_ _09376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_220_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18461_ rbzero.tex_g1\[46\] rbzero.tex_g1\[45\] _11538_ _11540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_213_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15673_ rbzero.spi_registers.buf_texadd2\[8\] _09317_ _09324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_198_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17412_ _10711_ _10713_ _10714_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14624_ rbzero.tex_g1\[35\] _07855_ _07613_ _08432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18392_ _11500_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14956__A2 _08753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17343_ rbzero.pov.spi_buffer\[40\] _10662_ _10659_ _10663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14555_ _07434_ _08364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13506_ _07261_ _07265_ _07317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17274_ _06897_ _10611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14486_ _07496_ _08295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_19013_ _11881_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16225_ _09737_ _09738_ _09734_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13437_ _07193_ _07247_ _07248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xrebuffer2 _04813_ net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_248_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_248_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22651__A1 _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16156_ _08926_ _09687_ _09688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13368_ gpout0.vpos\[1\] _07180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_41_i_clk clknet_5_16__leaf_i_clk clknet_leaf_41_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_23_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15107_ _08894_ _08895_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_16087_ _09600_ _09635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_228_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13299_ _07110_ _07112_ _07113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19915_ _12684_ _12686_ _12687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15038_ _08830_ _08831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_236_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_209_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_56_i_clk clknet_5_23__leaf_i_clk clknet_leaf_56_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19846_ _12470_ _12411_ _12561_ _12475_ _12618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_108_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19777_ _12548_ _12491_ _12549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16989_ _10395_ _10396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__23903__A1 _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18728_ _11649_ _11692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_88_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19583__A1 _08041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18659_ _11653_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_121_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25656__A1 _05333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24459__A2 _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20193__A2 _12223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21670_ _11334_ _02729_ _02735_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20621_ _12706_ _01712_ _01599_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19886__A2 _12301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13521__I _07331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23340_ _04171_ _04070_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20552_ _01482_ _01485_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_154_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23271_ _04008_ _04009_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20483_ _01574_ _01575_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_119_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer25_I _05098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22222_ _03182_ _03183_ _03194_ _03165_ rbzero.wall_tracer.rcp_fsm.i_data\[10\] _03195_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_25010_ _05584_ _05586_ _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_89_Left_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22153_ _03119_ _03139_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_3_7_0_i_clk clknet_0_i_clk clknet_3_7_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__24270__B _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21104_ _02190_ _02191_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_100_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26961_ _00871_ clknet_leaf_114_i_clk rbzero.texV\[-9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_22084_ _03078_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_196_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17663__I _10872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25912_ _06902_ _06694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21035_ _02110_ _02123_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_245_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26892_ _00802_ clknet_leaf_176_i_clk rbzero.tex_r0\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_227_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19810__A2 _12578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25843_ _06626_ _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_98_Left_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_25774_ _05976_ _05989_ _06558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_198_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22986_ _12662_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_241_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24725_ _05407_ _05307_ _05509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21937_ _10483_ _11092_ _02975_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_210_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27444_ _01349_ clknet_leaf_73_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24656_ _05362_ _05439_ _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_26_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21868_ _02910_ _02911_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_139_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23607_ _04451_ _04454_ _04458_ _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_38_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27375_ _01280_ clknet_leaf_81_i_clk rbzero.wall_tracer.trackDistY\[-5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20819_ _01904_ _01908_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_24587_ _05129_ _05371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_154_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21799_ _09989_ _02847_ _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_166_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14340_ _08149_ _08078_ _08150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26326_ _00236_ clknet_leaf_234_i_clk rbzero.spi_registers.buf_mapdy\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_231_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23538_ _04381_ _04390_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_231_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26072__A1 _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17838__I _07166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14271_ rbzero.debug_overlay.facingX\[-7\] _08081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26257_ _00167_ clknet_leaf_239_i_clk rbzero.spi_registers.texadd3\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23469_ _04221_ _04224_ _04322_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_243_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26609__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16010_ rbzero.spi_registers.buf_mapdy\[3\] _09572_ _09577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25208_ _05988_ _05991_ _05992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13222_ _07009_ _07036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26188_ _00098_ clknet_leaf_242_i_clk rbzero.spi_registers.texadd0\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25139_ _05920_ _05922_ _05923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13153_ rbzero.texu_hot\[1\] _06961_ _06967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_55_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17961_ _11103_ _11104_ _11105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13084_ _06898_ _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_226_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19700_ _12471_ _12472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16912_ _07698_ _10330_ _10331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_236_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17892_ _08075_ rbzero.wall_tracer.rayAddendX\[10\] _11036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_233_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_218_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19631_ _12402_ _12403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16843_ _10268_ _10270_ _10214_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_217_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14626__A1 rbzero.tex_g1\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19562_ rbzero.wall_tracer.stepDistX\[-7\] _12161_ _12333_ _12334_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_16774_ rbzero.pov.ready_buffer\[64\] _10208_ _10209_ _10210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_205_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13986_ _07219_ _06875_ _07796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19565__A1 _08042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18513_ rbzero.tex_r0\[4\] rbzero.tex_r0\[3\] _11566_ _11570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15725_ rbzero.spi_registers.texadd2\[21\] _09362_ _09363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19493_ _12261_ _12264_ _12265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_198_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18444_ _11530_ _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_158_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15656_ _09310_ _09311_ _09301_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_199_Right_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14607_ _08411_ _08412_ _08414_ _07867_ _07868_ _08415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_8_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18375_ _11480_ _11491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__21124__A1 _12231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15587_ _09256_ _09260_ _09253_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_83_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17326_ _10649_ _10650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_173_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14538_ rbzero.tex_g0\[56\] _07901_ _08347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20883__B1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17257_ rbzero.pov.spi_buffer\[18\] _10598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_183_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14469_ rbzero.tex_g0\[38\] _08277_ _08278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25965__I _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16208_ rbzero.spi_registers.buf_texadd1\[18\] _09719_ _09726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13365__A1 _07176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17188_ _10546_ _10547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16139_ _09674_ _09675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_228_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24377__A1 _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18579__I _11564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_242_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19829_ _12567_ _12600_ _12601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_166_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22840_ _03680_ _03698_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_224_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21733__I _11409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22771_ _03627_ _03628_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13840__A2 _07576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24510_ _05292_ _05291_ _05293_ _05294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_52_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21722_ _02779_ _11118_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_25490_ _05521_ _06024_ _05967_ _06274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_8_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_166_Right_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24441_ _05041_ _05042_ _05136_ _05043_ _05122_ _05088_ _05225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_21653_ _02692_ _08194_ _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13251__I _07040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20604_ _12423_ _12646_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_27160_ _01065_ clknet_leaf_204_i_clk rbzero.map_rom.f4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_24372_ _05105_ _05106_ _05154_ _05155_ _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_21584_ _02261_ _01380_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22564__I _09973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26111_ _00021_ clknet_leaf_242_i_clk rbzero.spi_registers.spi_buffer\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20535_ _01477_ _01489_ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23323_ _04065_ _04177_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__16542__A1 _09989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27091_ _01001_ clknet_leaf_140_i_clk rbzero.tex_b1\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_134_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13356__A1 _07164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_226_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26042_ _06720_ _06725_ _06815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22615__A1 _11131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13356__B2 _07167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23254_ _04027_ _04109_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_20466_ _01464_ _01543_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19873__I _12644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15178__I _08933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22205_ _03176_ _03181_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23185_ _02595_ _03660_ _04039_ _12428_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_20397_ _01465_ _01490_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_203_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22136_ _03087_ _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14305__B1 _08016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17393__I _10665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_184_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22067_ rbzero.wall_tracer.stepDistY\[5\] _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_199_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26944_ _00854_ clknet_leaf_177_i_clk rbzero.tex_r1\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_21018_ _01921_ _01928_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26875_ _00785_ clknet_leaf_164_i_clk rbzero.tex_r0\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_50_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_221_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25826_ _06573_ _06589_ _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_221_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13840_ rbzero.tex_r0\[19\] _07576_ _07651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19541__C _12005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23343__A2 _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25757_ _06487_ _06540_ _06541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13771_ _07481_ _07582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_230_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22969_ _03823_ _03826_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15510_ _09200_ _09201_ _09202_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24708_ _05411_ _05492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16490_ _09942_ _08099_ _08100_ _09946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_69_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25688_ _06470_ _06471_ _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_195_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27427_ _01332_ clknet_leaf_83_i_clk rbzero.wall_tracer.rcp_fsm.operand\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15441_ _08883_ _09153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_24639_ _05409_ _05412_ _05414_ _05423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_167_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16781__A1 rbzero.debug_overlay.playerX\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18160_ _11301_ _11303_ _11304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_27358_ _01263_ clknet_leaf_106_i_clk rbzero.wall_tracer.trackDistX\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15372_ _09074_ _09101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21657__A2 _08491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17111_ _10395_ _10489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26309_ _00219_ clknet_leaf_233_i_clk rbzero.spi_registers.buf_vshift\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14323_ rbzero.debug_overlay.vplaneX\[-4\] _08133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_208_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18091_ _11159_ _11233_ _11234_ _11235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27289_ _01194_ clknet_leaf_210_i_clk gpout0.hpos\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13347__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17042_ _10385_ _10436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22606__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14254_ _08063_ _08064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13205_ _07013_ _07018_ _07019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_14185_ gpout0.hpos\[8\] _07994_ _07995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13136_ rbzero.texu_hot\[3\] _06949_ _06950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18993_ rbzero.tex_g0\[32\] rbzero.tex_g0\[31\] _11866_ _11870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14847__A1 _08315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23031__A1 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17944_ _08073_ rbzero.wall_tracer.rayAddendX\[8\] _11088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13067_ _06882_ _06883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_206_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19786__A1 _12422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17875_ _11008_ _11016_ _11018_ _11019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13336__I _07065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19614_ _12282_ _12386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16826_ _10255_ _10256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__22649__I _11399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14075__A2 _07884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23334__A2 _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19545_ rbzero.wall_tracer.visualWallDist\[-8\] _12198_ _12316_ _12317_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_45_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16757_ _10193_ _10188_ _10189_ _10195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_13969_ _07204_ _07720_ _07229_ _07779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__19023__I _11871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_175_i_clk_I clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15708_ _09349_ _09350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_158_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19476_ _12175_ _12248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16688_ _10066_ _10131_ _10024_ _10132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_152_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15639_ _09297_ _09298_ _09290_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18427_ _11520_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16772__A1 rbzero.debug_overlay.playerX\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18358_ rbzero.tex_g1\[1\] rbzero.tex_g1\[0\] _11481_ _11482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17309_ rbzero.pov.spi_buffer\[31\] _10637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16524__A1 _08105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18289_ rbzero.wall_tracer.mapX\[10\] _11406_ _11428_ _11429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_43_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20320_ _12486_ _12645_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19693__I _12464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20251_ _12280_ _13021_ _13022_ _13023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20182_ _12873_ _12925_ _12954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21820__A2 _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25011__A2 _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15726__I _09352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24990_ _05761_ _05771_ _05772_ _05773_ _05774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_235_Right_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23941_ _04721_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_209_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21584__A1 _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26660_ _00570_ clknet_leaf_158_i_clk rbzero.tex_b0\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23872_ rbzero.wall_tracer.rcp_fsm.o_data\[-7\] _04696_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_193_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_162_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input15_I i_gpout2_sel[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25611_ _06349_ _06393_ _06394_ _06395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_223_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22823_ _03667_ _02614_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26591_ _00501_ clknet_leaf_33_i_clk rbzero.pov.spi_buffer\[60\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25542_ _06277_ _06292_ _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22754_ _03586_ _02567_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_94_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21705_ _02765_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_25473_ _06219_ _06248_ _06256_ _06257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_109_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22685_ _03548_ _03552_ _03553_ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27212_ _01117_ clknet_leaf_76_i_clk rbzero.wall_tracer.stepDistY\[-3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24424_ _05087_ _05019_ _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_19_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21636_ rbzero.wall_tracer.rayAddendX\[-6\] _02689_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19701__A1 _12472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17388__I _10542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27143_ _00004_ clknet_leaf_73_i_clk rbzero.wall_tracer.rcp_fsm.state\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24355_ _05063_ _05064_ _05110_ _05111_ _05139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_180_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21567_ _02260_ _02403_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13849__C _07603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13329__A1 _06884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23306_ _03651_ _04159_ _04160_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20518_ _12283_ _01436_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27074_ _00984_ clknet_leaf_143_i_clk rbzero.tex_b1\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24286_ _05069_ _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_21498_ _02462_ _02494_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_169_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26025_ _06769_ _06799_ _06682_ _06785_ _06743_ _06800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_23237_ _04091_ _04092_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20449_ _01491_ _01542_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_28_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23168_ _04020_ _04021_ _04022_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_182_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14829__B2 _08502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_223_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22119_ _03110_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23099_ _03935_ _03955_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_15990_ _09550_ _09562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_147_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14941_ rbzero.vga_sync.vsync _08744_ _08745_ net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_26927_ _00837_ clknet_leaf_172_i_clk rbzero.tex_r1\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XFILLER_0_246_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_237_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_202_Right_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_17660_ _10866_ rbzero.pov.ready_buffer\[10\] _10871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26858_ _00768_ clknet_leaf_187_i_clk rbzero.tex_r0\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14872_ _07889_ _08659_ _08664_ _08669_ _08677_ _08678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_173_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16611_ _10044_ _10045_ _10043_ _10059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25809_ _06579_ _06586_ _06593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_215_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13823_ rbzero.tex_r0\[25\] _07633_ _07634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_203_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_201_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17591_ _10826_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_201_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26789_ _00699_ clknet_leaf_128_i_clk rbzero.tex_g1\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_67_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16542_ _09989_ _09994_ _09995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19330_ _12127_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_197_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13754_ rbzero.tex_r0\[45\] _07543_ _07565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19261_ _12072_ _12088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16473_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] _09912_
+ _09930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18682__I _11650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15557__A2 _09232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13685_ _07495_ _07496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__20550__A2 _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18212_ _11341_ _11335_ _11353_ _11355_ _11356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_80_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15424_ _09139_ _09140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22827__A1 _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19192_ _12035_ _12036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_14_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_234_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18143_ rbzero.wall_tracer.visualWallDist\[-2\] _11287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15355_ _09054_ _09089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16506__A1 _08106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14715__I _07613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14306_ rbzero.debug_overlay.vplaneY\[-1\] _08116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18074_ _11211_ _11215_ _11217_ _11218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_151_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15286_ _09037_ _09038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17025_ _10407_ _10421_ _10422_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_22_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14237_ _08046_ _08047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16930__I rbzero.debug_overlay.playerY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20066__A1 _12816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20066__B2 _12675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14168_ _06888_ _07141_ _07195_ _07977_ _07978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_111_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15546__I _09190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13119_ _06912_ _06931_ _06932_ _06933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_226_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14099_ _07523_ _07909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18976_ _11860_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_238_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17927_ _08072_ _11025_ _11059_ _11071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__21566__A1 _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_17858_ rbzero.debug_overlay.facingX\[-2\] _11001_ _11002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__14048__A2 _07857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16809_ _10238_ _10239_ _10240_ _10241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__16377__I _09819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25911__C _10992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17789_ _10951_ _10702_ _10954_ _10956_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_19528_ _12299_ _12300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_152_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21869__A2 _10466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19459_ _12202_ _12231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__16745__A1 _10168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22470_ _07983_ _03403_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_173_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14220__A2 _07995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21421_ _12780_ _01918_ _02388_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_146_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17545__I0 rbzero.tex_b0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24140_ _04719_ _04913_ _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_142_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21352_ _02325_ _02438_ _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19637__B _12408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20303_ _12982_ _13030_ _01397_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_141_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24071_ rbzero.wall_tracer.rcp_fsm.operand\[-2\] rbzero.wall_tracer.rcp_fsm.operand\[-3\]
+ _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_21283_ _02368_ _02369_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23022_ _03776_ _03879_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20234_ _12986_ _13005_ _13006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_203_Left_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__24418__S1 _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20165_ _12926_ _12936_ _12937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_164_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14287__A2 _08078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15484__A1 _06958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20096_ _12611_ _12655_ _12868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_24973_ _05635_ _05755_ _05756_ _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_129_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26712_ _00622_ clknet_leaf_30_i_clk rbzero.pov.ready_buffer\[42\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23924_ _04726_ _04729_ _10508_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22289__I _10048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14039__A2 _07845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26643_ _00553_ clknet_leaf_147_i_clk rbzero.tex_b0\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_98_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23855_ _04683_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13704__I _07340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22806_ _03659_ _03664_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_212_Left_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_26574_ _00484_ clknet_leaf_27_i_clk rbzero.pov.spi_buffer\[43\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23786_ _03612_ _04622_ _04623_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_179_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20998_ _12698_ _01967_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_179_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25525_ _06272_ _06083_ _06309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22737_ rbzero.wall_tracer.stepDistX\[0\] _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_138_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15539__A2 _09030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25456_ _05696_ _05822_ _06225_ _06240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_62_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13470_ _07279_ _07280_ _07281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24009__I _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22668_ _03538_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_216_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24407_ _05039_ _05054_ _05117_ _05191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_192_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15140__B _08887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21619_ _02694_ _02696_ _02698_ _10036_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_25387_ _06130_ _06132_ _06171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_129_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22599_ _07241_ _08752_ _03086_ _03484_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_36_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15140_ _08919_ _08921_ _08887_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27126_ _01036_ clknet_leaf_120_i_clk rbzero.traced_texVinit\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24338_ _04966_ _05122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15071_ _08809_ rbzero.spi_registers.ss_buffer\[1\] _08864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_27057_ _00967_ clknet_leaf_133_i_clk rbzero.tex_b1\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA_clkbuf_leaf_123_i_clk_I clknet_5_18__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_221_Left_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_24269_ _04720_ _04913_ _05052_ _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26008_ _06737_ _06785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14022_ _07831_ _07832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__17067__B _10436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20599__A2 _12587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18110__B1 _11251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18830_ _11752_ _11756_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22701__B _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18761_ rbzero.tex_r1\[47\] rbzero.tex_r1\[46\] _11708_ _11711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15973_ rbzero.spi_registers.buf_mapdx\[0\] _09548_ _09549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_235_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_199_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17712_ _10905_ _10906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14924_ _08215_ _08222_ _07472_ _08360_ _08730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__22199__I _10151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_199_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18692_ _11671_ _11672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_231_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14855_ rbzero.tex_b1\[9\] _08568_ _08289_ _08661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17643_ _10858_ _10554_ _10851_ _10860_ _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_19_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13806_ _07594_ _07617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_236_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17574_ _10816_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14786_ _08565_ _08589_ _08592_ _08593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_48_i_clk_I clknet_5_17__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14450__A2 _08258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16525_ _09914_ _09978_ _09979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_19313_ rbzero.tex_b1\[35\] rbzero.tex_b1\[34\] _12115_ _12118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13737_ rbzero.tex_r0\[37\] _07532_ _07548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16456_ _08100_ _09914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19244_ rbzero.tex_b1\[5\] rbzero.tex_b1\[4\] _12078_ _12079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13668_ _07417_ _07479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15407_ rbzero.spi_registers.buf_sky\[4\] _09119_ _09128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19175_ _11252_ _12007_ _12019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16387_ _09859_ _09860_ _09856_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13599_ _06867_ _07391_ _07409_ _06857_ _07410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__20891__B _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20287__A1 _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18126_ rbzero.debug_overlay.playerY\[0\] _11269_ _11270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_15338_ _08883_ _09077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17756__I _10847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18057_ rbzero.wall_tracer.trackDistX\[-8\] _11201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__23225__A1 _12949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15269_ rbzero.spi_registers.buf_otherx\[2\] _09021_ _09024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17008_ _10374_ _10410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15276__I _09028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21539__A1 _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18959_ _11850_ _11851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_225_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25922__B _05880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21970_ _03000_ _02998_ _03001_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer12 _05181_ net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer23 _04992_ net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_20921_ _01875_ _01876_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_5_15__f_i_clk_I clknet_3_3_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer34 _04862_ net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_1
XFILLER_0_179_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16966__A1 _08876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20762__A2 _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23640_ _04223_ _04054_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_124_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20852_ _01940_ _01941_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_76_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23700__A2 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23571_ _04410_ _04422_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20783_ _01683_ _01684_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25310_ _06072_ _06093_ _06094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_119_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22522_ _09972_ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26290_ _00200_ clknet_leaf_228_i_clk rbzero.spi_registers.buf_floor\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25241_ _06024_ _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22453_ _03385_ _03388_ _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17518__I0 rbzero.tex_b0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20278__A1 _12979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Left_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21404_ _02214_ _02488_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25172_ _05950_ _05953_ _05955_ _05956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__17143__A1 rbzero.pov.ready_buffer\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22384_ _01550_ _03329_ _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24123_ _04737_ _04906_ _04907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_103_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21335_ _02226_ _02229_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__17694__A2 rbzero.pov.ready_buffer\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24054_ _04781_ _04837_ _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__23767__A2 _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21266_ _02351_ _02352_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__21778__A1 _12216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15186__I _08916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23005_ _03861_ _03862_ _03738_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_20217_ _12480_ _12989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13180__A2 _06913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21197_ _02269_ _02284_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_229_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20148_ _12523_ _12919_ _12920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22578__I0 rbzero.wall_tracer.wall\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15914__I _09504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20079_ _12843_ _12848_ _12850_ _12851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_24956_ _05696_ _05739_ _05740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23907_ _04351_ _04696_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_231_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24887_ _05659_ _05669_ _05670_ _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16957__A1 _08066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21950__A1 _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14640_ _07513_ _08448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_26626_ _00536_ clknet_leaf_160_i_clk rbzero.tex_b0\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23838_ rbzero.wall_tracer.trackDistY\[8\] _03074_ _04664_ _04669_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_218_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14968__C2 _07179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_218_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_194_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14571_ rbzero.trace_state\[3\] _08379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
X_26557_ _00467_ clknet_leaf_67_i_clk rbzero.pov.spi_buffer\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23769_ _04605_ _04608_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_170_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__20505__A2 _12917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21702__A1 _08066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16310_ _09741_ _09802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25508_ _06280_ _06289_ _06291_ _06292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_13522_ _07332_ _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_60_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17290_ rbzero.pov.spi_buffer\[26\] _10623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26488_ _00398_ clknet_leaf_57_i_clk rbzero.debug_overlay.facingX\[-1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Left_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_231_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_231_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16241_ _08913_ _09748_ _09752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25439_ _06187_ _06182_ _06223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_97_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13453_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] _07264_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16681__S _10125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20269__A1 _13037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16172_ _09660_ _09700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13384_ _07189_ _07194_ _07195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__22482__I _09938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17134__A1 rbzero.pov.ready_buffer\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15123_ _08906_ _08907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_27109_ _01019_ clknet_leaf_142_i_clk rbzero.tex_b1\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_105_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18882__A1 rbzero.traced_texa\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19931_ _12687_ _12702_ _12695_ _12703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__23758__A2 _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15054_ rbzero.spi_registers.spi_counter\[3\] _08846_ _08847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__24403__S _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14005_ _07806_ _07809_ _07813_ _07814_ _07648_ _07815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_120_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_246_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19862_ _12549_ _12550_ _12634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__22430__A2 _07700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15448__A1 rbzero.spi_registers.vshift\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_118_Left_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_18813_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] _11742_ _11743_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_19793_ _12556_ _12564_ _12565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_37_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18744_ _11701_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15956_ _09534_ _09535_ _09536_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_223_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14907_ _08709_ _08710_ _08712_ _08558_ _08595_ _08713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_15887_ _09483_ _09484_ _09473_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16948__A1 _10295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18675_ _11662_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25132__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17626_ rbzero.pov.spi_done _10847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_106_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14838_ rbzero.tex_b1\[18\] _08528_ _08643_ _08644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_188_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14769_ rbzero.tex_b0\[19\] _08340_ _08576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17557_ _10801_ _10807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_127_Left_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16508_ _09927_ _09960_ _09962_ _09963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20177__I _12760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17488_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _10765_ _10768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19227_ rbzero.wall_tracer.mapY\[10\] _12067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_16439_ _09896_ _09897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19158_ _11915_ _11980_ _12001_ _12002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_143_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18109_ rbzero.debug_overlay.playerY\[1\] _11252_ _11253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19089_ _11927_ _11931_ _11932_ _11933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21120_ _02091_ _02207_ _01839_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__23749__A2 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_136_Left_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21051_ _02136_ _02139_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20002_ _12768_ _12772_ _12773_ _12774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_226_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20983__A2 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24810_ _05557_ _05593_ _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__19206__I _12044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25790_ _06553_ _06568_ _06574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14662__A2 _07940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24741_ _05468_ _05475_ _05479_ _05524_ _05525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_94_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21953_ _02988_ _02984_ _02989_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_193_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16939__A1 _08057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21932__A1 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21932__B2 _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20904_ _01993_ _11390_ _12583_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_29_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24672_ _05396_ _05404_ _05456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21884_ _08122_ _08143_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_178_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_145_Left_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_3_3_0_i_clk clknet_0_i_clk clknet_3_3_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_194_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26411_ _00321_ clknet_leaf_15_i_clk rbzero.spi_registers.buf_texadd3\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23623_ _04471_ _04472_ _04474_ _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_27391_ _01296_ clknet_leaf_107_i_clk rbzero.wall_tracer.stepDistX\[-11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20835_ _01804_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_194_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26342_ _00252_ clknet_leaf_11_i_clk rbzero.spi_registers.buf_texadd0\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23554_ _04402_ _04403_ _04406_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_119_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20766_ _01855_ _01856_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_42_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26886__CLKN clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22505_ _03425_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_213_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26273_ _00183_ clknet_leaf_17_i_clk rbzero.spi_registers.texadd3\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23485_ _04302_ _04338_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20697_ _01786_ _01787_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25224_ _05718_ _06007_ _06008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_220_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23988__A2 _08813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22436_ _03346_ _03378_ _03347_ _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_220_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20815__I _12950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17116__A1 _09933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25155_ _05878_ _05883_ _05939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22367_ rbzero.mapdyw\[1\] _12038_ _03314_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24106_ _04868_ _04889_ _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_231_i_clk clknet_5_0__leaf_i_clk clknet_leaf_231_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_92_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21318_ _02249_ _02404_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25086_ _05864_ _05870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22298_ _11177_ _03239_ _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24037_ _04775_ _04817_ _04819_ _04779_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_202_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21249_ _01954_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_229_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_246_i_clk clknet_5_0__leaf_i_clk clknet_leaf_246_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15810_ _09424_ _09425_ _09417_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_70_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16790_ rbzero.debug_overlay.playerX\[-2\] _10223_ _10224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_244_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25988_ _06752_ _06765_ _06766_ _06745_ _06767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_245_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14653__A2 _07807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15850__A1 _08942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15741_ _09352_ _09375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_198_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24939_ _05642_ _05722_ _05723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_99_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19592__A2 _12172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18460_ _11539_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15672_ rbzero.spi_registers.texadd2\[8\] _09315_ _09323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_197_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14623_ rbzero.tex_g1\[34\] _07890_ _08431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_17411_ rbzero.pov.spi_buffer\[57\] _10709_ _10706_ _10714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_200_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26609_ _00519_ clknet_leaf_168_i_clk rbzero.tex_b0\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_68_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18391_ rbzero.tex_g1\[16\] rbzero.tex_g1\[15\] _11496_ _11500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_201_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17342_ _10649_ _10662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14554_ _07467_ _08362_ _07474_ _08363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__23810__B _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13505_ _07261_ _07265_ _07315_ _07316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17273_ rbzero.pov.spi_buffer\[22\] _10610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14485_ _07819_ _08294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16224_ _09011_ _09732_ _09738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19012_ rbzero.tex_g0\[40\] rbzero.tex_g0\[39\] _11877_ _11881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13916__A1 rbzero.map_overlay.i_otherx\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13436_ _07244_ _07246_ _07247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17107__A1 rbzero.pov.ready_buffer\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer3 _05143_ net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_248_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16155_ _09675_ _09687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_248_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13367_ _07178_ _07179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__17658__A2 rbzero.pov.ready_buffer\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_248_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20662__A1 _12237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15106_ _08857_ _08892_ _08895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16086_ rbzero.spi_registers.buf_texadd0\[12\] _09633_ _09634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13298_ rbzero.spi_registers.texadd3\[4\] _07111_ _07035_ rbzero.spi_registers.texadd0\[4\]
+ _07112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_19914_ _12685_ _12686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15037_ _08825_ _08829_ _08830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_121_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__16881__A3 _08048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19845_ _12552_ _12565_ _12616_ _12617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__20460__I _09939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_235_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19776_ _12259_ _12548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16988_ _10377_ _10395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_147_Right_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18727_ _11691_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15939_ _09521_ _09523_ _09520_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18658_ rbzero.tex_r1\[2\] rbzero.tex_r1\[1\] _11651_ _11653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_121_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24459__A3 _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17609_ _10836_ _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_18589_ _11607_ _11613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13802__I _07586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20620_ _01704_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_171_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23720__B _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20551_ _01482_ _01485_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23270_ rbzero.wall_tracer.stepDistX\[7\] _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__19099__A1 rbzero.debug_overlay.facingY\[-1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20482_ _01518_ _01537_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22221_ _11297_ _03091_ _03125_ _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17649__A2 rbzero.pov.ready_buffer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__20653__A1 _12661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22152_ rbzero.wall_tracer.rcp_fsm.i_data\[-4\] _03126_ _03138_ _03139_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__22850__I _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19645__B _12255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13249__I _07062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21103_ _12413_ _01436_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26960_ _00870_ clknet_leaf_112_i_clk rbzero.texV\[-10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_22083_ rbzero.wall_tracer.rcp_fsm.o_data\[10\] rbzero.wall_tracer.stepDistY\[10\]
+ _03033_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25911_ _06903_ _02988_ _06661_ _06693_ _10992_ _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_21034_ _02117_ _02122_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13693__B _07493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26891_ _00801_ clknet_leaf_177_i_clk rbzero.tex_r0\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_25842_ _06625_ _06626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_35_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17821__A2 rbzero.pov.ready_buffer\[65\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14635__A2 _07906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25773_ _06520_ _06524_ _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_222_i_clk_I clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22985_ _12760_ _03842_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__18775__I _11713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20708__A2 _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_153_Left_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__19574__A2 _11993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24724_ _05503_ _05504_ _05507_ _05508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_21936_ _02972_ _02973_ _02974_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__21381__A2 _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27443_ _01348_ clknet_leaf_70_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24655_ _05306_ _05439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16295__I _09741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21867_ _02897_ _02896_ _02894_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_195_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13712__I _07340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23606_ _04359_ _04456_ _04457_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_139_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27374_ _01279_ clknet_leaf_89_i_clk rbzero.wall_tracer.trackDistY\[-6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20818_ _01905_ _01859_ _01868_ _01907_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_24586_ _05362_ _05365_ _05368_ _05369_ _05370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_148_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21798_ _10477_ _02845_ _02846_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_26325_ _00235_ clknet_leaf_234_i_clk rbzero.spi_registers.buf_mapdy\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23537_ _04384_ _04389_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20749_ rbzero.wall_tracer.size_full\[7\] _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__26072__A2 rbzero.wall_tracer.rcp_fsm.o_data\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15899__A1 _08942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14270_ _08079_ _08011_ _08080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26256_ _00166_ clknet_leaf_8_i_clk rbzero.spi_registers.texadd2\[23\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23468_ _04321_ _04217_ _04225_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_80_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_162_Left_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_59_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25207_ _05915_ _05990_ _05991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_190_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13221_ _07020_ _07035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_170_i_clk clknet_5_11__leaf_i_clk clknet_leaf_170_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_22419_ _08061_ _08176_ _03341_ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26187_ _00097_ clknet_leaf_241_i_clk rbzero.spi_registers.texadd0\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_189_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23399_ _04137_ _04139_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_25138_ _05840_ _05921_ _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13152_ rbzero.texu_hot\[0\] _06965_ _06966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_103_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25069_ _05845_ _05852_ _05853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13083_ _06897_ _06898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17960_ _11101_ _11104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_226_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_243_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14874__A2 _08298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_185_i_clk clknet_5_3__leaf_i_clk clknet_leaf_185_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16911_ _07705_ _08061_ _10316_ _10330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_17891_ _10996_ _11032_ _11034_ _11035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_217_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25335__A1 _05996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19630_ _12401_ _12402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16842_ rbzero.pov.ready_buffer\[72\] _10260_ _10269_ _10266_ _10264_ _10270_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__17812__A2 rbzero.pov.ready_buffer\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_171_Left_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_205_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15823__A1 rbzero.spi_registers.texadd3\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14626__A2 _07894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19561_ _12331_ _12332_ _12333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13985_ _07204_ _06865_ _07795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_16773_ _10167_ _10209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_204_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18512_ _11569_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_232_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15724_ _09349_ _09362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19492_ _12263_ _12264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_232_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18443_ rbzero.tex_g1\[38\] rbzero.tex_g1\[37\] _11528_ _11530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15655_ rbzero.spi_registers.buf_texadd2\[3\] _09306_ _09311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15051__A2 _08843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14606_ rbzero.tex_g1\[12\] _07821_ _08413_ _08414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_123_i_clk clknet_5_18__leaf_i_clk clknet_leaf_123_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15586_ rbzero.spi_registers.buf_texadd1\[9\] _09259_ _09260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18374_ _11490_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14537_ _07551_ _08346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17325_ _10542_ _10649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_166_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14468_ _08276_ _08277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17256_ _10596_ _10594_ _10597_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_181_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_138_i_clk clknet_5_15__leaf_i_clk clknet_leaf_138_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_16207_ _09724_ _09725_ _09723_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13419_ _07175_ _07229_ _07178_ _07230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_180_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14453__I _07333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17187_ _10541_ _10546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14399_ rbzero.tex_g0\[30\] _08207_ _08208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20635__A1 _12596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16138_ _08843_ _09669_ _09674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_216_Right_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_171_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24377__A2 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16069_ _09620_ _09621_ _09615_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__26700__CLK clknet_leaf_63_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14865__A2 _07633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19828_ _12573_ _12599_ _12600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_166_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19759_ _12524_ _12529_ _12531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22770_ _03627_ _03628_ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22560__A1 _11290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22560__B2 rbzero.traced_texa\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21721_ _02739_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_177_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17004__I _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24301__A2 _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24440_ _05118_ _05183_ _05224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_96_i_clk_I clknet_5_26__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21652_ _02692_ _07772_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20603_ _01693_ _01694_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24371_ _04947_ _05107_ _05108_ _05109_ _05155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_191_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21583_ _02258_ _02546_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26110_ _00020_ clknet_leaf_242_i_clk rbzero.spi_registers.spi_buffer\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20874__A1 _12789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23322_ _04063_ _04067_ _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20534_ _01572_ _01626_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_27090_ _01000_ clknet_leaf_152_i_clk rbzero.tex_b1\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_145_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26041_ _06777_ _06787_ _06813_ _06738_ _06814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_23253_ _04073_ _04108_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__14553__A1 _08360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19867__I0 _11067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20465_ _01458_ _01461_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22204_ _03162_ _03164_ _03179_ _03180_ rbzero.wall_tracer.rcp_fsm.i_data\[6\] _03181_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_23184_ _12428_ _02595_ _03660_ _04039_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_20396_ _01477_ _01489_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_242_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25565__A1 _06271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22135_ _03119_ _03124_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14856__A2 _08448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13659__A3 _07468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22066_ _03066_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26943_ _00853_ clknet_leaf_177_i_clk rbzero.tex_r1\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__23040__A2 _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21017_ _02060_ _02105_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_233_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26874_ _00784_ clknet_leaf_165_i_clk rbzero.tex_r0\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_50_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14608__A2 _07597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25825_ _06573_ _06589_ _06609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_226_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_221_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23879__A1 rbzero.wall_tracer.rcp_fsm.o_data\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_242_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25756_ _06488_ _06502_ _06540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13770_ rbzero.tex_r0\[2\] _07579_ _07580_ _07581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_22968_ _03824_ _03825_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_241_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40_i_clk clknet_5_16__leaf_i_clk clknet_leaf_40_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_168_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24707_ _05434_ _05451_ _05491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_21919_ _10113_ _02959_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_25687_ _06434_ _06463_ _06471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22899_ _03753_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15440_ rbzero.spi_registers.vshift\[1\] _09151_ _09152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27426_ _01331_ clknet_leaf_82_i_clk rbzero.wall_tracer.rcp_fsm.operand\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24638_ _05419_ _05303_ _05421_ _05351_ _05422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_139_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15371_ _09098_ _09099_ _09100_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27357_ _01262_ clknet_leaf_105_i_clk rbzero.wall_tracer.trackDistX\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24569_ _05246_ _05250_ _05244_ _05245_ _05353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_154_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_55_i_clk clknet_5_25__leaf_i_clk clknet_leaf_55_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__26045__A2 _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17110_ _09915_ _10487_ _10488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14322_ _08131_ _08132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18090_ _11149_ _11152_ _11154_ _11157_ _11234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_26308_ _00218_ clknet_leaf_236_i_clk rbzero.spi_registers.buf_othery\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_27288_ _01193_ clknet_leaf_210_i_clk gpout0.hpos\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_208_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17041_ rbzero.pov.ready_buffer\[28\] _10434_ _10435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14544__A1 _08346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13347__A2 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26239_ _00149_ clknet_leaf_14_i_clk rbzero.spi_registers.texadd2\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14253_ _08030_ _08054_ _08063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22606__A2 _11391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13204_ _07008_ _07016_ _07017_ _07018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_61_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14184_ _07987_ _07993_ _07211_ _07994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__18286__A2 _11420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17584__I _10758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13135_ _06910_ _06947_ _06948_ _06949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18992_ _11869_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_238_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14847__A2 _08652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17943_ _10997_ _11087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13066_ gpout0.hpos\[9\] _06882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__23031__A2 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_206_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16049__A1 _09518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_206_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17874_ rbzero.debug_overlay.facingX\[-6\] _11017_ _11018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_206_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_206_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19613_ _12299_ _12264_ _12385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16825_ _08805_ _10255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_45_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19544_ _11385_ _12316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_232_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16756_ _10170_ _10194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13968_ _07254_ _07198_ _07777_ _07778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22542__A1 rbzero.wall_tracer.visualWallDist\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_118_i_clk_I clknet_5_19__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15707_ _09204_ _09349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19475_ _12246_ _12247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16687_ _08116_ _10131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13899_ _07707_ _07706_ _07709_ _07060_ _07710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_88_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13352__I gpout0.vinf vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15024__A2 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18426_ rbzero.tex_g1\[31\] rbzero.tex_g1\[30\] _11517_ _11520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15638_ rbzero.spi_registers.buf_texadd1\[23\] _09293_ _09298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23098__A2 _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18357_ _11480_ _11481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15569_ _09244_ _09246_ _09242_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20856__A1 _12733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17308_ _10634_ _10630_ _10636_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18288_ _11426_ _11422_ _11427_ _11428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16524__A2 _08107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15279__I _09029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14535__A1 _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13338__A2 _07147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17239_ rbzero.pov.spi_buffer\[13\] _10585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_116_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20608__A1 _12206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19907__C _12369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20250_ rbzero.wall_tracer.stepDistX\[2\] _12316_ _13022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_9__f_i_clk clknet_3_2_0_i_clk clknet_5_9__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20181_ _12873_ _12925_ _12953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_228_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14838__A2 _08528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23940_ rbzero.wall_tracer.rcp_fsm.operand\[-6\] _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_32_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23871_ _04684_ _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_162_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25610_ _06336_ _06345_ _06394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_233_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22822_ _03668_ _02613_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__26608__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26590_ _00500_ clknet_leaf_33_i_clk rbzero.pov.spi_buffer\[59\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25541_ _06312_ _06323_ _06324_ _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22753_ _03612_ _03613_ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16212__A1 _09000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21704_ _11913_ _02764_ _02728_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_25472_ _06250_ _06254_ _06255_ _06256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_177_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22684_ _02737_ _01550_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_165_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_27211_ _01116_ clknet_leaf_80_i_clk rbzero.wall_tracer.stepDistY\[-4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_192_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24423_ _05206_ _05207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14774__A1 _07624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21635_ _08128_ rbzero.wall_tracer.rayAddendX\[-6\] _02711_ _02712_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_164_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27142_ _01052_ clknet_leaf_59_i_clk rbzero.wall_tracer.rayAddendY\[-6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24354_ _05136_ _05062_ _05105_ _05106_ _05137_ _05138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_133_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24038__A1 _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21566_ _02257_ _02250_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16515__A2 _09956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23305_ _04151_ _04159_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20517_ _01510_ _01511_ _01609_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27073_ _00983_ clknet_leaf_138_i_clk rbzero.tex_b1\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_127_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24285_ _04990_ _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_16_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21497_ _02519_ _02558_ _02581_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_169_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26024_ _06752_ _06765_ _06766_ _06720_ _06799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_31_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23236_ _03981_ _03989_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20448_ _01493_ _01541_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18268__A2 _11410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_4__f_i_clk_I clknet_3_1_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23167_ _04020_ _04021_ _04022_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_30_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20379_ _01471_ _01472_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22118_ _09897_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_246_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_223_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24210__A1 _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23098_ _03938_ _03954_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_246_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21024__A1 _12427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22049_ rbzero.wall_tracer.stepDistY\[-2\] _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14940_ _08744_ reg_vsync _08745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26926_ _00836_ clknet_leaf_129_i_clk rbzero.tex_r1\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__21654__I _10255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22772__A1 _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26857_ _00767_ clknet_leaf_187_i_clk rbzero.tex_r0\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14871_ _08315_ _08676_ _08677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_242_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16610_ _10057_ _10058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14696__C _08346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25808_ _06591_ _06588_ _06592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13822_ _07632_ _07633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_201_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17590_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _10823_ _10826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_67_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26788_ _00698_ clknet_leaf_128_i_clk rbzero.tex_g1\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_97_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16541_ _09990_ _09992_ _09993_ _09994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_13753_ rbzero.tex_r0\[46\] _07563_ _07489_ _07564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25739_ _05979_ _05988_ _06523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19260_ _12087_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_168_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16472_ _08109_ rbzero.wall_tracer.rayAddendY\[-5\] _09929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13684_ _07444_ _07495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_214_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__17951__A1 _11039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18211_ _11263_ _11308_ _11354_ _11109_ _11355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_27409_ _01314_ clknet_leaf_107_i_clk rbzero.wall_tracer.stepDistX\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13568__A2 _06873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15423_ _06898_ _09139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_183_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19191_ _11137_ _12035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__16483__I _09939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14765__B2 _08284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22827__A2 _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18142_ rbzero.wall_tracer.visualWallDist\[-1\] _11286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15354_ rbzero.spi_registers.buf_mapdxw\[1\] _09078_ _09088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14305_ _08103_ _08010_ _08016_ _08104_ _08114_ _08115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_18073_ _11205_ _11216_ _11217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15285_ _09028_ _09037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_124_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17024_ rbzero.pov.ready_buffer\[24\] _10403_ _10422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14236_ _08005_ _08034_ _08046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_111_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14167_ _06860_ _06870_ _07977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_44_i_clk_I clknet_5_16__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13118_ rbzero.spi_registers.texadd0\[12\] _06912_ _06932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14098_ rbzero.tex_r1\[41\] _07906_ _07907_ _07908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18975_ rbzero.tex_g0\[24\] rbzero.tex_g0\[23\] _11856_ _11860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_225_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17926_ _08079_ _11069_ _11027_ _11070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_56_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13049_ gpout0.hpos\[7\] _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19462__C _11390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13791__B _07601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17857_ rbzero.wall_tracer.rayAddendX\[6\] _11001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15245__A2 _08917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16808_ _08171_ _10232_ _10240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17788_ _10952_ rbzero.pov.ready_buffer\[53\] _10956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_221_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19527_ _12298_ _12299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_178_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16739_ _10178_ _10179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_220_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19458_ rbzero.wall_tracer.visualWallDist\[-2\] _12229_ _12230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18409_ _11510_ _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16393__I _09818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19389_ _12160_ _12161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21420_ _02500_ _02503_ _02505_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_29_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21351_ _02436_ _02437_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20302_ _12984_ _13029_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24070_ _04757_ _04853_ _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15181__A1 _08955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21282_ _02332_ _02334_ _02367_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_31_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24440__A1 _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23243__A2 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21254__A1 _12439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23021_ _03835_ _03878_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15737__I _09336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20233_ _12997_ _13004_ _13005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20164_ _12927_ _12935_ _12936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_164_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_129_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20095_ _12665_ _12669_ _12867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_228_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24972_ _05545_ _05597_ _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_157_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26711_ _00621_ clknet_leaf_30_i_clk rbzero.pov.ready_buffer\[41\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_243_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23923_ rbzero.wall_tracer.rcp_fsm.i_data\[-10\] _04728_ _04729_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15472__I _09111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23854_ _09896_ _02981_ _03085_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_26642_ _00552_ clknet_leaf_147_i_clk rbzero.tex_b0\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_98_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22506__A1 rbzero.wall_tracer.size\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22805_ _02600_ _03663_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_200_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14088__I _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23785_ _04620_ _04621_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26573_ _00483_ clknet_leaf_27_i_clk rbzero.pov.spi_buffer\[42\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20997_ _01946_ _01959_ _01955_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_223_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_179_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25524_ _06144_ _06147_ _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22736_ _03598_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25455_ _06183_ _06237_ _06238_ _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_149_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22667_ _03537_ _11205_ _11400_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_62_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13720__I _07482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_216_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24406_ _05099_ _05157_ _05185_ net55 _05189_ _05190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_11_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21618_ _02697_ _02694_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25386_ _06161_ _06164_ _06169_ _06170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_192_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22598_ _07236_ _11394_ _03483_ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_164_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24337_ _04905_ _05121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27125_ _01035_ clknet_leaf_120_i_clk rbzero.traced_texVinit\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_21549_ _12728_ _02633_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15070_ _08856_ _08862_ _08863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27056_ _00966_ clknet_leaf_133_i_clk rbzero.tex_b1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_132_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24268_ _04966_ _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_160_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26007_ _06694_ _03000_ _06776_ _06784_ _06719_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_205_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14021_ _07508_ _07831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15647__I _09257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19989__A2 _12760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23219_ _03978_ _03990_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__18023__I rbzero.wall_tracer.trackDistY\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13722__A2 _07532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24199_ _04923_ _04882_ _04885_ _04983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_120_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__18110__B2 rbzero.debug_overlay.playerY\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18760_ _11710_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15972_ _09547_ _09548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22745__A1 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17711_ _10843_ _10905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_199_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14923_ _07433_ _07446_ _08729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26909_ _00819_ clknet_leaf_126_i_clk rbzero.tex_r1\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_199_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18691_ _11649_ _11671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_188_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17642_ _10859_ rbzero.pov.ready_buffer\[3\] _10860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_215_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14854_ rbzero.tex_b1\[8\] _08258_ _08660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_215_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_203_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13805_ rbzero.tex_r0\[15\] _07592_ _07616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_236_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17573_ rbzero.tex_b0\[44\] rbzero.tex_b0\[43\] _10812_ _10816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14785_ _07912_ _08590_ _08591_ _08592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__18177__A1 rbzero.map_overlay.i_othery\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19312_ _12117_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16524_ _08105_ _08107_ rbzero.debug_overlay.vplaneY\[-8\] _09978_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_13736_ rbzero.tex_r0\[38\] _07545_ _07546_ _07547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_168_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19243_ _12072_ _12078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16455_ _09902_ rbzero.wall_tracer.rayAddendY\[-5\] _09912_ _09913_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14738__B2 _08284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13667_ _07348_ _07478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_128_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15406_ rbzero.color_sky\[4\] _09115_ _09127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19174_ _11354_ _12008_ _12018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16386_ rbzero.spi_registers.spi_buffer\[14\] _09853_ _09860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13598_ rbzero.row_render.size\[8\] _07389_ _07409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_137_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17527__I1 rbzero.tex_b0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18125_ rbzero.map_rom.d6 _11269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_206_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15337_ _07751_ _09075_ _09076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_27__f_i_clk clknet_3_6_0_i_clk clknet_5_27__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_18056_ _11195_ _11196_ _11198_ _11199_ _11200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__15163__A1 _08939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_1 _07804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15268_ rbzero.map_overlay.i_otherx\[2\] _09019_ _09023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17007_ _10407_ _10408_ _10409_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14219_ _08028_ _08029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_22_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15199_ _08933_ _08971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18958_ _11828_ _11850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17909_ _11046_ _11051_ _11052_ _11053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18889_ _11769_ _11804_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_241_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_20920_ _02008_ _01880_ _02009_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xrebuffer13 _06160_ net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer24 _04979_ net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer35 _05207_ net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__20762__A3 _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20851_ _12429_ _01712_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_124_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18168__A1 rbzero.map_overlay.i_mapdy\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23570_ _04410_ _04422_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_20782_ _01871_ _01872_ _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_147_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21711__A2 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22521_ _03434_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__25989__A1 _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25240_ _05466_ _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_162_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22452_ _03383_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__19668__A1 rbzero.wall_tracer.visualWallDist\[-3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21403_ _02488_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25171_ _05918_ _05927_ _05954_ _05955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13952__A2 rbzero.map_overlay.i_mapdy\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22383_ _03327_ _08042_ _03328_ _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17143__A2 _10485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24122_ _04819_ _04869_ _04906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21334_ _02279_ _02280_ _02420_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_40_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24053_ _04831_ _04830_ _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21265_ _12790_ _01971_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23004_ _03727_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21778__A2 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20216_ _12274_ _12988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_21196_ _02273_ _02283_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20147_ _12918_ _12919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_239_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_217_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22727__A1 _11134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22578__I1 _08364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20078_ _12811_ _12849_ _12850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24955_ _05729_ _05738_ _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13715__I _07331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23906_ _03024_ _04711_ _04715_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__24319__I2 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24886_ _05666_ _05668_ _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_170_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26625_ _00535_ clknet_leaf_160_i_clk rbzero.tex_b0\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__14968__A1 _07180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23837_ _03296_ _03074_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_218_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_194_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14570_ _08378_ net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23768_ _04606_ _04601_ _04607_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20548__I _12527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26556_ _00466_ clknet_leaf_67_i_clk rbzero.pov.spi_buffer\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17906__A1 _08084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25507_ _06133_ _06134_ _06290_ _06151_ _06158_ _06291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_13521_ _07331_ _07332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_211_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22719_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] _03578_
+ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14546__I _07349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23699_ rbzero.wall_tracer.trackDistY\[-9\] _03037_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26487_ _00397_ clknet_leaf_57_i_clk rbzero.debug_overlay.facingX\[-2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_231_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16240_ rbzero.spi_registers.buf_texadd2\[1\] _09743_ _09751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13452_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] _07263_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_231_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25438_ _06184_ _06102_ _06222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_97_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24652__A1 _05275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24652__B2 _05257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25369_ _05720_ _06012_ _06153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13383_ _07193_ _07194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16171_ _08948_ _09698_ _09699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15122_ _08905_ _08906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_217_i_clk_I clknet_5_3__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27108_ _01018_ clknet_leaf_142_i_clk rbzero.tex_b1\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_90_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24404__A1 _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18882__A2 rbzero.texV\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19930_ _12695_ _12701_ _12702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15053_ _08835_ _08840_ _08845_ _08846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_27039_ _00949_ clknet_leaf_158_i_clk rbzero.tex_g0\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XFILLER_0_32_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23808__B _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14004_ _07501_ _07814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19861_ _12588_ _12598_ _12589_ _12633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_246_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18812_ _11735_ _11740_ _11741_ _11742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15448__A2 _09151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19792_ _12558_ _12559_ _12563_ _12564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_208_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18743_ rbzero.tex_r1\[39\] rbzero.tex_r1\[38\] _11698_ _11701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__25380__A2 _06129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15955_ _09504_ _09536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14906_ rbzero.tex_b1\[52\] _08698_ _08711_ _08712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_216_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18674_ rbzero.tex_r1\[9\] rbzero.tex_r1\[8\] _11661_ _11662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15886_ _08920_ _09477_ _09484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14959__A1 _07074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17625_ _10228_ _10846_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__25132__A2 _05321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14837_ rbzero.tex_b1\[19\] _08529_ _08643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14959__B2 _07153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17556_ _10806_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__19898__A1 _12665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14768_ _08339_ _08573_ _08574_ _08575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13631__A1 _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23694__A2 rbzero.wall_tracer.stepDistY\[-10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16507_ _09945_ _09961_ _09962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13719_ _07480_ _07506_ _07529_ _07530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_184_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17487_ _10767_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14699_ _07566_ _08506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19226_ _12061_ _12049_ _12050_ _12066_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_16438_ _09895_ _09896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_27_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19157_ _08149_ rbzero.wall_tracer.rayAddendY\[9\] _12001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_143_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16369_ rbzero.spi_registers.buf_texadd3\[10\] _09840_ _09847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18108_ rbzero.map_rom.c6 _11252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_19088_ _08156_ _10007_ _11932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21209__A1 _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16884__A1 _10293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18039_ _11176_ _11180_ _11182_ _11183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14344__C1 _08022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21050_ _02137_ _02138_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20001_ _12769_ _12771_ _12773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_238_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_240_Left_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__22709__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25371__A2 _05998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14111__A2 _07920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21952_ rbzero.wall_tracer.size_full\[-10\] _02986_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24740_ _05473_ _05474_ _05469_ _05471_ _05524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_2_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20903_ rbzero.wall_tracer.stepDistX\[-1\] _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_24671_ _05396_ _05404_ _05455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_29_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21883_ _02910_ _02911_ _02915_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_23622_ _04397_ _04400_ _04473_ _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_26410_ _00320_ clknet_leaf_13_i_clk rbzero.spi_registers.buf_texadd3\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_159_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20834_ _01682_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_166_i_clk_I clknet_5_8__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27390_ _01295_ clknet_leaf_95_i_clk rbzero.wall_tracer.trackDistY\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20499__A2 _12518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23553_ _04404_ _04405_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26341_ _00251_ clknet_leaf_237_i_clk rbzero.spi_registers.buf_texadd0\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__21696__A1 _07693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20765_ _01755_ _01764_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14366__I rbzero.debug_overlay.playerX\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23679__I _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22504_ rbzero.wall_tracer.size\[8\] _03423_ _03424_ _07354_ _03425_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26272_ _00182_ clknet_leaf_17_i_clk rbzero.spi_registers.texadd3\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_213_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23484_ _04305_ _04307_ _04337_ _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_18_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20696_ _01673_ _01769_ _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25223_ _06006_ _06007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22435_ _03374_ _03377_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_137_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19361__I0 rbzero.tex_b1\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25154_ _05885_ _05902_ _05937_ _05938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_22366_ _11330_ _11367_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24105_ _04753_ _04870_ _04889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__15197__I _08951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21317_ _02403_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_92_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16875__A1 _10293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24937__A2 _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25085_ _05824_ _05866_ _05868_ _05869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__20671__A2 _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22297_ _03253_ _03256_ _03258_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_229_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24036_ _04819_ _04817_ _04775_ _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_57_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21248_ _02196_ _02201_ _02194_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24303__I _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__20423__A2 _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14969__C _08747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21179_ _02156_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25987_ _06703_ _06724_ _06766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_217_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13310__B1 _07109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15740_ rbzero.spi_registers.texadd3\[1\] _09373_ _09374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24938_ _05687_ _05719_ _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22758__I _11409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21662__I _12044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15671_ _09321_ _09322_ _09314_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_24869_ _05328_ _05413_ _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_213_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17410_ _10712_ _10713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_29_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26608_ _00518_ clknet_leaf_168_i_clk rbzero.tex_b0\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14622_ _08405_ _08429_ _07928_ _08430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_201_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18390_ _11499_ _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_185_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17341_ rbzero.pov.spi_buffer\[39\] _10661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14553_ _08360_ _07472_ _08361_ _08362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26539_ _00449_ clknet_leaf_23_i_clk rbzero.pov.spi_buffer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13504_ _07266_ _07271_ _07314_ _07315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22493__I _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17272_ _10608_ _10606_ _10609_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_181_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24625__A1 _05296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14484_ rbzero.tex_g0\[35\] _08288_ _08292_ _08293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19011_ _11880_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_180_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__21439__A1 _12238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16223_ rbzero.spi_registers.buf_texadd1\[22\] _09730_ _09737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13435_ _07201_ _07245_ _07246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_64_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__17107__A2 _10485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer4 net58 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_248_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13366_ gpout0.vpos\[9\] _07178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16154_ rbzero.spi_registers.buf_texadd1\[4\] _09685_ _09686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_248_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_248_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15105_ _08864_ _08894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__20662__A2 _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16085_ _09596_ _09633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13297_ _06928_ _07111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_19913_ _12304_ _12685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15036_ _08826_ _08828_ _08829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_239_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19844_ _12556_ _12564_ _12616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19775_ _12487_ _12527_ _12547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16987_ _08087_ _10393_ _10394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_218_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13355__I _07166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13301__B1 _07026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18726_ rbzero.tex_r1\[32\] rbzero.tex_r1\[31\] _11687_ _11691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15938_ _09522_ _09507_ _09523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13852__A1 _07624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21914__A2 _10474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18657_ _11652_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15869_ _09462_ _09469_ _09470_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_121_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23116__A1 _12949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19042__I _11892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25979__I _10255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24459__A4 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17608_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _10833_ _10836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18588_ _11612_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17539_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _10796_ _10797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22617__B _09927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20550_ _12235_ _01642_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19209_ rbzero.wall_tracer.mapY\[6\] _12009_ _12034_ _12052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__13907__A2 rbzero.map_overlay.i_othery\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20481_ _01520_ _01573_ _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20137__B _12172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22220_ _09989_ _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14580__A2 _07818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22151_ _11989_ _03134_ _03137_ _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__20653__A2 _12448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22352__B _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21102_ _12483_ _13025_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__25219__I _05388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22082_ _03026_ _03034_ _03077_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__20651__I _12590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25592__A2 _06329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_92_i_clk_I clknet_5_24__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25910_ _06662_ _06682_ _06692_ _05007_ _06693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_21033_ _02118_ _02119_ _02121_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__13540__B1 _07349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26890_ _00800_ clknet_leaf_176_i_clk rbzero.tex_r0\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_22_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25841_ _06618_ _06601_ _06625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_226_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25772_ _06555_ _06556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_22984_ _02075_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24723_ _05505_ _05506_ _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_21935_ _02951_ _02963_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23107__A1 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21381__A3 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25889__I _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27442_ _01347_ clknet_leaf_70_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_195_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24654_ _05327_ _05437_ _05438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_167_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21866_ _02895_ _02898_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_26_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19887__I _12658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23605_ _04361_ _04455_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20817_ _01906_ _01867_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14096__I _07498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21669__A1 _08018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27373_ _01278_ clknet_leaf_98_i_clk rbzero.wall_tracer.trackDistY\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_139_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24585_ _05357_ _05349_ _05355_ _05369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_21797_ rbzero.debug_overlay.vplaneX\[-1\] _11080_ _02833_ _02846_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_154_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26324_ _00234_ clknet_leaf_234_i_clk rbzero.spi_registers.buf_mapdy\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20748_ _01526_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23536_ _04385_ _04388_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23202__I _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23467_ _03862_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26255_ _00165_ clknet_leaf_9_i_clk rbzero.spi_registers.texadd2\[22\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20679_ _01668_ _01770_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14020__A1 rbzero.tex_r1\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13220_ _07024_ _07032_ _07034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17200__I _10555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25206_ _05985_ _05990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_59_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22418_ _03360_ _03362_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23398_ _04133_ _04240_ _04251_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_26186_ _00096_ clknet_leaf_235_i_clk rbzero.spi_registers.texadd0\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23830__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13151_ _06962_ _06953_ _06963_ _06964_ _06965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_25137_ _05301_ _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_22349_ _03210_ _03298_ _03300_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__19555__C _12159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25068_ _05846_ _05851_ _05852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_72_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13082_ _06896_ _06897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_237_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_226_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_243_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24019_ _04749_ rbzero.wall_tracer.rcp_fsm.operand\[-5\] rbzero.wall_tracer.rcp_fsm.operand\[-6\]
+ rbzero.wall_tracer.rcp_fsm.operand\[-7\] _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA__23594__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16910_ _10327_ _10329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_17890_ _08075_ _11033_ _11034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_208_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16841_ _08184_ _07687_ _10250_ _10269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_205_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15823__A2 _09032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19560_ rbzero.wall_tracer.stepDistY\[-7\] _12271_ _11384_ _12332_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_16772_ rbzero.debug_overlay.playerX\[-4\] _10203_ _10208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_13984_ _07227_ _07078_ _07794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_18511_ rbzero.tex_r0\[3\] rbzero.tex_r0\[2\] _11566_ _11569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_232_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15723_ _09359_ _09360_ _09361_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19491_ _12262_ _12263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16486__I _08107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15390__I _09064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18442_ _11529_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15654_ rbzero.spi_registers.texadd2\[3\] _09303_ _09310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14605_ rbzero.tex_g1\[13\] _07811_ _08413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_18373_ rbzero.tex_g1\[8\] rbzero.tex_g1\[7\] _11486_ _11490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15585_ _09258_ _09259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17324_ rbzero.pov.spi_buffer\[35\] _10648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14536_ _08334_ _08338_ _08344_ _08345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20883__A2 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17255_ rbzero.pov.spi_buffer\[18\] _10591_ _10588_ _10597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14734__I _07566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14467_ _07486_ _08276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_154_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16206_ _08994_ _09721_ _09725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13418_ _07228_ _07229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_17186_ _10544_ _10545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__23821__A2 _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14398_ _08206_ _08207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_180_Right_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16137_ rbzero.spi_registers.buf_texadd1\[0\] _09672_ _09673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__21832__A1 _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_114_i_clk_I clknet_5_31__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13349_ _07157_ net12 _07161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14314__A2 _08078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16068_ _08950_ _09612_ _09621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_227_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15019_ _08807_ net20 _08816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__20399__A1 _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19827_ _12588_ _12598_ _12599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_235_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13085__I _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24385__I0 _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_208_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19758_ _12524_ _12529_ _12530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_223_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18709_ _11681_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19689_ _12458_ _12459_ _12460_ _12461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_189_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13813__I _07608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21720_ _11113_ _11115_ _11117_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_182_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_230_i_clk clknet_5_2__leaf_i_clk clknet_leaf_230_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_177_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_39_i_clk_I clknet_5_16__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21651_ _02708_ _02721_ _02723_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18367__I1 rbzero.tex_g1\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20602_ _12987_ _12585_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24370_ _05066_ _05068_ _05070_ _04942_ _05154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_21582_ _02530_ _12959_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23321_ _04172_ _04175_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_20533_ _01582_ _01625_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20874__A2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_245_i_clk clknet_5_0__leaf_i_clk clknet_leaf_245_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_144_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26040_ _06811_ _06812_ _06813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22076__A1 _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23252_ _04076_ _04107_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_134_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20464_ _01544_ _01548_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23812__A2 _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22203_ _03108_ _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21823__A1 _10471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23183_ _03669_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20395_ _01488_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_101_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_242_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22134_ rbzero.wall_tracer.rcp_fsm.i_data\[-7\] _03088_ _03123_ _03124_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14305__A2 _08010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25565__A2 _06348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22065_ rbzero.wall_tracer.rcp_fsm.o_data\[4\] _03065_ _03033_ _03066_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_184_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26942_ _00852_ clknet_leaf_186_i_clk rbzero.tex_r1\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_184_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21016_ _02084_ _02104_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_215_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26873_ _00783_ clknet_leaf_165_i_clk rbzero.tex_r0\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_226_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23328__B2 _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25824_ _06549_ _06570_ _06608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_226_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_221_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25755_ _06484_ _06503_ _06539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22101__I _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22967_ _02504_ _02114_ _02633_ _01383_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13723__I _07418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24706_ _05345_ _05488_ _05489_ _05490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_69_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21918_ _02955_ _02939_ _02957_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_25686_ _06428_ _06462_ _06470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_195_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22898_ _02571_ _02687_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_210_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27425_ _01330_ clknet_leaf_83_i_clk rbzero.wall_tracer.rcp_fsm.operand\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_242_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24637_ _05371_ _05420_ _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21849_ _08138_ _08132_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_195_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27356_ _01261_ clknet_leaf_105_i_clk rbzero.wall_tracer.trackDistX\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15370_ _09054_ _09100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__21511__B1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24568_ _05205_ _05352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_182_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26307_ _00217_ clknet_leaf_235_i_clk rbzero.spi_registers.buf_othery\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14321_ rbzero.debug_overlay.vplaneX\[-5\] _08131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23519_ _04368_ _04370_ _04371_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_135_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27287_ _01192_ clknet_leaf_212_i_clk gpout0.hpos\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24499_ _05282_ _05283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23867__I _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17040_ _10378_ _10434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26238_ _00148_ clknet_leaf_14_i_clk rbzero.spi_registers.texadd2\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14252_ rbzero.debug_overlay.playerY\[-5\] _08062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_208_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13203_ rbzero.spi_registers.texadd0\[20\] _07008_ _07017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26169_ _00079_ clknet_leaf_227_i_clk rbzero.color_sky\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14183_ _07992_ _07990_ _07993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13134_ rbzero.spi_registers.texadd0\[9\] _06910_ _06948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18991_ rbzero.tex_g0\[31\] rbzero.tex_g0\[30\] _11866_ _11869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15385__I _08986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17942_ _11041_ _11067_ _11068_ _11085_ _11086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_13065_ _06860_ _06881_ net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__23816__B _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23031__A3 _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_206_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17873_ rbzero.wall_tracer.rayAddendX\[2\] _11017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17797__A2 rbzero.pov.ready_buffer\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_233_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19612_ _12383_ _12304_ _12384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16824_ rbzero.pov.ready_buffer\[70\] _10183_ _10212_ _10253_ _10254_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_21_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_19543_ _12314_ _12315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_233_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16755_ rbzero.debug_overlay.playerX\[-6\] _10193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_13967_ _07197_ _07078_ _07777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_85_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15706_ _09346_ _09347_ _09348_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_186_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19474_ _12179_ _12246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16686_ _10127_ _10128_ _10129_ _10130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_158_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13898_ _07708_ _07709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_40_i_clk_I clknet_5_16__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18425_ _11519_ _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15637_ rbzero.spi_registers.texadd1\[23\] _09291_ _09297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18356_ _11479_ _11480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_185_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14783__A2 _08300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15568_ rbzero.spi_registers.buf_texadd1\[5\] _09245_ _09246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15980__A1 _08968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17307_ rbzero.pov.spi_buffer\[31\] _10627_ _10635_ _10636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__20856__A2 _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14519_ _08316_ _08326_ _08327_ _08328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_151_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18287_ _11419_ _11406_ _11427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15499_ rbzero.spi_registers.buf_texadd0\[11\] _09194_ _09195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16524__A3 rbzero.debug_overlay.vplaneY\[-8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17238_ _10582_ _10583_ _10584_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_116_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20608__A2 _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22614__C _10049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17169_ _10512_ _10530_ _10531_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_101_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25992__I _05212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_20180_ _12948_ _12951_ _12952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_161_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_209_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17788__A2 rbzero.pov.ready_buffer\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23870_ _02994_ _04690_ _04695_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_162_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_22821_ _03677_ _03678_ _03679_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_193_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25540_ _06269_ _06169_ _06306_ _06324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_22752_ _03607_ _03610_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_177_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_190_Left_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_177_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21703_ _02761_ _02762_ _02763_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_25471_ _06063_ _06094_ _06104_ _06255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_22683_ _11238_ _12499_ _03551_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__16854__I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27210_ _01115_ clknet_leaf_76_i_clk rbzero.wall_tracer.stepDistY\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24422_ _05129_ _05182_ _05196_ _05205_ _05206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_21634_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] _02710_
+ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_184_i_clk clknet_5_2__leaf_i_clk clknet_leaf_184_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27141_ _01051_ clknet_leaf_44_i_clk rbzero.wall_tracer.rayAddendY\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24353_ _04896_ _05066_ _05068_ _05070_ _05137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_21565_ _12211_ _02524_ _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14374__I rbzero.debug_overlay.playerX\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23304_ _04150_ _04157_ _04158_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_20516_ _12706_ _01608_ _01512_ _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24284_ _05067_ _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_27072_ _00982_ clknet_leaf_138_i_clk rbzero.tex_b1\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_34_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21496_ _02460_ _02518_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_105_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26023_ _06903_ _03004_ _10988_ _06798_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_23235_ _03983_ _03988_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20447_ _01496_ _01540_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_199_i_clk clknet_5_12__leaf_i_clk clknet_leaf_199_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23166_ _03966_ _03971_ _03973_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_20378_ _01467_ _01470_ _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_246_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22117_ _03108_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_246_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_223_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23097_ _03943_ _03953_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__24210__A2 _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_122_i_clk clknet_5_13__leaf_i_clk clknet_leaf_122_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_22048_ _03004_ _03045_ _03055_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__22221__A1 _11297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21024__A2 _12433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26925_ _00835_ clknet_leaf_129_i_clk rbzero.tex_r1\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_238_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__17779__A2 rbzero.pov.ready_buffer\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26856_ _00766_ clknet_leaf_187_i_clk rbzero.tex_r0\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14870_ _08295_ _08672_ _08675_ _08676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_203_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25807_ _06576_ _06591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13821_ _07582_ _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_187_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_137_i_clk clknet_5_15__leaf_i_clk clknet_leaf_137_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26787_ _00697_ clknet_leaf_128_i_clk rbzero.tex_g1\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23999_ _04787_ _04776_ _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_203_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_201_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23721__A1 _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16540_ rbzero.debug_overlay.vplaneY\[-1\] _09965_ _09970_ _09993_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_67_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25738_ _05986_ _06521_ _06522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13752_ _07534_ _07563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_238_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16471_ _08112_ _09928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25669_ _06407_ _06452_ _06453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13683_ rbzero.tex_r0\[48\] _07487_ _07493_ _07494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_183_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18210_ _11256_ _11354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_27408_ _01313_ clknet_leaf_113_i_clk rbzero.wall_tracer.stepDistX\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22288__A1 _11288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15422_ _08197_ _09124_ _09138_ _09126_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_39_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19190_ _12031_ _12032_ _12034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_167_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19153__A1 _11986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18141_ _11281_ _11282_ _11283_ _11284_ _11285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_182_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15353_ rbzero.mapdxw\[1\] _09075_ _09087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_27339_ _01244_ clknet_leaf_37_i_clk rbzero.texu_hot\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17703__A2 rbzero.pov.ready_buffer\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18900__A1 rbzero.traced_texa\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14304_ _07719_ _08108_ _08113_ _08114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_18072_ _11207_ _11216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14517__A2 _07617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15284_ _09027_ _09031_ _09033_ _09036_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_123_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23788__A1 _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17023_ _08156_ _10401_ _10421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14235_ _08044_ _08045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_180_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22460__A1 _07150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14166_ _06878_ _07975_ _07976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_81_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13117_ rbzero.spi_registers.texadd3\[12\] _06921_ _06925_ rbzero.spi_registers.texadd2\[12\]
+ _06917_ rbzero.spi_registers.texadd1\[12\] _06931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__16004__I _09547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14097_ _07492_ _07907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18974_ _11859_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22450__B _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22212__A1 _11279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24221__I _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17925_ rbzero.wall_tracer.rayAddendX\[6\] _11069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13048_ _06864_ _06865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_218_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17856_ _10998_ _10999_ _11000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_206_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16807_ rbzero.debug_overlay.playerX\[0\] _10232_ _10239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_17787_ _10951_ _10699_ _10954_ _10955_ _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_221_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14999_ net86 _08797_ _08800_ _08801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__23712__A1 _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19526_ _12297_ _12298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16738_ net16 _10177_ _08882_ _10178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_241_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19457_ _12228_ _12229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16669_ _10109_ _10111_ _10113_ _10114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_220_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0_0_i_clk_I clknet_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17942__A2 _11067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18408_ rbzero.tex_g1\[23\] rbzero.tex_g1\[22\] _11507_ _11510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__20196__I _12553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19388_ _12159_ _12160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18339_ _07176_ _11466_ _11464_ _11468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_115_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21350_ _02327_ _02435_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23779__A1 _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20301_ _01375_ _01395_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21281_ _02332_ _02334_ _02367_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15181__A2 _08940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24440__A2 _05183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23020_ _03838_ _03877_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_229_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20232_ _13002_ _13003_ _13004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_228_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13538__I _07348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20163_ _12932_ _12934_ _12935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_164_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20094_ _12775_ _12864_ _12865_ _12866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_24971_ _05684_ _05753_ _05754_ _05755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_129_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13495__A2 _07305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_54_i_clk clknet_5_25__leaf_i_clk clknet_leaf_54_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_146_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22754__A2 _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26710_ _00620_ clknet_leaf_30_i_clk rbzero.pov.ready_buffer\[40\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23922_ _04727_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input20_I i_reg_mosi vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16433__A2 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26641_ _00551_ clknet_leaf_146_i_clk rbzero.tex_b0\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_93_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23853_ _04682_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_240_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22804_ _03661_ _03662_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_49_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22586__I _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26572_ _00482_ clknet_leaf_27_i_clk rbzero.pov.spi_buffer\[41\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20996_ _01974_ _01983_ _01968_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_23784_ _04620_ _04621_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_69_i_clk clknet_5_29__leaf_i_clk clknet_leaf_69_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_179_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25523_ _06161_ _06164_ _06307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_179_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22735_ _03597_ rbzero.wall_tracer.trackDistX\[-1\] _03569_ _03598_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__16197__A1 _08983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21190__A1 _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__25456__A1 _05696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25454_ _06192_ _06198_ _06238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22666_ _02773_ _03535_ _03536_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_62_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__19895__I _12666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24405_ _05186_ _05187_ _05188_ _05163_ _05189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_216_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21617_ _10448_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_233_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25385_ _06165_ _06168_ _06169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_192_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22597_ _11135_ _07238_ _12229_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_146_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27124_ _01034_ clknet_leaf_117_i_clk rbzero.traced_texVinit\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24336_ _05015_ _05051_ _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24306__I _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21548_ _02233_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__20834__I _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27055_ _00965_ clknet_leaf_133_i_clk rbzero.tex_b1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24267_ _04933_ _05037_ _04987_ _05051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_105_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21479_ _02323_ _02564_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_133_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_26006_ _06738_ _06783_ _06743_ _06784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14020_ rbzero.tex_r1\[16\] _07829_ _07830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23218_ _03978_ _03990_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_8_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22442__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24198_ _04902_ _04981_ _04956_ _04880_ _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__18110__A2 _11249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23149_ _02766_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19563__C _12334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24195__A1 _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25137__I _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21665__I _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15971_ _08822_ _08831_ _09547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__14683__A1 _07222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17710_ _10903_ _10904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14922_ _07802_ _08679_ _08727_ _08728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_26908_ _00818_ clknet_leaf_126_i_clk rbzero.tex_r1\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_18690_ _11670_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_215_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17641_ _10844_ _10859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14853_ _08655_ _08656_ _08658_ _08502_ _08346_ _08659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_26839_ _00749_ clknet_leaf_200_i_clk rbzero.tex_r0\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA_clkbuf_leaf_213_i_clk_I clknet_5_6__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13183__I _06922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13804_ _07610_ _07611_ _07612_ _07614_ _07589_ _07615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_17572_ _10815_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14784_ rbzero.tex_b0\[10\] _07629_ _08591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19311_ rbzero.tex_b1\[34\] rbzero.tex_b1\[33\] _12115_ _12117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__18177__A2 _11269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18195__B _11338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16523_ _09920_ _09977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13735_ _07336_ _07546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15612__B _09278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19242_ _12077_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_168_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16454_ _09903_ _09910_ _09911_ _09912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13666_ _07326_ _07477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__19126__A1 _08161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15405_ _08485_ _09124_ _09125_ _09126_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_94_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19173_ _11251_ _12015_ _12017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_213_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16385_ rbzero.spi_registers.buf_texadd3\[14\] _09851_ _09859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13410__A2 _07218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13597_ _06863_ _07388_ _07391_ _06867_ _07407_ _07408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_183_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18124_ rbzero.wall_tracer.mapY\[6\] rbzero.wall_tracer.mapY\[9\] rbzero.wall_tracer.mapY\[8\]
+ rbzero.wall_tracer.mapY\[10\] _11268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_136_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15336_ _09074_ _09075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15838__I _09429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18055_ rbzero.wall_tracer.trackDistX\[-7\] _11199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_124_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15163__A2 _08940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15267_ _09020_ _09022_ _09018_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_2 _08379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__26607__CLKN clknet_leaf_168_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17006_ rbzero.pov.ready_buffer\[41\] _10403_ _10409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14218_ rbzero.debug_overlay.playerY\[-8\] _08028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_238_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15198_ _08968_ _08969_ _08970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14910__A2 _08698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14149_ _07888_ _07927_ _07958_ _07477_ _07959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_21_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24186__A1 _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18957_ _11849_ _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17908_ _08081_ _11014_ _11052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_207_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18888_ rbzero.traced_texa\[5\] _07279_ _11803_ _11804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_206_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17839_ _10987_ _10988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_222_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer14 net59 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13307__B _07028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer25 _05098_ net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_222_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer36 _05207_ net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_20850_ _01938_ _01939_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14977__A2 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18168__A2 _11301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19509_ _08181_ _12280_ _12281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20781_ _01758_ _01759_ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22520_ rbzero.wall_tracer.texu\[4\] _03429_ _03430_ rbzero.row_render.texu\[4\]
+ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_187_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14729__A2 _08529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22451_ _03391_ _03392_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19668__A2 _11381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21402_ _02485_ _02486_ _02487_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_199_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25170_ _05919_ _05925_ _05954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22382_ _03327_ _10188_ _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24121_ _04904_ _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_21333_ _02278_ _02281_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_40_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23216__A3 _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24052_ _04787_ _04835_ _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_21264_ _12498_ _01723_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14901__A2 _07829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_162_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17963__I _11106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20215_ _12884_ _12987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23003_ _03860_ _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16103__A1 _08990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21195_ _02276_ _02282_ _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20146_ _12917_ _12918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_244_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22727__A2 _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20077_ _12193_ _12224_ _12807_ _12837_ _12849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_24954_ _05724_ _05728_ _05613_ _05738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_231_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23905_ _04246_ _04696_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__18651__I0 _07171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24885_ _05666_ _05668_ _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_213_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26624_ _00534_ clknet_leaf_159_i_clk rbzero.tex_b0\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_68_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23836_ _04660_ _04536_ _04667_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_200_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_218_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26555_ _00465_ clknet_leaf_66_i_clk rbzero.pov.spi_buffer\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23767_ rbzero.wall_tracer.trackDistY\[-1\] _03058_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_184_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20979_ _12482_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_196_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_25506_ _06152_ _06156_ _06290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13520_ _07305_ _07322_ _07330_ _07331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_22718_ _03582_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26486_ _00396_ clknet_leaf_49_i_clk rbzero.debug_overlay.facingX\[-3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23698_ _11216_ _04529_ _04546_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_211_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14048__B _07646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_231_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25437_ _06187_ _06182_ _06220_ _06221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_36_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13451_ rbzero.texV\[8\] _07262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_22649_ _11399_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_97_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16170_ _09675_ _09698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_25368_ _06034_ _06006_ _06152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13382_ _07190_ _07191_ _07192_ _07193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_152_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15121_ rbzero.spi_registers.ss_buffer\[1\] _08867_ _08904_ _08905_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_27107_ _01017_ clknet_leaf_142_i_clk rbzero.tex_b1\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24319_ _04896_ _04898_ _05035_ _05034_ _05060_ _05079_ _05103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_51_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25299_ _06082_ _06083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24255__I2 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14353__B1 _08060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15052_ _08844_ _08845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_27038_ _00948_ clknet_leaf_138_i_clk rbzero.tex_g0\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_120_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14003_ rbzero.tex_r1\[28\] _07810_ _07812_ _07813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__22966__A2 _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_248_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_19860_ _12617_ _12631_ _12632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__26759__CLK clknet_5_3__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18811_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] _11741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19791_ _12476_ _12562_ _12563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16489__I _09944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22179__B1 _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15393__I _09117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18742_ _11700_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15954_ _09518_ _09528_ _09535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23824__B _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14905_ rbzero.tex_b1\[53\] _07561_ _08711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_18673_ _11650_ _11661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15885_ rbzero.spi_registers.buf_leak\[1\] _09482_ _09483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20744__A4 _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14836_ rbzero.tex_b1\[17\] _08250_ _07826_ _08642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17624_ _10845_ rbzero.pov.ready _10256_ _10846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__17070__A2 _10434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24340__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17555_ rbzero.tex_b0\[36\] rbzero.tex_b0\[35\] _10802_ _10806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__21154__A1 _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14767_ rbzero.tex_b0\[17\] _08340_ _08574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13631__A2 _07334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17113__I _08932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16506_ _08106_ _09946_ _09961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13718_ _07507_ _07528_ _07529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22954__I _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17486_ rbzero.tex_b0\[6\] rbzero.tex_b0\[5\] _10765_ _10767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14698_ rbzero.tex_b0\[49\] _08496_ _08335_ _08505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16437_ rbzero.vga_sync.vsync net23 _09895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
X_19225_ _12061_ _12062_ _12065_ _12066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_144_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13649_ _07459_ _07460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_186_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__24643__A2 _05425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19156_ _08149_ _10150_ _12000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_147_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16368_ _09845_ _09846_ _09844_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18107_ _11250_ _11251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_26_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15319_ _07743_ _09058_ _09062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19087_ _11928_ _11929_ _11930_ _11931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_140_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16299_ _09761_ _09795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13147__A1 _06958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18038_ _11181_ rbzero.wall_tracer.trackDistY\[0\] _11177_ _11178_ _11182_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14344__B1 _08010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21209__A2 _13012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14344__C2 _08153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14895__B2 _08564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20000_ _12769_ _12771_ _12772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19989_ _12193_ _12760_ _12761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_185_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23906__A1 _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14140__C _07464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21951_ rbzero.wall_tracer.rcp_fsm.o_data\[-10\] _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_97_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__17061__A2 _10443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20902_ _01801_ _01809_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24670_ _05384_ _05453_ _05454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21882_ _10477_ _10466_ _02914_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_29_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_109_i_clk_I clknet_5_31__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23621_ _03849_ _04259_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_159_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_176_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20833_ _12432_ _12704_ _01682_ _01804_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_49_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26340_ _00250_ clknet_leaf_237_i_clk rbzero.spi_registers.buf_texadd0\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23552_ _04199_ _04259_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__21696__A2 _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_194_Right_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20764_ _01637_ _01763_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_193_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22503_ _03411_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26271_ _00181_ clknet_leaf_17_i_clk rbzero.spi_registers.texadd3\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23483_ _04318_ _04336_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20695_ _01676_ _01768_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25831__A1 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_213_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23896__S _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25222_ _06005_ _06006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20384__I _12260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22434_ _03375_ _03376_ _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25153_ _05884_ _05904_ _05937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22365_ _03312_ _03313_ _03079_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24104_ _04887_ _04888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_102_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14335__B1 _08046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_248_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_21316_ _01712_ _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25084_ _05867_ _05807_ _05863_ _05864_ _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_22296_ _11287_ _03237_ _03257_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_92_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24035_ _04795_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_21247_ _02203_ _02333_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_228_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_228_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21178_ _02252_ _02265_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_229_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14638__B2 _07912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20129_ _12636_ _12637_ _12901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__16102__I _09599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25986_ _06627_ _06622_ _06688_ _06765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_70_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19577__A1 _12255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_24937_ _05718_ _05720_ _05643_ _05721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_169_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15670_ rbzero.spi_registers.buf_texadd2\[7\] _09317_ _09322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24868_ _05647_ _05648_ _05652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_198_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26607_ _00517_ clknet_leaf_168_i_clk rbzero.tex_b0\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14621_ _07803_ _08410_ _08415_ _08420_ _08428_ _08429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_197_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23819_ _11151_ _04619_ _04652_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_240_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24799_ _05579_ _05581_ _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17340_ _10657_ _10653_ _10660_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_200_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14552_ _07461_ _07445_ _08361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_26538_ _00448_ clknet_leaf_23_i_clk rbzero.pov.spi_buffer\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__26075__A1 _06842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_161_Right_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13503_ _07312_ _07313_ _07314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17271_ rbzero.pov.spi_buffer\[22\] _10603_ _10599_ _10609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_101_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14483_ rbzero.tex_g0\[34\] _08291_ _08292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_101_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26469_ _00379_ clknet_leaf_45_i_clk rbzero.debug_overlay.playerY\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24625__A2 _05408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19010_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _11877_ _11880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_16222_ _09735_ _09736_ _09734_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_181_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13434_ gpout0.vpos\[7\] _07226_ _07245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15388__I _06898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer5 _04861_ net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16153_ _09671_ _09685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13365_ _07176_ _07161_ net14 _07177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_248_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_248_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_248_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15104_ _08865_ _08892_ _08893_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_51_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16084_ _09631_ _09632_ _09626_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16866__A2 _10289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13296_ rbzero.spi_registers.texadd2\[4\] _07108_ _07109_ rbzero.spi_registers.texadd1\[4\]
+ _07110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_121_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19912_ _12683_ _12684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15035_ _08827_ _08828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_248_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_236_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19843_ _12612_ _12613_ _12614_ _12615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__22014__I _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_19774_ _12504_ _12544_ _12545_ _12546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_108_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16986_ _10392_ _10393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13301__A1 rbzero.spi_registers.texadd2\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18725_ _11690_ _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15937_ rbzero.spi_registers.spi_buffer\[3\] _09522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14895__C _07839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21914__A3 _10471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15868_ _08928_ _09460_ _09470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18656_ rbzero.tex_r1\[1\] rbzero.tex_r1\[0\] _11651_ _11652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_110_i_clk_I clknet_5_31__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_121_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17607_ _10835_ _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14819_ _07971_ _08625_ _08626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14467__I _07486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18587_ rbzero.tex_r0\[36\] rbzero.tex_r0\[35\] _11608_ _11612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15799_ _09415_ _09416_ _09417_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17538_ _10780_ _10796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_200_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17469_ rbzero.pov.spi_buffer\[73\] _10544_ _10751_ _10756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16554__A1 _09945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25813__A1 _05949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_154_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_154_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19208_ _12016_ _12051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_20480_ _01523_ _01536_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_171_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20638__B1 _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19139_ _11944_ _11982_ _11983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_144_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22150_ rbzero.wall_tracer.visualWallDist\[-4\] _03135_ _03130_ _11073_ _03136_ _03137_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_30_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_11__f_i_clk clknet_3_2_0_i_clk clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21101_ _12465_ _01954_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22081_ _03076_ _03070_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_196_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_35_i_clk_I clknet_5_5__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21989__I0 rbzero.wall_tracer.rcp_fsm.o_data\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_58_Left_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_227_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16609__A2 _08112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21032_ _12689_ _02120_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13540__A1 rbzero.floor_leak\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_238_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25840_ _06623_ _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_226_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19559__A1 rbzero.wall_tracer.size\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25771_ _06527_ _06536_ _06554_ _06555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_22983_ _03839_ _03840_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_24722_ _05239_ _05299_ _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_21934_ _02966_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__17181__C _10357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27441_ _01346_ clknet_leaf_69_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_210_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24653_ net53 _05436_ _05437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21865_ _02905_ _02908_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_26_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Left_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23604_ _04361_ _04455_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27372_ _01277_ clknet_leaf_90_i_clk rbzero.wall_tracer.trackDistY\[-8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20816_ _01862_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_139_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21669__A2 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24584_ _05362_ _05367_ _05368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_21796_ _11047_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26323_ _00233_ clknet_leaf_236_i_clk rbzero.spi_registers.buf_mapdy\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23535_ _04386_ _04387_ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_231_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20747_ _01530_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_135_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26254_ _00164_ clknet_leaf_8_i_clk rbzero.spi_registers.texadd2\[21\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23466_ _04319_ _04303_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20678_ _01673_ _01769_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14020__A2 _07829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25205_ _05979_ _05988_ _05989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22417_ rbzero.wall_tracer.texu\[1\] _03361_ _02715_ _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26185_ _00095_ clknet_leaf_235_i_clk rbzero.spi_registers.texadd0\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23397_ _04236_ _04239_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_104_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25136_ _05408_ _05233_ _05920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13150_ rbzero.spi_registers.texadd3\[6\] _06920_ _06923_ rbzero.spi_registers.texadd2\[6\]
+ _06953_ _06964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_22348_ _11279_ _03290_ _03299_ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Left_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__19408__I _12179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25067_ _05847_ _05850_ _05851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13081_ net23 _06896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_237_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22279_ _03225_ _03241_ _03242_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_72_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_243_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24018_ _04801_ _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14061__B _07587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_208_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16840_ _08184_ _10267_ _10268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_208_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25966__S1 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14087__A2 _07834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15284__A1 _09027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_230_Right_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__24543__A1 _05275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16771_ _10200_ _10180_ _10207_ _10187_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_25969_ _05058_ _06749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13983_ _07244_ _07254_ _07793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_244_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15722_ _09336_ _09361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_18510_ _11568_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_19490_ rbzero.wall_tracer.visualWallDist\[-10\] _12198_ _12262_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Left_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15653_ _09308_ _09309_ _09301_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18441_ rbzero.tex_g1\[37\] rbzero.tex_g1\[36\] _11528_ _11529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21109__A1 _12731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__16784__A1 rbzero.pov.ready_buffer\[65\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14604_ rbzero.tex_g1\[15\] _07807_ _07642_ _08412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18372_ _11489_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_205_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22857__A1 _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15584_ _09257_ _09258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__26048__A1 _05242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19722__A1 _12355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20868__B1 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17323_ _10645_ _10641_ _10647_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_83_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14535_ _08339_ _08341_ _08343_ _08344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_83_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15620__B _09278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17254_ rbzero.pov.spi_buffer\[17\] _10596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14466_ _08201_ _08239_ _08274_ _07802_ _08275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_43_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16205_ rbzero.spi_registers.buf_texadd1\[17\] _09719_ _09724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13417_ _07213_ _07226_ _07227_ _07228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_4_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17185_ _10543_ _10544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14397_ _07628_ _08206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_94_Left_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16136_ _09671_ _09672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_24__f_i_clk_I clknet_3_6_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13348_ _06892_ _07160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__20635__A3 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16067_ rbzero.spi_registers.buf_texadd0\[7\] _09610_ _09620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15511__A2 _09030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13279_ _07053_ _07090_ _07091_ _07092_ _07057_ _07093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__13794__C _07604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15018_ _08815_ _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_209_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19826_ _12589_ _12597_ _12598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22679__I _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19757_ _12526_ _12528_ _12529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_16969_ rbzero.pov.ready_buffer\[33\] _10379_ _10380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15581__I _09254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18708_ rbzero.tex_r1\[24\] rbzero.tex_r1\[23\] _11677_ _11681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_223_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19688_ _12425_ _12447_ _12460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19988__I _12238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18639_ _11641_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14197__I _08006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21650_ rbzero.wall_tracer.rayAddendY\[-6\] _02722_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23896__I0 rbzero.wall_tracer.rcp_fsm.o_data\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20601_ _12989_ _12519_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_21581_ _02663_ _02664_ _02665_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16527__B2 _09918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23320_ _04173_ _04174_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20532_ _01584_ _01603_ _01624_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_90_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14002__A2 _07811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23251_ _04079_ _04106_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20463_ _01457_ _01554_ _01555_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_134_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15750__A2 _09373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22202_ _03177_ _03178_ _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13761__A1 _07478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23182_ _03923_ _03924_ _04034_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_20394_ _01479_ _01481_ _01487_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_247_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22133_ _11992_ _03121_ _03094_ _03122_ _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_30_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26941_ _00851_ clknet_leaf_184_i_clk rbzero.tex_r1\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_22064_ rbzero.wall_tracer.stepDistY\[4\] _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_218_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21015_ _02085_ _02103_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26872_ _00782_ clknet_leaf_165_i_clk rbzero.tex_r0\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__25317__A3 _06100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_25823_ _06571_ _06590_ _06601_ _06606_ _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_215_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__17192__B _10174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21339__A1 _12382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_221_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13816__A2 _07626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18204__A1 _11338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25754_ _06526_ _06537_ _06538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22966_ _02146_ _01383_ _02114_ _02633_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__20011__A1 _12705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_203_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24705_ _05433_ _05487_ _05489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21917_ _02955_ _02939_ _02957_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_25685_ _06424_ _06467_ _06468_ _06469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_85_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22897_ _03754_ _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_27424_ _01329_ clknet_leaf_84_i_clk rbzero.wall_tracer.rcp_fsm.operand\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24636_ _05190_ _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_183_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21848_ _02879_ _10040_ _02886_ _02887_ _02893_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_139_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23500__A2 _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27355_ _01260_ clknet_leaf_80_i_clk rbzero.wall_tracer.trackDistX\[-3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24567_ _05350_ _05351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18307__I _08869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21511__A1 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21779_ rbzero.debug_overlay.vplaneX\[-1\] _11080_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__21511__B2 _12414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17211__I _08805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26306_ _00216_ clknet_leaf_236_i_clk rbzero.spi_registers.buf_othery\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14320_ _08128_ _08039_ _08044_ _08129_ _08130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_23518_ _04272_ _04369_ _04277_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_27286_ _01191_ clknet_leaf_213_i_clk gpout0.hpos\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__20865__A3 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24498_ _05280_ _05281_ _05282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_52_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26237_ _00147_ clknet_leaf_14_i_clk rbzero.spi_registers.texadd2\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14251_ rbzero.debug_overlay.playerY\[-4\] _08061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_162_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23449_ _04212_ _04227_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13202_ rbzero.spi_registers.texadd3\[20\] _07014_ _07009_ rbzero.spi_registers.texadd2\[20\]
+ _07015_ rbzero.spi_registers.texadd1\[20\] _07016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_26168_ _00078_ clknet_leaf_228_i_clk rbzero.color_sky\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14182_ _06871_ _06861_ _07992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25119_ _05885_ _05902_ _05903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13133_ rbzero.spi_registers.texadd3\[9\] _06920_ _06924_ rbzero.spi_registers.texadd2\[9\]
+ _06916_ rbzero.spi_registers.texadd1\[9\] _06947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_26099_ _00009_ clknet_leaf_243_i_clk rbzero.spi_registers.spi_done vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_18990_ _11868_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21027__B1 _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17941_ _11070_ _11071_ _11073_ _11084_ _11085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_13064_ _06870_ _06880_ _06881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19582__B _10305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__18977__I _11850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_218_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17872_ _11009_ _11013_ _11015_ _11016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__20250__A1 rbzero.wall_tracer.stepDistX\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19611_ _12382_ _12383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_16823_ _10250_ _10251_ _10252_ _10253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__16497__I _09926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13807__A2 _07617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19542_ _08029_ _12014_ _12311_ _12313_ _12314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_13966_ _07735_ _07750_ _07776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16754_ _10188_ _10180_ _10192_ _10187_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_220_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15705_ _09336_ _09348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_19473_ _12244_ _12245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16685_ _10115_ _10122_ _10129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13897_ rbzero.debug_overlay.playerX\[-1\] _07708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_186_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18424_ rbzero.tex_g1\[30\] rbzero.tex_g1\[29\] _11517_ _11519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_152_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15636_ _09295_ _09296_ _09290_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16509__A1 _09956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15567_ _09208_ _09245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18355_ _11478_ _11479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17306_ _10611_ _10635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14518_ rbzero.tex_g0\[49\] _07890_ _08327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15498_ _09153_ _09194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__17182__A1 rbzero.pov.ss_buffer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18286_ _11419_ _11420_ _11426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14449_ _08226_ _08258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17237_ rbzero.pov.spi_buffer\[13\] _10580_ _10577_ _10584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13743__A1 _07480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_208_i_clk_I clknet_5_7__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17168_ rbzero.pov.spi_counter\[4\] _10529_ _10531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16119_ _08931_ _09659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14480__I _07549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17099_ _10478_ _10458_ _10479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24755__A1 _05460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20241__A1 _12592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19809_ _12171_ _12579_ _12580_ _12581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_32_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22820_ _02631_ _02637_ _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__23742__B _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22751_ _02739_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_189_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21741__A1 _08175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19511__I _12282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21702_ _08066_ _02740_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25470_ _06002_ _06252_ _06253_ _06254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_22682_ _03549_ _03550_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_192_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24421_ _05201_ _05204_ _05205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_192_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21633_ _02705_ _02709_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_158_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22297__A2 _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15971__A2 _08831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17031__I _06899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27140_ _01050_ clknet_leaf_31_i_clk rbzero.wall_tracer.rayAddendY\[-8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24352_ _05135_ _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21564_ _02529_ _02533_ _02648_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_34_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23303_ _03656_ _03654_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20515_ _01607_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_173_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_27071_ _00981_ clknet_leaf_143_i_clk rbzero.tex_b1\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__24294__I0 _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24283_ _04989_ _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_160_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21495_ _02577_ _02579_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_144_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26022_ _06795_ _06797_ _06798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_144_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23234_ _04081_ _04089_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_127_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20446_ _01498_ _01539_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_127_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14604__B _07642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_23165_ _03962_ _03992_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__25538__A3 _06311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20377_ _01467_ _01470_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_207_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__20480__A1 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22116_ _03087_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23096_ _03951_ _03952_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_223_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24210__A3 _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22047_ _03053_ _03054_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26924_ _00834_ clknet_leaf_126_i_clk rbzero.tex_r1\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_238_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23208__I _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22112__I _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26855_ _00765_ clknet_leaf_187_i_clk rbzero.tex_r0\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_13820_ rbzero.tex_r0\[26\] _07629_ _07630_ _07631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_25806_ _06573_ _06589_ _06590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_230_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26786_ _00696_ clknet_leaf_127_i_clk rbzero.tex_g1\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_23998_ rbzero.wall_tracer.rcp_fsm.operand\[7\] _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_201_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25737_ _05981_ _06089_ _05985_ _05984_ _06521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13751_ rbzero.tex_r0\[47\] _07561_ _07562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_67_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22949_ _03690_ _03806_ _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__21732__A1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_4_i_clk_I clknet_5_4__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_238_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19421__I _12192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_197_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16470_ _09926_ _09927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_157_i_clk_I clknet_5_10__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25668_ _05910_ _05945_ _05965_ _05890_ _06452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_13682_ _07492_ _07493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_211_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15421_ rbzero.spi_registers.buf_floor\[2\] _09137_ _09138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_27407_ _01312_ clknet_leaf_113_i_clk rbzero.wall_tracer.stepDistX\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24619_ _05401_ _05402_ _05403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_167_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25599_ _06381_ _06382_ _06383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19153__A2 _11988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18140_ rbzero.wall_tracer.visualWallDist\[4\] _11284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15352_ _09085_ _09086_ _09073_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_27338_ _01243_ clknet_leaf_36_i_clk rbzero.texu_hot\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14303_ _08110_ _08063_ _08059_ _08112_ _08113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_18071_ _11211_ _11214_ _11215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27269_ _01174_ clknet_leaf_100_i_clk rbzero.wall_tracer.visualWallDist\[9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15283_ _09035_ _09036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__16911__A1 _07705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17022_ _10419_ _10420_ _10414_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14234_ _08043_ _08034_ _08044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_180_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21799__A1 _09989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13909__I _07719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14165_ gpout0.hpos\[3\] _07974_ _07975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22460__A2 _08887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13116_ rbzero.spi_registers.texadd3\[13\] _06928_ _06917_ rbzero.spi_registers.texadd1\[13\]
+ _06930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_111_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__24502__I _05257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14096_ _07498_ _07906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18973_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _11856_ _11859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14150__A1 _07802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17924_ _11000_ _11063_ _11068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_13047_ _06863_ _06864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_219_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17855_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] _10999_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_245_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_244_i_clk clknet_5_0__leaf_i_clk clknet_leaf_244_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__25162__A1 _05871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16806_ _10209_ _10238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22957__I _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17786_ _10952_ rbzero.pov.ready_buffer\[52\] _10955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14998_ _08798_ _08799_ _08800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_220_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19525_ _12296_ _12297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16737_ rbzero.pov.ready _10162_ _10177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13949_ _07216_ _07760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_163_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19456_ _12200_ _12228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16668_ _09917_ _10113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17942__A3 _11068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18407_ _11509_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15619_ rbzero.spi_registers.buf_texadd1\[18\] _09281_ _09284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14475__I _07642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19387_ _12158_ _12159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_174_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16599_ _09988_ _10048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_173_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18338_ _11466_ _11465_ _11467_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13312__C _07052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__17155__A1 _07167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4_0_i_clk_I clknet_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23228__A1 _12212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18269_ _11402_ _11408_ _11411_ _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__16902__A1 rbzero.debug_overlay.playerY\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20300_ _01382_ _01394_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21280_ _02356_ _02366_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25936__C _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19447__A3 _12218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13819__I _07520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20231_ _13000_ _13001_ _12998_ _13003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_229_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24728__A1 _05292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20162_ _12933_ _12667_ _12934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_181_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20093_ _12673_ _12776_ _12865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24970_ _05632_ _05633_ _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__21972__S _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23921_ _11392_ _06895_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_157_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_26640_ _00550_ clknet_leaf_171_i_clk rbzero.tex_b0\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_240_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23852_ rbzero.wall_tracer.trackDistY\[10\] _04681_ _04535_ _04682_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I i_gpout2_sel[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14444__A2 _08206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22803_ _12791_ _02485_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_197_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26571_ _00481_ clknet_leaf_27_i_clk rbzero.pov.spi_buffer\[40\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23783_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] _04616_
+ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_49_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20995_ _02063_ _02083_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25522_ _06305_ _06297_ _06306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_22734_ _03590_ _03596_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_179_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25456__A2 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25453_ _06192_ _06198_ _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14385__I _07185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22665_ _02746_ _03334_ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_192_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24404_ _05080_ _05147_ _05150_ _05114_ _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_62_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_216_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21616_ _09920_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13955__A1 _07750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_233_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25384_ _06166_ _06167_ _06168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_11_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22596_ _07241_ _11132_ _12225_ _03481_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_146_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_233_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_27123_ _01033_ clknet_leaf_117_i_clk rbzero.traced_texVinit\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24335_ net92 _05118_ _05119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_146_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21547_ _02501_ _01919_ _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__18894__A1 _11769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22690__A2 _12499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20336__B _12912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27054_ _00964_ clknet_leaf_133_i_clk rbzero.tex_b1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24266_ _05026_ _05039_ _05049_ _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_16_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21478_ _02450_ _02563_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_26005_ _06777_ _06780_ _06782_ _06783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_95_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23217_ _04029_ _04072_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14380__A1 _07980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20429_ _01521_ _01522_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_24197_ _04827_ _04882_ _04885_ _04980_ _04981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_31_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__26023__B _10988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_248_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_23148_ _03548_ _03897_ _04004_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__24322__I _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22043__S _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_83_i_clk_I clknet_5_28__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14988__C net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23079_ _02621_ _03802_ _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15970_ _08911_ _09545_ _09546_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20205__A1 _12962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23942__A2 _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19071__A1 rbzero.debug_overlay.facingY\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14921_ _08201_ _08703_ _08726_ _08357_ _08727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_26907_ _00817_ clknet_leaf_125_i_clk rbzero.tex_r1\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_199_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold50 _08802_ net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_117_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__21953__A1 _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17640_ _10857_ _10858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_243_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_199_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14852_ rbzero.tex_b1\[12\] _08631_ _08657_ _08658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_26838_ _00748_ clknet_leaf_199_i_clk rbzero.tex_r0\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_89_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13803_ rbzero.tex_r0\[8\] _07579_ _07613_ _07614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14783_ rbzero.tex_b0\[11\] _08300_ _08590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_17571_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _10812_ _10815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_216_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26769_ _00679_ clknet_leaf_125_i_clk rbzero.tex_g1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_231_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19310_ _12116_ _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_16522_ _09974_ _09975_ _09976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13734_ _07534_ _07545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19241_ rbzero.tex_b1\[4\] rbzero.tex_b1\[3\] _12073_ _12077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16453_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] _09911_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13665_ _07441_ _07457_ _07467_ _07474_ _07475_ _07476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_156_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15404_ _09067_ _09126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_213_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16384_ _09857_ _09858_ _09856_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_19172_ _12015_ _12016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_171_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13596_ _07405_ _07406_ _07407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17137__A1 rbzero.pov.ready_buffer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15335_ _08877_ _09074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18123_ rbzero.wall_tracer.mapX\[9\] rbzero.wall_tracer.mapX\[8\] rbzero.wall_tracer.mapX\[10\]
+ rbzero.wall_tracer.mapY\[7\] _11267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__22681__A2 _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18054_ _11197_ _11198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_15266_ rbzero.spi_registers.buf_otherx\[1\] _09021_ _09022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22017__I _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17005_ _08071_ _10401_ _10408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14217_ _07706_ _08023_ _08026_ _07685_ _08027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_15197_ _08951_ _08969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14148_ _07928_ _07944_ _07957_ _07958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__22180__C _09918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__25383__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__24186__A2 _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14079_ _07608_ _07889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18956_ rbzero.tex_g0\[16\] rbzero.tex_g0\[15\] _11845_ _11849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_207_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_183_i_clk clknet_5_2__leaf_i_clk clknet_leaf_183_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input5_I i_gpout0_sel[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17907_ _11048_ _11049_ _11050_ _11051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_18887_ rbzero.traced_texa\[4\] rbzero.texV\[4\] _11802_ _11803_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__21944__A1 _09925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13374__I net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17838_ _07166_ _10987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_179_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_175_Right_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer15 _05814_ net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14426__A2 _07872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer26 _05001_ net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_156_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer37 _05013_ net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_83_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23697__A1 _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17769_ _10934_ _10943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_124_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_198_i_clk clknet_5_13__leaf_i_clk clknet_leaf_198_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_19508_ _11385_ _12280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20780_ _01756_ _01757_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_159_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25438__A2 _06102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14419__B _08220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19439_ _12210_ _12211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15926__A2 _09498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_121_i_clk clknet_5_18__leaf_i_clk clknet_leaf_121_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_44_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22450_ rbzero.wall_tracer.texu\[4\] _03323_ _03111_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__17128__A1 _09928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13937__B2 _07743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_199_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21401_ _12807_ _12699_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_174_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22381_ _12907_ _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24120_ _04733_ _04903_ _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_21332_ _02417_ _02282_ _02418_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_136_i_clk clknet_5_15__leaf_i_clk clknet_leaf_136_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_248_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24051_ _04829_ _04834_ _04794_ _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__24264__I3 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21263_ _12732_ _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19825__B1 _12594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_105_i_clk_I clknet_5_30__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23621__A1 _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22371__B rbzero.wall_tracer.wall\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23002_ _02251_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_20214_ _12893_ _12898_ _12985_ _12986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_21194_ _02278_ _02281_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20145_ _11386_ _12915_ _12916_ _12917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_110_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14665__A2 _07916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24953_ _05727_ _05732_ _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20076_ _12841_ _12817_ _12842_ _12848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_231_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23904_ _03022_ _04711_ _04714_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24884_ _05618_ _05667_ _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23835_ _04348_ _04666_ _04528_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_26623_ _00533_ clknet_leaf_157_i_clk rbzero.tex_b0\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_213_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_218_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26554_ _00464_ clknet_leaf_66_i_clk rbzero.pov.spi_buffer\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_235_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_23766_ rbzero.wall_tracer.trackDistY\[-1\] _03058_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_194_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20978_ _02066_ _12483_ _12919_ _01704_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_32_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22360__A1 rbzero.mapdyw\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25505_ _06281_ _06285_ _06288_ _06289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_22717_ _03581_ rbzero.wall_tracer.trackDistX\[-3\] _03569_ _03582_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13233__B _07046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26485_ _00395_ clknet_leaf_52_i_clk rbzero.debug_overlay.facingX\[-4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23697_ _04542_ _04545_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_193_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25436_ _06194_ _06188_ _06220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13928__A1 _07736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13450_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] _07261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_193_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22648_ _02731_ _03518_ _03520_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__17119__A1 _09942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25367_ _06149_ _06150_ _06151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_13381_ gpout0.vpos\[0\] _07192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__23860__A1 _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22663__A2 _12214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22579_ _03469_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15120_ rbzero.spi_registers.spi_counter\[6\] rbzero.spi_registers.spi_counter\[5\]
+ _08848_ _08904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_91_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24318_ _05061_ _05101_ _05045_ _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__20674__A1 _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27106_ _01016_ clknet_leaf_142_i_clk rbzero.tex_b1\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25298_ _06079_ _06080_ _06081_ _05728_ _06082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_16_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24255__I3 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14353__A1 _08161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15051_ _08842_ _08843_ _08844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_27037_ _00947_ clknet_leaf_137_i_clk rbzero.tex_g0\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24249_ net54 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__14353__B2 _08162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14002_ rbzero.tex_r1\[29\] _07811_ _07812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_75_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput40 net40 o_tex_csb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__15674__I _09289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_246_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18810_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] _11740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_248_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_208_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19790_ _12561_ _12562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__22179__B2 _11291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14656__A2 _08448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18741_ rbzero.tex_r1\[38\] rbzero.tex_r1\[37\] _11698_ _11700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15953_ rbzero.spi_registers.buf_vshift\[2\] _09531_ _09534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_216_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14904_ rbzero.tex_b1\[55\] _07597_ _08603_ _08710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_18672_ _11660_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15884_ _09481_ _09482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_216_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_17623_ _10844_ _10845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__15623__B _09278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14835_ rbzero.tex_b1\[16\] _08248_ _08641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_231_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_106_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17554_ _10805_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14766_ rbzero.tex_b0\[16\] _08342_ _08573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16505_ _08103_ _09956_ _09959_ _09960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_13717_ _07517_ _07527_ _07528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_128_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17485_ _10766_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14697_ rbzero.tex_b0\[48\] _08277_ _08504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__20901__A2 _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16030__A1 _09591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19224_ _12055_ _12063_ _12064_ _12065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_16436_ _09894_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_184_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13648_ _07419_ _07459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_85_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__22103__A1 _09948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22103__B2 _12834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19155_ _11998_ _11999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_143_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13395__A2 _07202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23851__A1 _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13579_ _07355_ _07356_ _07387_ _07390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_16367_ _08955_ _09842_ _09846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_186_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__20665__A1 _12472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18106_ rbzero.map_rom.i_row\[4\] _11250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_15318_ _09059_ _09061_ _09055_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19086_ _08157_ _09991_ _11930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16298_ _08990_ _09793_ _09794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14344__A1 _08151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18037_ _11169_ _11181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14344__B2 _08152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15249_ rbzero.spi_registers.spi_buffer\[23\] _08917_ _09010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_244_Right_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15584__I _09257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19988_ _12238_ _12760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14647__A2 _08300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15844__A1 _08928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18939_ _11839_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_126_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Left_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21950_ _02980_ _02984_ _02987_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_207_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22590__A1 rbzero.wall_tracer.wall\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20901_ _01760_ _01762_ _01881_ _01882_ _01869_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_TAPCELL_ROW_2_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21881_ _02918_ _02923_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_29_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23620_ _04214_ _04217_ _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20832_ _12780_ _01578_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_176_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22342__A1 _11281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14280__B1 _08060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_31_i_clk_I clknet_5_22__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23551_ _03849_ _04080_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_65_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20763_ _01798_ _01853_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_65_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__26084__A2 _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22502_ _03409_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_174_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26270_ _00180_ clknet_leaf_17_i_clk rbzero.spi_registers.texadd3\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23482_ _04335_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_190_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20694_ _01669_ _01672_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_114_Left_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_174_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23041__I _12035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_213_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25221_ _05869_ _05909_ _06005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22433_ _03364_ _03367_ _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_220_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14583__B2 _07826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23842__A1 _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22645__A2 _12395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20656__A1 _12658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25152_ _05932_ _05935_ _05936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22364_ _02784_ _03248_ rbzero.wall_tracer.wall\[0\] _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_190_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24103_ _04875_ _04886_ _04825_ _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_21315_ _02223_ _02240_ _02401_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__14335__A1 _08143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25083_ _05825_ _05867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_20_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_22295_ _03110_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_92_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_211_Right_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14886__A2 _07577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_248_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_24034_ _04812_ _04775_ _04817_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_21246_ _02220_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_57_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__16088__A1 _08973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15494__I _09190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_228_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_228_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21177_ _02255_ _02264_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_123_Left_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20128_ _12883_ _12899_ _12900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_25985_ _06752_ _06761_ _06763_ _06707_ _06764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_70_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__26020__C _06737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13310__A2 _07108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_20059_ _12825_ _12831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_24936_ _05719_ _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_99_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output44_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24867_ _05650_ _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_240_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16260__A1 _08939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_26606_ _00516_ clknet_leaf_170_i_clk rbzero.tex_b0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_14620_ _07608_ _08427_ _08428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23818_ _04121_ _04651_ _04625_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_24798_ _05579_ _05581_ _05582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_67_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14551_ rbzero.row_render.texu\[0\] _08360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_23749_ rbzero.wall_tracer.trackDistY\[-3\] _03053_ _04583_ _04591_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26537_ _00447_ clknet_leaf_22_i_clk rbzero.pov.spi_buffer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_200_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19569__C _12325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_132_Left_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_166_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13502_ _07266_ _07271_ _07313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14482_ _07523_ _08291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17270_ rbzero.pov.spi_buffer\[21\] _10608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_153_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26468_ _00378_ clknet_leaf_44_i_clk rbzero.debug_overlay.playerY\[-6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25822__A2 _06605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16221_ _09008_ _09732_ _09736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13433_ gpout0.vpos\[3\] _07244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_25419_ _06202_ _06042_ _06203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_26399_ _00309_ clknet_leaf_3_i_clk rbzero.spi_registers.buf_texadd2\[19\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19501__A2 _12267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16152_ _09683_ _09684_ _09678_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13364_ _07175_ _07176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__19585__B _12245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer6 _05196_ net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_248_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_14__f_i_clk_I clknet_3_3_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_248_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15103_ rbzero.spi_registers.spi_counter\[1\] _08891_ _08893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_248_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16083_ _08968_ _09624_ _09632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13295_ _07015_ _07109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_146_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19911_ _12489_ _12683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15034_ rbzero.spi_registers.spi_cmd\[0\] _08827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_121_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_141_Left_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19842_ _12546_ _12566_ _12614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_208_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23835__B _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14629__A2 _07898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19773_ _12468_ _12485_ _12545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_16985_ _10391_ _10392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13301__A2 _07108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18724_ rbzero.tex_r1\[31\] rbzero.tex_r1\[30\] _11687_ _11690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15936_ rbzero.spi_registers.buf_othery\[3\] _09510_ _09521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22572__A1 _11279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22572__B2 rbzero.traced_texa\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18655_ _11650_ _11651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15867_ rbzero.spi_registers.buf_floor\[3\] _09464_ _09469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13652__I _07462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17606_ rbzero.tex_b0\[58\] rbzero.tex_b0\[57\] _10833_ _10835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14818_ _07697_ _08624_ _08625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_121_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18586_ _11611_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__21127__A2 _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15798_ _09383_ _09417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_147_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17537_ _10795_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16963__I _10373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14749_ rbzero.tex_b0\[25\] _07499_ _08556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_50_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19740__A2 _11070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17468_ rbzero.pov.spi_buffer\[72\] _10755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_184_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19207_ _12045_ _12050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_154_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_16419_ _09667_ _09876_ _09884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_171_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17399_ rbzero.pov.spi_buffer\[54\] _10704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19138_ _11945_ _11917_ _11982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__25577__A1 _05977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19069_ rbzero.wall_tracer.mapY\[5\] _11913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21100_ _02070_ _02072_ _02067_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14868__A2 _07595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22080_ rbzero.wall_tracer.stepDistY\[9\] _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_125_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__21989__I1 rbzero.wall_tracer.size\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13827__I _07449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21031_ _01924_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16203__I _09711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13540__A2 _07325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15817__A1 rbzero.spi_registers.texadd3\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16490__A1 _09942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25770_ _06528_ _06535_ _06554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_22982_ _03680_ _03698_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_179_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24721_ _05257_ _05231_ _05505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_21933_ _02921_ _02963_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15045__A2 _08831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_27440_ _01345_ clknet_leaf_70_i_clk rbzero.wall_tracer.rcp_fsm.o_data\[-7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24652_ _05275_ _05232_ _05300_ _05257_ _05436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__26494__D _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__22875__I _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21864_ _02906_ _02907_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_210_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22315__A1 _11291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25251__I _06034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23603_ _04440_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_139_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20815_ _12950_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24583_ _05366_ _05367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_27371_ _01276_ clknet_leaf_90_i_clk rbzero.wall_tracer.trackDistY\[-9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21795_ _02840_ _02843_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_166_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26322_ _00232_ clknet_leaf_236_i_clk rbzero.spi_registers.buf_mapdy\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23534_ _04292_ _04382_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_20746_ _01835_ _01836_ _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26253_ _00163_ clknet_leaf_8_i_clk rbzero.spi_registers.texadd2\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14556__A1 _07433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23465_ _04216_ _04226_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14393__I _07916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20677_ _01676_ _01768_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25204_ _05986_ _05987_ _05988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_163_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22416_ _03322_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26184_ _00094_ clknet_leaf_235_i_clk rbzero.spi_registers.vshift\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23291__A2 _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23396_ _04245_ _04246_ _04249_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_162_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25568__A1 _06328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25135_ _05895_ _05898_ _05919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_189_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22347_ _09926_ _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_131_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14859__A2 _08248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13080_ rbzero.wall_tracer.rcp_fsm.state\[0\] _06895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_25066_ _05848_ _05849_ _05850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22278_ rbzero.wall_tracer.visualWallDist\[-4\] _03237_ _03229_ _03242_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_72_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24017_ rbzero.wall_tracer.rcp_fsm.operand\[-8\] rbzero.wall_tracer.rcp_fsm.operand\[-9\]
+ rbzero.wall_tracer.rcp_fsm.operand\[-10\] rbzero.wall_tracer.rcp_fsm.operand\[-11\]
+ _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA__13531__A2 _07337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21229_ _02290_ _02300_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_243_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_208_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_208_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__24543__A2 _05296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16770_ rbzero.pov.ready_buffer\[63\] _10201_ _10202_ _10206_ _10207_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_25968_ _06683_ _06732_ _06747_ _06699_ _06748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_13982_ _06891_ _07080_ _07780_ _07792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_244_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15721_ rbzero.spi_registers.buf_texadd2\[20\] _09353_ _09360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24919_ _05694_ _05700_ _05703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_198_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_25899_ _06634_ _06665_ _06671_ _06681_ _06682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_213_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18440_ _11522_ _11528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15652_ rbzero.spi_registers.buf_texadd2\[2\] _09306_ _09309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_103_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14603_ rbzero.tex_g1\[14\] _07805_ _08411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14795__A1 _08595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18371_ rbzero.tex_g1\[7\] rbzero.tex_g1\[6\] _11486_ _11489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__22857__A2 _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15583_ _08882_ _09257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_139_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19722__A2 _12357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20868__A1 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17322_ rbzero.pov.spi_buffer\[35\] _10638_ _10646_ _10647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_83_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14534_ rbzero.tex_g0\[60\] _08342_ _08343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14547__A1 _08333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17253_ _10593_ _10594_ _10595_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14465_ _08201_ _08273_ _08274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16204_ _09720_ _09722_ _09723_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_221_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13416_ gpout0.vpos\[5\] _07227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14396_ _07463_ _08203_ _08204_ _08205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_17184_ _10542_ _10543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_181_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_221_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16135_ _09670_ _09671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_13347_ net13 net12 _07159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13770__A2 _07579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20635__A4 _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16066_ _09618_ _09619_ _09615_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13278_ _06906_ _06976_ _07092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_228_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_219_Left_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_114_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__21045__A1 _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13647__I rbzero.row_render.side vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15017_ _08807_ rbzero.wall_tracer.rcp_fsm.state\[4\] _08815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_20_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__16023__I _09564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21596__A2 _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19825_ _12590_ _12593_ _12594_ _12596_ _12597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_235_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_19756_ _12527_ _12386_ _12528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_16968_ _10378_ _10379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_34_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18707_ _11680_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_189_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15919_ _08962_ _09508_ _09509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19687_ _12425_ _12447_ _12459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_190_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_204_i_clk_I clknet_5_13__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16899_ _08061_ _10301_ _10319_ _10320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__20020__A2 _12788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18638_ rbzero.tex_r0\[58\] rbzero.tex_r0\[57\] _11639_ _11641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_228_Left_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_177_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14786__A1 _08565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18569_ _11601_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23896__I1 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20600_ _01591_ _01592_ _01691_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21580_ _02503_ _02505_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_191_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__16527__A2 _09977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20531_ _01606_ _01623_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14538__A1 rbzero.tex_g0\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19937__C _12192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23250_ _04090_ _04105_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20462_ _01455_ _01549_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_134_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22201_ _11282_ _03166_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__21284__A1 _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23181_ _03920_ _04034_ _04035_ _03926_ _04036_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XPHY_EDGE_ROW_237_Left_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_20393_ _01482_ _01485_ _01486_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer16_I _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22132_ rbzero.wall_tracer.visualWallDist\[-7\] _03100_ _03117_ _11078_ _03122_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_112_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23025__A2 _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_22063_ _03064_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_26940_ _00850_ clknet_leaf_184_i_clk rbzero.tex_r1\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_225_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__25246__I _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21014_ _02101_ _02102_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_199_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26871_ _00781_ clknet_leaf_165_i_clk rbzero.tex_r0\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_96_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15772__I _09117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25822_ _06602_ _06605_ _06606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__24525__A2 _05308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__22536__A1 rbzero.wall_tracer.visualWallDist\[-7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25753_ _06527_ _06536_ _06537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22965_ _02271_ _01919_ _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_246_Left_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_223_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19952__A2 _12430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_203_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24704_ _05433_ _05487_ _05488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_21916_ _10477_ _02956_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_25684_ _06426_ _06466_ _06468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__24289__A1 _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22896_ _02571_ _02687_ _03753_ _03754_ _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_222_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_27423_ _01328_ clknet_leaf_82_i_clk rbzero.wall_tracer.rcp_fsm.operand\[-1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24635_ _05418_ _05310_ _05419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_167_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21847_ _02891_ _02892_ _09899_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27354_ _01259_ clknet_leaf_81_i_clk rbzero.wall_tracer.trackDistX\[-4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24566_ _05305_ _05350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16518__A2 _09971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21778_ _12216_ _02703_ _02828_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__18763__I0 rbzero.tex_r1\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26305_ _00215_ clknet_leaf_215_i_clk rbzero.spi_registers.buf_othery\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_23517_ _04272_ _04369_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_20729_ _12423_ _12918_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_24497_ _05033_ _05185_ _05281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27285_ _01190_ clknet_leaf_211_i_clk gpout0.hpos\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15012__I _08810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14250_ _08059_ _08060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_208_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_23448_ _04268_ _04301_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_26236_ _00146_ clknet_leaf_246_i_clk rbzero.spi_registers.texadd2\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__24325__I _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13201_ _06998_ _07015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__21275__A1 _12692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14181_ _07985_ _07987_ _07990_ _07991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_23379_ _04140_ _04233_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__18323__I _10271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26167_ _00077_ clknet_leaf_227_i_clk rbzero.color_sky\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13132_ _06945_ _06946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_25118_ _05887_ _05901_ _05902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_clkbuf_leaf_0_i_clk_I clknet_5_1__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24213__A1 _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26098_ _00008_ clknet_leaf_229_i_clk rbzero.spi_registers.ss_buffer\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_237_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_153_i_clk_I clknet_5_11__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__21027__A1 _12816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__21027__B2 _12675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25049_ _05773_ _05832_ _05791_ _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_17940_ _11074_ _11076_ _11078_ _11083_ _11084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_13063_ _06875_ _06876_ _06879_ _06880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_237_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__22775__A1 _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17871_ rbzero.debug_overlay.facingX\[-7\] _11014_ _11015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__16778__I _09855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19610_ _12381_ _12382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_16822_ _10181_ _10252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_219_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_217_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19541_ _11954_ _11999_ _12312_ _12005_ _12313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_16753_ rbzero.pov.ready_buffer\[61\] _10183_ _10179_ _10191_ _10192_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_13965_ _07774_ _07775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__16206__A1 _08994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15704_ rbzero.spi_registers.buf_texadd2\[16\] _09340_ _09347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_85_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19943__A2 _12692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19472_ _11382_ _12244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_16684_ rbzero.wall_tracer.rayAddendY\[8\] _10128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_158_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13896_ _07192_ _07707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_18423_ _11518_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_201_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15635_ rbzero.spi_registers.buf_texadd1\[22\] _09293_ _09296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14768__A1 _08339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_78_i_clk_I clknet_5_28__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18354_ _07041_ _06876_ _06860_ _11478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_51_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15566_ rbzero.spi_registers.texadd1\[5\] _09243_ _09244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17305_ rbzero.pov.spi_buffer\[30\] _10634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_138_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14517_ rbzero.tex_g0\[48\] _07617_ _08326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18285_ _11402_ _11423_ _11425_ _00660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_151_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15497_ rbzero.spi_registers.texadd0\[11\] _09192_ _09193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_151_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15193__A1 _08965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17236_ _10571_ _10583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14448_ rbzero.tex_g0\[13\] _08202_ _08257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14761__I _07835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17167_ rbzero.pov.spi_counter\[4\] _10529_ _10530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_80_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__18131__A1 rbzero.debug_overlay.playerY\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14379_ _08179_ _08188_ _07195_ _08189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_16118_ _09005_ _09657_ _09658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__26444__CLK clknet_5_25__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17098_ _10477_ _10478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__16693__A1 _10015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16049_ _09518_ _09601_ _09607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__20241__A2 _13012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19808_ rbzero.wall_tracer.size\[7\] _12514_ _12580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22518__A1 rbzero.wall_tracer.texu\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19739_ rbzero.wall_tracer.stepDistX\[-2\] _12511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_193_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22750_ _03607_ _03610_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_144_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__18993__I0 rbzero.tex_g0\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21701_ _11913_ _12051_ _12028_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__21741__A2 _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22681_ rbzero.wall_tracer.trackDistX\[-8\] _03539_ _03542_ _03550_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14759__B2 _08564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24420_ _05025_ _05169_ _05203_ net55 _05204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21632_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] _02709_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19698__A1 _12267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__23494__A2 _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13431__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_24351_ _04742_ _04897_ _05135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_180_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21563_ _02531_ _02532_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_23302_ _12428_ _02595_ _04039_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_20514_ _12917_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27070_ _00980_ clknet_leaf_144_i_clk rbzero.tex_b1\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24282_ _05065_ _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__24443__A1 _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_21494_ _02528_ _02534_ _02578_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__24294__I1 _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26021_ _06659_ _06796_ _06797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_23233_ _04083_ _04088_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_127_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_20445_ _01515_ _01538_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_166_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23164_ _03964_ _03991_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__19870__A1 _12172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20376_ _12398_ _01469_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__23917__C _11473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_219_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_189_Right_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_22115_ _11994_ _03095_ _03105_ rbzero.wall_tracer.visualWallDist\[-9\] _03106_ _03107_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__20480__A2 _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23095_ _03945_ _03950_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22757__A1 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__24210__A4 _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22046_ _03038_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_26923_ _00833_ clknet_leaf_135_i_clk rbzero.tex_r1\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_205_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_26854_ _00764_ clknet_leaf_191_i_clk rbzero.tex_r0\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__21009__I _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25805_ _06576_ _06588_ _06589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_243_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26785_ _00695_ clknet_leaf_127_i_clk rbzero.tex_g1\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_97_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23997_ _04784_ _04785_ _04786_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_214_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25736_ _05235_ _06007_ _06520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_202_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13750_ _07483_ _07561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22948_ _03695_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_168_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13670__A1 _07321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_238_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23224__I _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_238_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_25667_ _06400_ _06449_ _06450_ _06451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13681_ _07442_ _07492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_22879_ _03735_ _03737_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13750__I _07483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27406_ _01311_ clknet_leaf_113_i_clk rbzero.wall_tracer.stepDistX\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15420_ _09029_ _09137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_24618_ _05361_ _05366_ _05374_ _05364_ _05352_ _05402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_195_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25598_ _06181_ _06187_ _06184_ _05990_ _06382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_80_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19153__A3 _11989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_27337_ _01242_ clknet_leaf_92_i_clk rbzero.trace_state\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15351_ rbzero.spi_registers.buf_mapdxw\[0\] _09078_ _09086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_24549_ _05332_ _05333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__22284__B _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14302_ _08111_ _08112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_202_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18070_ _11212_ _11209_ rbzero.wall_tracer.trackDistY\[-11\] _11213_ _11214_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_164_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27268_ _01173_ clknet_leaf_100_i_clk rbzero.wall_tracer.visualWallDist\[8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15282_ _09034_ _09035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16911__A2 _08061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17021_ rbzero.pov.ready_buffer\[23\] _10412_ _10420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14922__A1 _07802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26219_ _00129_ clknet_leaf_6_i_clk rbzero.spi_registers.texadd1\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14233_ _08037_ _08020_ _08043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_124_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27199_ _01104_ clknet_leaf_74_i_clk rbzero.wall_tracer.size_full\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14164_ gpout0.hpos\[2\] _07187_ _07974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_22_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_156_Right_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13115_ rbzero.spi_registers.texadd3\[14\] _06928_ _06925_ rbzero.spi_registers.texadd2\[14\]
+ _06929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_237_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14095_ rbzero.tex_r1\[40\] _07641_ _07905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_18972_ _11858_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13489__A1 rbzero.texV\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17923_ _10997_ _11066_ _11067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_13046_ _06862_ _06863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_219_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19613__A1 _12299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14150__A2 _07887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__20223__A2 _12296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17854_ _08071_ rbzero.wall_tracer.rayAddendX\[7\] _10998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16805_ _08171_ _10215_ _10237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_205_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__25162__A2 _05908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__17841__B _10988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17785_ _10946_ _10954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_227_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14997_ gpout0.vpos\[0\] _08776_ _08782_ _07180_ _07178_ _08781_ _08799_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_89_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19524_ _12287_ _12288_ _12293_ _12295_ _12296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_16736_ _08180_ _10176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13948_ _07220_ _07757_ _07758_ _07759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_152_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__21723__A2 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19455_ _07698_ _12007_ _12226_ _12227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__24348__S1 _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16667_ _10109_ _10111_ _10112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13879_ _07200_ rbzero.debug_overlay.playerY\[1\] _07690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_202_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18406_ rbzero.tex_g1\[22\] rbzero.tex_g1\[21\] _11507_ _11509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15618_ rbzero.spi_registers.texadd1\[18\] _09279_ _09283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19386_ _12157_ _12158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16598_ _10043_ _10046_ _10047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__23476__A2 _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_18337_ _11466_ _11465_ _10751_ _11467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15549_ rbzero.spi_registers.texadd1\[1\] _09230_ _09231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__17155__A2 rbzero.pov.ss_buffer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20707__B _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18268_ _11403_ _11410_ _11411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__24425__A1 _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__23228__A2 _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17219_ rbzero.pov.spi_buffer\[8\] _10570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14913__B2 _08558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18199_ _11111_ _11343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_142_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20230_ _12998_ _13000_ _13001_ _13002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_168_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__24728__A2 _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20161_ _12209_ _12933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14141__A2 _07460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20092_ _12776_ _12861_ _12862_ _12863_ _12864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_243_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13835__I _07524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23920_ _04724_ _04725_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_146_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__23753__B _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_23851_ _04514_ _04680_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22802_ _01956_ _03660_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_26570_ _00480_ clknet_leaf_64_i_clk rbzero.pov.spi_buffer\[39\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_211_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23782_ _11184_ rbzero.wall_tracer.stepDistY\[2\] _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_20994_ _02074_ _02082_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__17918__A1 _08079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_101_i_clk_I clknet_5_27__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_25521_ _06298_ _06304_ _06305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22733_ _02737_ _03594_ _03595_ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_179_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__23979__I _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25452_ _06200_ _06210_ _06236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_22664_ _11205_ _03533_ _03534_ _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_149_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24403_ _05158_ _05179_ _05036_ _05187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_62_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_21615_ _10449_ _02694_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_192_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_25383_ _05921_ _06032_ _06167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_22595_ _12170_ _03082_ _03480_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_35_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_233_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_233_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_27122_ _01032_ clknet_leaf_115_i_clk rbzero.traced_texVinit\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_24334_ _05117_ _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_21546_ _02629_ _02630_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15157__A1 _08935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__24416__A1 _05186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13168__B1 _06981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24265_ _05026_ _05048_ _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27053_ _00963_ clknet_leaf_144_i_clk rbzero.tex_b1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_209_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_21477_ _02457_ _02562_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__23928__B _10508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26004_ _06672_ _06781_ _06782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_23216_ _04033_ _04046_ _04071_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_133_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_20428_ _12262_ _01435_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_24196_ _04905_ _04944_ _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_95_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23147_ _03898_ _04003_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_20359_ rbzero.traced_texVinit\[0\] _10020_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_219_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_26_i_clk_I clknet_5_20__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14132__A2 _07940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23078_ _03820_ _03828_ _03934_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_140_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22029_ _03041_ _03039_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14920_ _08355_ _08714_ _08725_ _08726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_26906_ _00816_ clknet_leaf_125_i_clk rbzero.tex_r1\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_175_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__16121__I _09660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold40 _01026_ net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__13891__A1 _07701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_199_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14851_ rbzero.tex_b1\[13\] _07906_ _08657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_26837_ _00747_ clknet_leaf_196_i_clk rbzero.tex_r0\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_215_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13802_ _07586_ _07613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_17570_ _10814_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14782_ _08459_ _08587_ _08588_ _08589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_26768_ _00678_ clknet_leaf_125_i_clk rbzero.tex_g1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_86_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16521_ _09966_ _09969_ _09975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_25719_ _06487_ _06488_ _06502_ _06503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_202_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13733_ rbzero.tex_r0\[39\] _07543_ _07544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_196_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_26699_ _00609_ clknet_leaf_63_i_clk rbzero.pov.ready_buffer\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19240_ _12076_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16452_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] _09909_
+ _09910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_13664_ _07436_ _07475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15403_ rbzero.spi_registers.buf_sky\[3\] _09080_ _09125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_19171_ _12014_ _12015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_94_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16383_ rbzero.spi_registers.spi_buffer\[13\] _09853_ _09858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_225_Right_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13595_ _06872_ _07394_ _07388_ _06862_ _07406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_213_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18122_ _11254_ _11258_ _11262_ _11265_ _11266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_108_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15334_ _09071_ _09072_ _09073_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__20141__A1 rbzero.wall_tracer.size\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18053_ rbzero.wall_tracer.trackDistY\[-7\] _11197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__16896__A1 rbzero.debug_overlay.playerY\[-4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15265_ _08884_ _09021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__22742__B _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17004_ _06899_ _10407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14216_ _07997_ _08025_ _08026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__24513__I _05296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15196_ rbzero.spi_registers.spi_buffer\[11\] _08968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14147_ _07555_ _07950_ _07956_ _07957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_6_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14123__A2 _07632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__25383__A2 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14078_ _07570_ _07888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_18955_ _11848_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_163_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17906_ _08084_ _11047_ _11050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18886_ _11786_ _11801_ _11802_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_206_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__17073__A1 _08128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17837_ _10845_ _10753_ _10982_ _10986_ _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__23146__A1 _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_169_Left_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_233_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer16 _04862_ net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_206_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer27 _05001_ net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xrebuffer38 _05195_ net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_156_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17768_ _10935_ _10681_ _10939_ _10942_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__13634__A1 _07443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_141_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_19507_ _08048_ _12168_ _12278_ _12279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__18022__B1 _11165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16719_ net16 _10160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_5_3__f_i_clk_I clknet_3_0_0_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14486__I _07496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_17699_ _10874_ _10897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19438_ _12209_ _12210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__19498__B _12269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13937__A2 _07678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19369_ _12149_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21400_ _12782_ _02362_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_174_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22380_ _01661_ _03325_ _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_178_Left_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_21331_ _02273_ _02283_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_199_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24050_ rbzero.wall_tracer.rcp_fsm.operand\[6\] rbzero.wall_tracer.rcp_fsm.operand\[5\]
+ _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_163_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_21262_ _01982_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_170_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19825__A1 _12590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__19825__B2 _12596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_23001_ _03735_ _03737_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__16639__A1 _09897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20213_ _12888_ _12892_ _12985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21193_ _02279_ _02280_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_198_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_229_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_20144_ rbzero.wall_tracer.stepDistX\[1\] _12316_ _12916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__22188__A2 _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_20075_ _12845_ _12846_ _12847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_24952_ _05721_ _05734_ _05735_ _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_225_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_187_Left_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_23903_ _04125_ _04696_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__25126__A2 _05869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_24883_ _05617_ _05614_ _05615_ _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__19252__I _12072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_26622_ _00532_ clknet_leaf_162_i_clk rbzero.tex_b0\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_174_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23834_ _04661_ _04664_ _04665_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_240_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__23688__A2 _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_252_i_clk_I clknet_5_0__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_2__f_i_clk clknet_3_0_0_i_clk clknet_5_2__leaf_i_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_26553_ _00463_ clknet_leaf_66_i_clk rbzero.pov.spi_buffer\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_20977_ _12477_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_23765_ _11170_ rbzero.wall_tracer.stepDistY\[0\] _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_235_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25504_ _06286_ _06287_ _06288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_221_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_22716_ _03556_ _03579_ _03580_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_26484_ _00394_ clknet_leaf_50_i_clk rbzero.debug_overlay.facingX\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_193_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_23696_ _02751_ _04544_ _03536_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_25435_ _06214_ _06218_ _06219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_211_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_22647_ _12775_ _12864_ _03519_ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__14050__A1 rbzero.tex_r1\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19364__I0 rbzero.tex_b1\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_196_Left_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13380_ gpout0.vpos\[1\] _07191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_25366_ _06109_ _06113_ _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__22118__I _09897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_22578_ rbzero.wall_tracer.wall\[0\] _08364_ _09900_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__23860__A2 _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27105_ _01015_ clknet_leaf_142_i_clk rbzero.tex_b1\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24317_ _04886_ _04970_ _05038_ _05101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_21529_ _02611_ _02613_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_243_i_clk clknet_5_0__leaf_i_clk clknet_leaf_243_i_clk vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_25297_ _05965_ _06081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_69_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__26034__B _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15050_ rbzero.spi_registers.spi_cmd\[1\] _08827_ _08843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_27036_ _00946_ clknet_leaf_137_i_clk rbzero.tex_g0\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_24248_ net70 _05030_ _05018_ _05008_ _05031_ _05032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_181_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14353__A2 _08064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15955__I _09504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14001_ _07575_ _07811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_24179_ _04931_ _04843_ _04883_ _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_75_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__22966__A4 _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 net30 o_gpout[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_75_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput41 net41 o_tex_oeb0 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_246_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15302__A1 _07732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_18740_ _11699_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15952_ _09532_ _09533_ _09520_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_235_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14903_ rbzero.tex_b1\[54\] _08506_ _08709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_216_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18671_ rbzero.tex_r1\[8\] rbzero.tex_r1\[7\] _11656_ _11660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15883_ _09437_ _09480_ _08852_ _09481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_231_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15690__I _09336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_17622_ _10843_ _10844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14834_ _08636_ _08637_ _08639_ _08294_ _08509_ _08640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_230_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_17553_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _10802_ _10805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_106_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14765_ _08567_ _08569_ _08571_ _08284_ _08285_ _08572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_169_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16504_ _09951_ _09957_ _09958_ _09959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13716_ _07519_ _07521_ _07522_ _07525_ _07526_ _07527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_169_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_17484_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _10765_ _10766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14696_ _08495_ _08498_ _08501_ _08502_ _08346_ _08503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_19223_ rbzero.wall_tracer.mapY\[8\] _12062_ _12064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_16435_ _09892_ rbzero.pov.ss_buffer\[0\] _09894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13647_ rbzero.row_render.side _07458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14041__A1 _07848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_19154_ _11981_ _11983_ _11985_ _11997_ _11998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__20114__A1 _12471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13395__A3 _07205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14592__A2 _07843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_16366_ rbzero.spi_registers.buf_texadd3\[9\] _09840_ _09845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20114__B2 _12885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13578_ _07356_ _07387_ _07355_ _07389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_109_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_18105_ rbzero.map_rom.f1 _11249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_136_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15317_ rbzero.spi_registers.buf_mapdx\[3\] _09060_ _09061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_19085_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] _11929_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_147_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_16297_ _09746_ _09793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__22472__B _07160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_18036_ _11177_ _11178_ _11173_ _11179_ _11180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_151_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__19807__A1 rbzero.wall_tracer.size\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_200_Left_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14344__A2 _08006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15248_ _09007_ _09009_ _09003_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__20417__A2 _12644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15179_ _08949_ _08953_ _08954_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19987_ _12742_ _12749_ _12758_ _12759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_226_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13385__I gpout0.vpos\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_18938_ rbzero.tex_g0\[8\] rbzero.tex_g0\[7\] _11835_ _11839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
.ends

