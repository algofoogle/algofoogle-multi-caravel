magic
tech gf180mcuD
magscale 1 5
timestamp 1702222798
<< obsm1 >>
rect 672 1538 239288 20873
<< metal2 >>
rect 6384 21600 6440 22000
rect 7056 21600 7112 22000
rect 7728 21600 7784 22000
rect 8400 21600 8456 22000
rect 9072 21600 9128 22000
rect 9744 21600 9800 22000
rect 10416 21600 10472 22000
rect 11088 21600 11144 22000
rect 11760 21600 11816 22000
rect 12432 21600 12488 22000
rect 13104 21600 13160 22000
rect 13776 21600 13832 22000
rect 14448 21600 14504 22000
rect 15120 21600 15176 22000
rect 15792 21600 15848 22000
rect 16464 21600 16520 22000
rect 17136 21600 17192 22000
rect 17808 21600 17864 22000
rect 18480 21600 18536 22000
rect 19152 21600 19208 22000
rect 19824 21600 19880 22000
rect 20496 21600 20552 22000
rect 21168 21600 21224 22000
rect 21840 21600 21896 22000
rect 22512 21600 22568 22000
rect 23184 21600 23240 22000
rect 23856 21600 23912 22000
rect 24528 21600 24584 22000
rect 25200 21600 25256 22000
rect 25872 21600 25928 22000
rect 26544 21600 26600 22000
rect 27216 21600 27272 22000
rect 27888 21600 27944 22000
rect 28560 21600 28616 22000
rect 29232 21600 29288 22000
rect 29904 21600 29960 22000
rect 30576 21600 30632 22000
rect 31248 21600 31304 22000
rect 31920 21600 31976 22000
rect 32592 21600 32648 22000
rect 33264 21600 33320 22000
rect 33936 21600 33992 22000
rect 34608 21600 34664 22000
rect 35280 21600 35336 22000
rect 35952 21600 36008 22000
rect 36624 21600 36680 22000
rect 37296 21600 37352 22000
rect 37968 21600 38024 22000
rect 38640 21600 38696 22000
rect 39312 21600 39368 22000
rect 39984 21600 40040 22000
rect 40656 21600 40712 22000
rect 41328 21600 41384 22000
rect 42000 21600 42056 22000
rect 42672 21600 42728 22000
rect 43344 21600 43400 22000
rect 44016 21600 44072 22000
rect 44688 21600 44744 22000
rect 45360 21600 45416 22000
rect 46032 21600 46088 22000
rect 46704 21600 46760 22000
rect 47376 21600 47432 22000
rect 48048 21600 48104 22000
rect 48720 21600 48776 22000
rect 49392 21600 49448 22000
rect 50064 21600 50120 22000
rect 50736 21600 50792 22000
rect 51408 21600 51464 22000
rect 52080 21600 52136 22000
rect 59472 21600 59528 22000
rect 60144 21600 60200 22000
rect 60816 21600 60872 22000
rect 61488 21600 61544 22000
rect 62160 21600 62216 22000
rect 62832 21600 62888 22000
rect 63504 21600 63560 22000
rect 64176 21600 64232 22000
rect 64848 21600 64904 22000
rect 65520 21600 65576 22000
rect 66192 21600 66248 22000
rect 66864 21600 66920 22000
rect 74256 21600 74312 22000
rect 74928 21600 74984 22000
rect 75600 21600 75656 22000
rect 76272 21600 76328 22000
rect 76944 21600 77000 22000
rect 77616 21600 77672 22000
rect 78288 21600 78344 22000
rect 78960 21600 79016 22000
rect 79632 21600 79688 22000
rect 80304 21600 80360 22000
rect 80976 21600 81032 22000
rect 81648 21600 81704 22000
rect 82320 21600 82376 22000
rect 82992 21600 83048 22000
rect 83664 21600 83720 22000
rect 84336 21600 84392 22000
rect 85008 21600 85064 22000
rect 85680 21600 85736 22000
rect 86352 21600 86408 22000
rect 87024 21600 87080 22000
rect 87696 21600 87752 22000
rect 88368 21600 88424 22000
rect 89040 21600 89096 22000
rect 89712 21600 89768 22000
rect 90384 21600 90440 22000
rect 91056 21600 91112 22000
rect 91728 21600 91784 22000
rect 92400 21600 92456 22000
rect 93072 21600 93128 22000
rect 93744 21600 93800 22000
rect 94416 21600 94472 22000
rect 95088 21600 95144 22000
rect 95760 21600 95816 22000
rect 96432 21600 96488 22000
rect 97104 21600 97160 22000
rect 97776 21600 97832 22000
rect 98448 21600 98504 22000
rect 99120 21600 99176 22000
rect 99792 21600 99848 22000
rect 100464 21600 100520 22000
rect 101136 21600 101192 22000
rect 101808 21600 101864 22000
rect 102480 21600 102536 22000
rect 103152 21600 103208 22000
rect 103824 21600 103880 22000
rect 104496 21600 104552 22000
rect 105168 21600 105224 22000
rect 105840 21600 105896 22000
rect 106512 21600 106568 22000
rect 107184 21600 107240 22000
rect 107856 21600 107912 22000
rect 108528 21600 108584 22000
rect 109200 21600 109256 22000
rect 109872 21600 109928 22000
rect 110544 21600 110600 22000
rect 111216 21600 111272 22000
rect 111888 21600 111944 22000
rect 112560 21600 112616 22000
rect 113232 21600 113288 22000
rect 113904 21600 113960 22000
rect 114576 21600 114632 22000
rect 115248 21600 115304 22000
rect 115920 21600 115976 22000
rect 116592 21600 116648 22000
rect 117264 21600 117320 22000
rect 117936 21600 117992 22000
rect 118608 21600 118664 22000
rect 119280 21600 119336 22000
rect 119952 21600 120008 22000
rect 127344 21600 127400 22000
rect 128016 21600 128072 22000
rect 128688 21600 128744 22000
rect 129360 21600 129416 22000
rect 130032 21600 130088 22000
rect 130704 21600 130760 22000
rect 131376 21600 131432 22000
rect 132048 21600 132104 22000
rect 132720 21600 132776 22000
rect 140112 21600 140168 22000
rect 140784 21600 140840 22000
rect 141456 21600 141512 22000
rect 142128 21600 142184 22000
rect 142800 21600 142856 22000
rect 143472 21600 143528 22000
rect 144144 21600 144200 22000
rect 144816 21600 144872 22000
rect 145488 21600 145544 22000
rect 146160 21600 146216 22000
rect 146832 21600 146888 22000
rect 147504 21600 147560 22000
rect 148176 21600 148232 22000
rect 148848 21600 148904 22000
rect 149520 21600 149576 22000
rect 150192 21600 150248 22000
rect 150864 21600 150920 22000
rect 151536 21600 151592 22000
rect 152208 21600 152264 22000
rect 152880 21600 152936 22000
rect 153552 21600 153608 22000
rect 154224 21600 154280 22000
rect 154896 21600 154952 22000
rect 155568 21600 155624 22000
rect 156240 21600 156296 22000
rect 156912 21600 156968 22000
rect 157584 21600 157640 22000
rect 158256 21600 158312 22000
rect 158928 21600 158984 22000
rect 159600 21600 159656 22000
rect 160272 21600 160328 22000
rect 160944 21600 161000 22000
rect 161616 21600 161672 22000
rect 162288 21600 162344 22000
rect 162960 21600 163016 22000
rect 163632 21600 163688 22000
rect 164304 21600 164360 22000
rect 164976 21600 165032 22000
rect 165648 21600 165704 22000
rect 166320 21600 166376 22000
rect 166992 21600 167048 22000
rect 167664 21600 167720 22000
rect 168336 21600 168392 22000
rect 169008 21600 169064 22000
rect 169680 21600 169736 22000
rect 170352 21600 170408 22000
rect 171024 21600 171080 22000
rect 171696 21600 171752 22000
rect 172368 21600 172424 22000
rect 173040 21600 173096 22000
rect 173712 21600 173768 22000
rect 174384 21600 174440 22000
rect 175056 21600 175112 22000
rect 175728 21600 175784 22000
rect 176400 21600 176456 22000
rect 177072 21600 177128 22000
rect 177744 21600 177800 22000
rect 178416 21600 178472 22000
rect 179088 21600 179144 22000
rect 179760 21600 179816 22000
rect 180432 21600 180488 22000
rect 181104 21600 181160 22000
rect 181776 21600 181832 22000
rect 182448 21600 182504 22000
rect 183120 21600 183176 22000
rect 190512 21600 190568 22000
rect 191184 21600 191240 22000
rect 191856 21600 191912 22000
rect 192528 21600 192584 22000
rect 193200 21600 193256 22000
rect 193872 21600 193928 22000
rect 194544 21600 194600 22000
rect 195216 21600 195272 22000
rect 195888 21600 195944 22000
rect 196560 21600 196616 22000
rect 197232 21600 197288 22000
rect 197904 21600 197960 22000
rect 198576 21600 198632 22000
rect 199248 21600 199304 22000
rect 199920 21600 199976 22000
rect 200592 21600 200648 22000
rect 201264 21600 201320 22000
rect 201936 21600 201992 22000
rect 202608 21600 202664 22000
rect 203280 21600 203336 22000
rect 203952 21600 204008 22000
rect 204624 21600 204680 22000
rect 205296 21600 205352 22000
rect 205968 21600 206024 22000
rect 206640 21600 206696 22000
rect 207312 21600 207368 22000
rect 207984 21600 208040 22000
rect 208656 21600 208712 22000
rect 209328 21600 209384 22000
rect 210000 21600 210056 22000
rect 210672 21600 210728 22000
rect 211344 21600 211400 22000
rect 212016 21600 212072 22000
rect 212688 21600 212744 22000
rect 213360 21600 213416 22000
rect 214032 21600 214088 22000
rect 214704 21600 214760 22000
rect 215376 21600 215432 22000
rect 216048 21600 216104 22000
rect 216720 21600 216776 22000
rect 217392 21600 217448 22000
rect 218064 21600 218120 22000
rect 218736 21600 218792 22000
rect 219408 21600 219464 22000
rect 220080 21600 220136 22000
rect 220752 21600 220808 22000
rect 221424 21600 221480 22000
rect 222096 21600 222152 22000
rect 222768 21600 222824 22000
rect 223440 21600 223496 22000
rect 224112 21600 224168 22000
rect 224784 21600 224840 22000
rect 225456 21600 225512 22000
rect 226128 21600 226184 22000
rect 226800 21600 226856 22000
rect 5040 0 5096 400
rect 5712 0 5768 400
rect 6384 0 6440 400
rect 7056 0 7112 400
rect 7728 0 7784 400
rect 8400 0 8456 400
rect 9072 0 9128 400
rect 9744 0 9800 400
rect 10416 0 10472 400
rect 11088 0 11144 400
rect 11760 0 11816 400
rect 12432 0 12488 400
rect 13104 0 13160 400
rect 13776 0 13832 400
rect 14448 0 14504 400
rect 15120 0 15176 400
rect 15792 0 15848 400
rect 16464 0 16520 400
rect 17136 0 17192 400
rect 17808 0 17864 400
rect 18480 0 18536 400
rect 19152 0 19208 400
rect 19824 0 19880 400
rect 20496 0 20552 400
rect 21168 0 21224 400
rect 21840 0 21896 400
rect 22512 0 22568 400
rect 23184 0 23240 400
rect 23856 0 23912 400
rect 24528 0 24584 400
rect 25200 0 25256 400
rect 25872 0 25928 400
rect 26544 0 26600 400
rect 27216 0 27272 400
rect 27888 0 27944 400
rect 28560 0 28616 400
rect 29232 0 29288 400
rect 29904 0 29960 400
rect 30576 0 30632 400
rect 31248 0 31304 400
rect 31920 0 31976 400
rect 32592 0 32648 400
rect 33264 0 33320 400
rect 33936 0 33992 400
rect 34608 0 34664 400
rect 35280 0 35336 400
rect 35952 0 36008 400
rect 36624 0 36680 400
rect 37296 0 37352 400
rect 37968 0 38024 400
rect 38640 0 38696 400
rect 39312 0 39368 400
rect 39984 0 40040 400
rect 40656 0 40712 400
rect 41328 0 41384 400
rect 42000 0 42056 400
rect 42672 0 42728 400
rect 43344 0 43400 400
rect 44016 0 44072 400
rect 44688 0 44744 400
rect 45360 0 45416 400
rect 46032 0 46088 400
rect 46704 0 46760 400
rect 47376 0 47432 400
rect 48048 0 48104 400
rect 48720 0 48776 400
rect 49392 0 49448 400
rect 50064 0 50120 400
rect 50736 0 50792 400
rect 51408 0 51464 400
rect 52080 0 52136 400
rect 52752 0 52808 400
rect 53424 0 53480 400
rect 54096 0 54152 400
rect 54768 0 54824 400
rect 55440 0 55496 400
rect 56112 0 56168 400
rect 56784 0 56840 400
rect 57456 0 57512 400
rect 58128 0 58184 400
rect 58800 0 58856 400
rect 59472 0 59528 400
rect 60144 0 60200 400
rect 67536 0 67592 400
rect 68208 0 68264 400
rect 68880 0 68936 400
rect 69552 0 69608 400
rect 70224 0 70280 400
rect 70896 0 70952 400
rect 71568 0 71624 400
rect 72240 0 72296 400
rect 72912 0 72968 400
rect 73584 0 73640 400
rect 74256 0 74312 400
rect 74928 0 74984 400
rect 75600 0 75656 400
rect 76272 0 76328 400
rect 76944 0 77000 400
rect 77616 0 77672 400
rect 78288 0 78344 400
rect 78960 0 79016 400
rect 79632 0 79688 400
rect 80304 0 80360 400
rect 80976 0 81032 400
rect 81648 0 81704 400
rect 82320 0 82376 400
rect 82992 0 83048 400
rect 83664 0 83720 400
rect 84336 0 84392 400
rect 85008 0 85064 400
rect 85680 0 85736 400
rect 86352 0 86408 400
rect 87024 0 87080 400
rect 87696 0 87752 400
rect 88368 0 88424 400
rect 89040 0 89096 400
rect 89712 0 89768 400
rect 90384 0 90440 400
rect 91056 0 91112 400
rect 91728 0 91784 400
rect 92400 0 92456 400
rect 93072 0 93128 400
rect 93744 0 93800 400
rect 94416 0 94472 400
rect 95088 0 95144 400
rect 95760 0 95816 400
rect 96432 0 96488 400
rect 97104 0 97160 400
rect 97776 0 97832 400
rect 98448 0 98504 400
rect 99120 0 99176 400
rect 99792 0 99848 400
rect 100464 0 100520 400
rect 101136 0 101192 400
rect 101808 0 101864 400
rect 102480 0 102536 400
rect 103152 0 103208 400
rect 103824 0 103880 400
rect 104496 0 104552 400
rect 105168 0 105224 400
rect 105840 0 105896 400
rect 106512 0 106568 400
rect 107184 0 107240 400
rect 107856 0 107912 400
rect 108528 0 108584 400
rect 109200 0 109256 400
rect 109872 0 109928 400
rect 110544 0 110600 400
rect 111216 0 111272 400
rect 111888 0 111944 400
rect 112560 0 112616 400
rect 113232 0 113288 400
rect 113904 0 113960 400
rect 114576 0 114632 400
rect 115248 0 115304 400
rect 115920 0 115976 400
rect 116592 0 116648 400
rect 117264 0 117320 400
rect 117936 0 117992 400
rect 118608 0 118664 400
rect 119280 0 119336 400
rect 119952 0 120008 400
rect 127344 0 127400 400
rect 128016 0 128072 400
rect 128688 0 128744 400
rect 129360 0 129416 400
rect 130032 0 130088 400
rect 130704 0 130760 400
rect 131376 0 131432 400
rect 132048 0 132104 400
rect 132720 0 132776 400
rect 133392 0 133448 400
rect 134064 0 134120 400
rect 134736 0 134792 400
rect 135408 0 135464 400
rect 136080 0 136136 400
rect 136752 0 136808 400
rect 137424 0 137480 400
rect 151536 0 151592 400
rect 152208 0 152264 400
rect 152880 0 152936 400
rect 153552 0 153608 400
rect 154224 0 154280 400
rect 154896 0 154952 400
rect 155568 0 155624 400
rect 156240 0 156296 400
rect 156912 0 156968 400
rect 157584 0 157640 400
rect 158256 0 158312 400
rect 158928 0 158984 400
rect 159600 0 159656 400
rect 160272 0 160328 400
rect 160944 0 161000 400
rect 161616 0 161672 400
rect 162288 0 162344 400
rect 162960 0 163016 400
rect 163632 0 163688 400
rect 164304 0 164360 400
rect 164976 0 165032 400
rect 165648 0 165704 400
rect 166320 0 166376 400
rect 166992 0 167048 400
rect 167664 0 167720 400
rect 168336 0 168392 400
rect 169008 0 169064 400
rect 169680 0 169736 400
rect 170352 0 170408 400
rect 171024 0 171080 400
rect 171696 0 171752 400
rect 172368 0 172424 400
rect 173040 0 173096 400
rect 173712 0 173768 400
rect 174384 0 174440 400
rect 175056 0 175112 400
rect 175728 0 175784 400
rect 176400 0 176456 400
rect 177072 0 177128 400
rect 177744 0 177800 400
rect 178416 0 178472 400
rect 179088 0 179144 400
rect 179760 0 179816 400
rect 180432 0 180488 400
rect 181104 0 181160 400
rect 181776 0 181832 400
rect 182448 0 182504 400
rect 183120 0 183176 400
rect 183792 0 183848 400
rect 184464 0 184520 400
rect 185136 0 185192 400
rect 185808 0 185864 400
rect 186480 0 186536 400
rect 187152 0 187208 400
rect 187824 0 187880 400
rect 188496 0 188552 400
rect 189168 0 189224 400
rect 189840 0 189896 400
rect 190512 0 190568 400
rect 191184 0 191240 400
rect 191856 0 191912 400
rect 192528 0 192584 400
rect 193200 0 193256 400
rect 193872 0 193928 400
rect 194544 0 194600 400
rect 195216 0 195272 400
rect 195888 0 195944 400
rect 196560 0 196616 400
rect 197232 0 197288 400
rect 197904 0 197960 400
rect 198576 0 198632 400
rect 199248 0 199304 400
rect 199920 0 199976 400
rect 200592 0 200648 400
rect 201264 0 201320 400
rect 201936 0 201992 400
rect 202608 0 202664 400
rect 203280 0 203336 400
rect 203952 0 204008 400
rect 204624 0 204680 400
rect 205296 0 205352 400
rect 205968 0 206024 400
rect 206640 0 206696 400
rect 207312 0 207368 400
rect 207984 0 208040 400
rect 208656 0 208712 400
rect 209328 0 209384 400
rect 210000 0 210056 400
rect 210672 0 210728 400
rect 211344 0 211400 400
rect 212016 0 212072 400
rect 212688 0 212744 400
rect 213360 0 213416 400
rect 214032 0 214088 400
rect 214704 0 214760 400
rect 215376 0 215432 400
rect 216048 0 216104 400
rect 216720 0 216776 400
rect 217392 0 217448 400
rect 218064 0 218120 400
rect 218736 0 218792 400
rect 219408 0 219464 400
rect 220080 0 220136 400
rect 220752 0 220808 400
rect 221424 0 221480 400
<< obsm2 >>
rect 854 21570 6354 21658
rect 6470 21570 7026 21658
rect 7142 21570 7698 21658
rect 7814 21570 8370 21658
rect 8486 21570 9042 21658
rect 9158 21570 9714 21658
rect 9830 21570 10386 21658
rect 10502 21570 11058 21658
rect 11174 21570 11730 21658
rect 11846 21570 12402 21658
rect 12518 21570 13074 21658
rect 13190 21570 13746 21658
rect 13862 21570 14418 21658
rect 14534 21570 15090 21658
rect 15206 21570 15762 21658
rect 15878 21570 16434 21658
rect 16550 21570 17106 21658
rect 17222 21570 17778 21658
rect 17894 21570 18450 21658
rect 18566 21570 19122 21658
rect 19238 21570 19794 21658
rect 19910 21570 20466 21658
rect 20582 21570 21138 21658
rect 21254 21570 21810 21658
rect 21926 21570 22482 21658
rect 22598 21570 23154 21658
rect 23270 21570 23826 21658
rect 23942 21570 24498 21658
rect 24614 21570 25170 21658
rect 25286 21570 25842 21658
rect 25958 21570 26514 21658
rect 26630 21570 27186 21658
rect 27302 21570 27858 21658
rect 27974 21570 28530 21658
rect 28646 21570 29202 21658
rect 29318 21570 29874 21658
rect 29990 21570 30546 21658
rect 30662 21570 31218 21658
rect 31334 21570 31890 21658
rect 32006 21570 32562 21658
rect 32678 21570 33234 21658
rect 33350 21570 33906 21658
rect 34022 21570 34578 21658
rect 34694 21570 35250 21658
rect 35366 21570 35922 21658
rect 36038 21570 36594 21658
rect 36710 21570 37266 21658
rect 37382 21570 37938 21658
rect 38054 21570 38610 21658
rect 38726 21570 39282 21658
rect 39398 21570 39954 21658
rect 40070 21570 40626 21658
rect 40742 21570 41298 21658
rect 41414 21570 41970 21658
rect 42086 21570 42642 21658
rect 42758 21570 43314 21658
rect 43430 21570 43986 21658
rect 44102 21570 44658 21658
rect 44774 21570 45330 21658
rect 45446 21570 46002 21658
rect 46118 21570 46674 21658
rect 46790 21570 47346 21658
rect 47462 21570 48018 21658
rect 48134 21570 48690 21658
rect 48806 21570 49362 21658
rect 49478 21570 50034 21658
rect 50150 21570 50706 21658
rect 50822 21570 51378 21658
rect 51494 21570 52050 21658
rect 52166 21570 59442 21658
rect 59558 21570 60114 21658
rect 60230 21570 60786 21658
rect 60902 21570 61458 21658
rect 61574 21570 62130 21658
rect 62246 21570 62802 21658
rect 62918 21570 63474 21658
rect 63590 21570 64146 21658
rect 64262 21570 64818 21658
rect 64934 21570 65490 21658
rect 65606 21570 66162 21658
rect 66278 21570 66834 21658
rect 66950 21570 74226 21658
rect 74342 21570 74898 21658
rect 75014 21570 75570 21658
rect 75686 21570 76242 21658
rect 76358 21570 76914 21658
rect 77030 21570 77586 21658
rect 77702 21570 78258 21658
rect 78374 21570 78930 21658
rect 79046 21570 79602 21658
rect 79718 21570 80274 21658
rect 80390 21570 80946 21658
rect 81062 21570 81618 21658
rect 81734 21570 82290 21658
rect 82406 21570 82962 21658
rect 83078 21570 83634 21658
rect 83750 21570 84306 21658
rect 84422 21570 84978 21658
rect 85094 21570 85650 21658
rect 85766 21570 86322 21658
rect 86438 21570 86994 21658
rect 87110 21570 87666 21658
rect 87782 21570 88338 21658
rect 88454 21570 89010 21658
rect 89126 21570 89682 21658
rect 89798 21570 90354 21658
rect 90470 21570 91026 21658
rect 91142 21570 91698 21658
rect 91814 21570 92370 21658
rect 92486 21570 93042 21658
rect 93158 21570 93714 21658
rect 93830 21570 94386 21658
rect 94502 21570 95058 21658
rect 95174 21570 95730 21658
rect 95846 21570 96402 21658
rect 96518 21570 97074 21658
rect 97190 21570 97746 21658
rect 97862 21570 98418 21658
rect 98534 21570 99090 21658
rect 99206 21570 99762 21658
rect 99878 21570 100434 21658
rect 100550 21570 101106 21658
rect 101222 21570 101778 21658
rect 101894 21570 102450 21658
rect 102566 21570 103122 21658
rect 103238 21570 103794 21658
rect 103910 21570 104466 21658
rect 104582 21570 105138 21658
rect 105254 21570 105810 21658
rect 105926 21570 106482 21658
rect 106598 21570 107154 21658
rect 107270 21570 107826 21658
rect 107942 21570 108498 21658
rect 108614 21570 109170 21658
rect 109286 21570 109842 21658
rect 109958 21570 110514 21658
rect 110630 21570 111186 21658
rect 111302 21570 111858 21658
rect 111974 21570 112530 21658
rect 112646 21570 113202 21658
rect 113318 21570 113874 21658
rect 113990 21570 114546 21658
rect 114662 21570 115218 21658
rect 115334 21570 115890 21658
rect 116006 21570 116562 21658
rect 116678 21570 117234 21658
rect 117350 21570 117906 21658
rect 118022 21570 118578 21658
rect 118694 21570 119250 21658
rect 119366 21570 119922 21658
rect 120038 21570 127314 21658
rect 127430 21570 127986 21658
rect 128102 21570 128658 21658
rect 128774 21570 129330 21658
rect 129446 21570 130002 21658
rect 130118 21570 130674 21658
rect 130790 21570 131346 21658
rect 131462 21570 132018 21658
rect 132134 21570 132690 21658
rect 132806 21570 140082 21658
rect 140198 21570 140754 21658
rect 140870 21570 141426 21658
rect 141542 21570 142098 21658
rect 142214 21570 142770 21658
rect 142886 21570 143442 21658
rect 143558 21570 144114 21658
rect 144230 21570 144786 21658
rect 144902 21570 145458 21658
rect 145574 21570 146130 21658
rect 146246 21570 146802 21658
rect 146918 21570 147474 21658
rect 147590 21570 148146 21658
rect 148262 21570 148818 21658
rect 148934 21570 149490 21658
rect 149606 21570 150162 21658
rect 150278 21570 150834 21658
rect 150950 21570 151506 21658
rect 151622 21570 152178 21658
rect 152294 21570 152850 21658
rect 152966 21570 153522 21658
rect 153638 21570 154194 21658
rect 154310 21570 154866 21658
rect 154982 21570 155538 21658
rect 155654 21570 156210 21658
rect 156326 21570 156882 21658
rect 156998 21570 157554 21658
rect 157670 21570 158226 21658
rect 158342 21570 158898 21658
rect 159014 21570 159570 21658
rect 159686 21570 160242 21658
rect 160358 21570 160914 21658
rect 161030 21570 161586 21658
rect 161702 21570 162258 21658
rect 162374 21570 162930 21658
rect 163046 21570 163602 21658
rect 163718 21570 164274 21658
rect 164390 21570 164946 21658
rect 165062 21570 165618 21658
rect 165734 21570 166290 21658
rect 166406 21570 166962 21658
rect 167078 21570 167634 21658
rect 167750 21570 168306 21658
rect 168422 21570 168978 21658
rect 169094 21570 169650 21658
rect 169766 21570 170322 21658
rect 170438 21570 170994 21658
rect 171110 21570 171666 21658
rect 171782 21570 172338 21658
rect 172454 21570 173010 21658
rect 173126 21570 173682 21658
rect 173798 21570 174354 21658
rect 174470 21570 175026 21658
rect 175142 21570 175698 21658
rect 175814 21570 176370 21658
rect 176486 21570 177042 21658
rect 177158 21570 177714 21658
rect 177830 21570 178386 21658
rect 178502 21570 179058 21658
rect 179174 21570 179730 21658
rect 179846 21570 180402 21658
rect 180518 21570 181074 21658
rect 181190 21570 181746 21658
rect 181862 21570 182418 21658
rect 182534 21570 183090 21658
rect 183206 21570 190482 21658
rect 190598 21570 191154 21658
rect 191270 21570 191826 21658
rect 191942 21570 192498 21658
rect 192614 21570 193170 21658
rect 193286 21570 193842 21658
rect 193958 21570 194514 21658
rect 194630 21570 195186 21658
rect 195302 21570 195858 21658
rect 195974 21570 196530 21658
rect 196646 21570 197202 21658
rect 197318 21570 197874 21658
rect 197990 21570 198546 21658
rect 198662 21570 199218 21658
rect 199334 21570 199890 21658
rect 200006 21570 200562 21658
rect 200678 21570 201234 21658
rect 201350 21570 201906 21658
rect 202022 21570 202578 21658
rect 202694 21570 203250 21658
rect 203366 21570 203922 21658
rect 204038 21570 204594 21658
rect 204710 21570 205266 21658
rect 205382 21570 205938 21658
rect 206054 21570 206610 21658
rect 206726 21570 207282 21658
rect 207398 21570 207954 21658
rect 208070 21570 208626 21658
rect 208742 21570 209298 21658
rect 209414 21570 209970 21658
rect 210086 21570 210642 21658
rect 210758 21570 211314 21658
rect 211430 21570 211986 21658
rect 212102 21570 212658 21658
rect 212774 21570 213330 21658
rect 213446 21570 214002 21658
rect 214118 21570 214674 21658
rect 214790 21570 215346 21658
rect 215462 21570 216018 21658
rect 216134 21570 216690 21658
rect 216806 21570 217362 21658
rect 217478 21570 218034 21658
rect 218150 21570 218706 21658
rect 218822 21570 219378 21658
rect 219494 21570 220050 21658
rect 220166 21570 220722 21658
rect 220838 21570 221394 21658
rect 221510 21570 222066 21658
rect 222182 21570 222738 21658
rect 222854 21570 223410 21658
rect 223526 21570 224082 21658
rect 224198 21570 224754 21658
rect 224870 21570 225426 21658
rect 225542 21570 226098 21658
rect 226214 21570 226770 21658
rect 226886 21570 239162 21658
rect 854 430 239162 21570
rect 854 177 5010 430
rect 5126 177 5682 430
rect 5798 177 6354 430
rect 6470 177 7026 430
rect 7142 177 7698 430
rect 7814 177 8370 430
rect 8486 177 9042 430
rect 9158 177 9714 430
rect 9830 177 10386 430
rect 10502 177 11058 430
rect 11174 177 11730 430
rect 11846 177 12402 430
rect 12518 177 13074 430
rect 13190 177 13746 430
rect 13862 177 14418 430
rect 14534 177 15090 430
rect 15206 177 15762 430
rect 15878 177 16434 430
rect 16550 177 17106 430
rect 17222 177 17778 430
rect 17894 177 18450 430
rect 18566 177 19122 430
rect 19238 177 19794 430
rect 19910 177 20466 430
rect 20582 177 21138 430
rect 21254 177 21810 430
rect 21926 177 22482 430
rect 22598 177 23154 430
rect 23270 177 23826 430
rect 23942 177 24498 430
rect 24614 177 25170 430
rect 25286 177 25842 430
rect 25958 177 26514 430
rect 26630 177 27186 430
rect 27302 177 27858 430
rect 27974 177 28530 430
rect 28646 177 29202 430
rect 29318 177 29874 430
rect 29990 177 30546 430
rect 30662 177 31218 430
rect 31334 177 31890 430
rect 32006 177 32562 430
rect 32678 177 33234 430
rect 33350 177 33906 430
rect 34022 177 34578 430
rect 34694 177 35250 430
rect 35366 177 35922 430
rect 36038 177 36594 430
rect 36710 177 37266 430
rect 37382 177 37938 430
rect 38054 177 38610 430
rect 38726 177 39282 430
rect 39398 177 39954 430
rect 40070 177 40626 430
rect 40742 177 41298 430
rect 41414 177 41970 430
rect 42086 177 42642 430
rect 42758 177 43314 430
rect 43430 177 43986 430
rect 44102 177 44658 430
rect 44774 177 45330 430
rect 45446 177 46002 430
rect 46118 177 46674 430
rect 46790 177 47346 430
rect 47462 177 48018 430
rect 48134 177 48690 430
rect 48806 177 49362 430
rect 49478 177 50034 430
rect 50150 177 50706 430
rect 50822 177 51378 430
rect 51494 177 52050 430
rect 52166 177 52722 430
rect 52838 177 53394 430
rect 53510 177 54066 430
rect 54182 177 54738 430
rect 54854 177 55410 430
rect 55526 177 56082 430
rect 56198 177 56754 430
rect 56870 177 57426 430
rect 57542 177 58098 430
rect 58214 177 58770 430
rect 58886 177 59442 430
rect 59558 177 60114 430
rect 60230 177 67506 430
rect 67622 177 68178 430
rect 68294 177 68850 430
rect 68966 177 69522 430
rect 69638 177 70194 430
rect 70310 177 70866 430
rect 70982 177 71538 430
rect 71654 177 72210 430
rect 72326 177 72882 430
rect 72998 177 73554 430
rect 73670 177 74226 430
rect 74342 177 74898 430
rect 75014 177 75570 430
rect 75686 177 76242 430
rect 76358 177 76914 430
rect 77030 177 77586 430
rect 77702 177 78258 430
rect 78374 177 78930 430
rect 79046 177 79602 430
rect 79718 177 80274 430
rect 80390 177 80946 430
rect 81062 177 81618 430
rect 81734 177 82290 430
rect 82406 177 82962 430
rect 83078 177 83634 430
rect 83750 177 84306 430
rect 84422 177 84978 430
rect 85094 177 85650 430
rect 85766 177 86322 430
rect 86438 177 86994 430
rect 87110 177 87666 430
rect 87782 177 88338 430
rect 88454 177 89010 430
rect 89126 177 89682 430
rect 89798 177 90354 430
rect 90470 177 91026 430
rect 91142 177 91698 430
rect 91814 177 92370 430
rect 92486 177 93042 430
rect 93158 177 93714 430
rect 93830 177 94386 430
rect 94502 177 95058 430
rect 95174 177 95730 430
rect 95846 177 96402 430
rect 96518 177 97074 430
rect 97190 177 97746 430
rect 97862 177 98418 430
rect 98534 177 99090 430
rect 99206 177 99762 430
rect 99878 177 100434 430
rect 100550 177 101106 430
rect 101222 177 101778 430
rect 101894 177 102450 430
rect 102566 177 103122 430
rect 103238 177 103794 430
rect 103910 177 104466 430
rect 104582 177 105138 430
rect 105254 177 105810 430
rect 105926 177 106482 430
rect 106598 177 107154 430
rect 107270 177 107826 430
rect 107942 177 108498 430
rect 108614 177 109170 430
rect 109286 177 109842 430
rect 109958 177 110514 430
rect 110630 177 111186 430
rect 111302 177 111858 430
rect 111974 177 112530 430
rect 112646 177 113202 430
rect 113318 177 113874 430
rect 113990 177 114546 430
rect 114662 177 115218 430
rect 115334 177 115890 430
rect 116006 177 116562 430
rect 116678 177 117234 430
rect 117350 177 117906 430
rect 118022 177 118578 430
rect 118694 177 119250 430
rect 119366 177 119922 430
rect 120038 177 127314 430
rect 127430 177 127986 430
rect 128102 177 128658 430
rect 128774 177 129330 430
rect 129446 177 130002 430
rect 130118 177 130674 430
rect 130790 177 131346 430
rect 131462 177 132018 430
rect 132134 177 132690 430
rect 132806 177 133362 430
rect 133478 177 134034 430
rect 134150 177 134706 430
rect 134822 177 135378 430
rect 135494 177 136050 430
rect 136166 177 136722 430
rect 136838 177 137394 430
rect 137510 177 151506 430
rect 151622 177 152178 430
rect 152294 177 152850 430
rect 152966 177 153522 430
rect 153638 177 154194 430
rect 154310 177 154866 430
rect 154982 177 155538 430
rect 155654 177 156210 430
rect 156326 177 156882 430
rect 156998 177 157554 430
rect 157670 177 158226 430
rect 158342 177 158898 430
rect 159014 177 159570 430
rect 159686 177 160242 430
rect 160358 177 160914 430
rect 161030 177 161586 430
rect 161702 177 162258 430
rect 162374 177 162930 430
rect 163046 177 163602 430
rect 163718 177 164274 430
rect 164390 177 164946 430
rect 165062 177 165618 430
rect 165734 177 166290 430
rect 166406 177 166962 430
rect 167078 177 167634 430
rect 167750 177 168306 430
rect 168422 177 168978 430
rect 169094 177 169650 430
rect 169766 177 170322 430
rect 170438 177 170994 430
rect 171110 177 171666 430
rect 171782 177 172338 430
rect 172454 177 173010 430
rect 173126 177 173682 430
rect 173798 177 174354 430
rect 174470 177 175026 430
rect 175142 177 175698 430
rect 175814 177 176370 430
rect 176486 177 177042 430
rect 177158 177 177714 430
rect 177830 177 178386 430
rect 178502 177 179058 430
rect 179174 177 179730 430
rect 179846 177 180402 430
rect 180518 177 181074 430
rect 181190 177 181746 430
rect 181862 177 182418 430
rect 182534 177 183090 430
rect 183206 177 183762 430
rect 183878 177 184434 430
rect 184550 177 185106 430
rect 185222 177 185778 430
rect 185894 177 186450 430
rect 186566 177 187122 430
rect 187238 177 187794 430
rect 187910 177 188466 430
rect 188582 177 189138 430
rect 189254 177 189810 430
rect 189926 177 190482 430
rect 190598 177 191154 430
rect 191270 177 191826 430
rect 191942 177 192498 430
rect 192614 177 193170 430
rect 193286 177 193842 430
rect 193958 177 194514 430
rect 194630 177 195186 430
rect 195302 177 195858 430
rect 195974 177 196530 430
rect 196646 177 197202 430
rect 197318 177 197874 430
rect 197990 177 198546 430
rect 198662 177 199218 430
rect 199334 177 199890 430
rect 200006 177 200562 430
rect 200678 177 201234 430
rect 201350 177 201906 430
rect 202022 177 202578 430
rect 202694 177 203250 430
rect 203366 177 203922 430
rect 204038 177 204594 430
rect 204710 177 205266 430
rect 205382 177 205938 430
rect 206054 177 206610 430
rect 206726 177 207282 430
rect 207398 177 207954 430
rect 208070 177 208626 430
rect 208742 177 209298 430
rect 209414 177 209970 430
rect 210086 177 210642 430
rect 210758 177 211314 430
rect 211430 177 211986 430
rect 212102 177 212658 430
rect 212774 177 213330 430
rect 213446 177 214002 430
rect 214118 177 214674 430
rect 214790 177 215346 430
rect 215462 177 216018 430
rect 216134 177 216690 430
rect 216806 177 217362 430
rect 217478 177 218034 430
rect 218150 177 218706 430
rect 218822 177 219378 430
rect 219494 177 220050 430
rect 220166 177 220722 430
rect 220838 177 221394 430
rect 221510 177 239162 430
<< metal3 >>
rect 239600 21504 240000 21560
rect 0 21280 400 21336
rect 239600 21168 240000 21224
rect 0 20832 400 20888
rect 239600 20832 240000 20888
rect 239600 20496 240000 20552
rect 0 20384 400 20440
rect 239600 20160 240000 20216
rect 0 19936 400 19992
rect 239600 19824 240000 19880
rect 0 19488 400 19544
rect 239600 19488 240000 19544
rect 239600 19152 240000 19208
rect 0 19040 400 19096
rect 239600 18816 240000 18872
rect 0 18592 400 18648
rect 239600 18480 240000 18536
rect 0 18144 400 18200
rect 239600 18144 240000 18200
rect 239600 17808 240000 17864
rect 0 17696 400 17752
rect 239600 17472 240000 17528
rect 0 17248 400 17304
rect 239600 17136 240000 17192
rect 0 16800 400 16856
rect 239600 16800 240000 16856
rect 239600 16464 240000 16520
rect 0 16352 400 16408
rect 239600 16128 240000 16184
rect 0 15904 400 15960
rect 239600 15792 240000 15848
rect 0 15456 400 15512
rect 239600 15456 240000 15512
rect 239600 15120 240000 15176
rect 0 15008 400 15064
rect 239600 14784 240000 14840
rect 0 14560 400 14616
rect 239600 14448 240000 14504
rect 0 14112 400 14168
rect 239600 14112 240000 14168
rect 239600 13776 240000 13832
rect 0 13664 400 13720
rect 239600 13440 240000 13496
rect 0 13216 400 13272
rect 239600 13104 240000 13160
rect 0 12768 400 12824
rect 239600 12768 240000 12824
rect 239600 12432 240000 12488
rect 0 12320 400 12376
rect 239600 12096 240000 12152
rect 0 11872 400 11928
rect 239600 11760 240000 11816
rect 0 11424 400 11480
rect 239600 11424 240000 11480
rect 239600 11088 240000 11144
rect 0 10976 400 11032
rect 239600 10752 240000 10808
rect 0 10528 400 10584
rect 239600 10416 240000 10472
rect 0 10080 400 10136
rect 239600 10080 240000 10136
rect 239600 9744 240000 9800
rect 0 9632 400 9688
rect 239600 9408 240000 9464
rect 0 9184 400 9240
rect 239600 9072 240000 9128
rect 0 8736 400 8792
rect 239600 8736 240000 8792
rect 239600 8400 240000 8456
rect 0 8288 400 8344
rect 239600 8064 240000 8120
rect 0 7840 400 7896
rect 239600 7728 240000 7784
rect 0 7392 400 7448
rect 239600 7392 240000 7448
rect 239600 7056 240000 7112
rect 0 6944 400 7000
rect 239600 6720 240000 6776
rect 0 6496 400 6552
rect 239600 6384 240000 6440
rect 0 6048 400 6104
rect 239600 6048 240000 6104
rect 239600 5712 240000 5768
rect 0 5600 400 5656
rect 239600 5376 240000 5432
rect 0 5152 400 5208
rect 239600 5040 240000 5096
rect 0 4704 400 4760
rect 239600 4704 240000 4760
rect 239600 4368 240000 4424
rect 0 4256 400 4312
rect 239600 4032 240000 4088
rect 0 3808 400 3864
rect 239600 3696 240000 3752
rect 0 3360 400 3416
rect 239600 3360 240000 3416
rect 239600 3024 240000 3080
rect 0 2912 400 2968
rect 239600 2688 240000 2744
rect 0 2464 400 2520
rect 239600 2352 240000 2408
rect 0 2016 400 2072
rect 239600 2016 240000 2072
rect 239600 1680 240000 1736
rect 0 1568 400 1624
rect 239600 1344 240000 1400
rect 0 1120 400 1176
rect 239600 1008 240000 1064
rect 0 672 400 728
rect 239600 672 240000 728
rect 239600 336 240000 392
<< obsm3 >>
rect 400 21474 239570 21546
rect 400 21366 239600 21474
rect 430 21254 239600 21366
rect 430 21250 239570 21254
rect 400 21138 239570 21250
rect 400 20918 239600 21138
rect 430 20802 239570 20918
rect 400 20582 239600 20802
rect 400 20470 239570 20582
rect 430 20466 239570 20470
rect 430 20354 239600 20466
rect 400 20246 239600 20354
rect 400 20130 239570 20246
rect 400 20022 239600 20130
rect 430 19910 239600 20022
rect 430 19906 239570 19910
rect 400 19794 239570 19906
rect 400 19574 239600 19794
rect 430 19458 239570 19574
rect 400 19238 239600 19458
rect 400 19126 239570 19238
rect 430 19122 239570 19126
rect 430 19010 239600 19122
rect 400 18902 239600 19010
rect 400 18786 239570 18902
rect 400 18678 239600 18786
rect 430 18566 239600 18678
rect 430 18562 239570 18566
rect 400 18450 239570 18562
rect 400 18230 239600 18450
rect 430 18114 239570 18230
rect 400 17894 239600 18114
rect 400 17782 239570 17894
rect 430 17778 239570 17782
rect 430 17666 239600 17778
rect 400 17558 239600 17666
rect 400 17442 239570 17558
rect 400 17334 239600 17442
rect 430 17222 239600 17334
rect 430 17218 239570 17222
rect 400 17106 239570 17218
rect 400 16886 239600 17106
rect 430 16770 239570 16886
rect 400 16550 239600 16770
rect 400 16438 239570 16550
rect 430 16434 239570 16438
rect 430 16322 239600 16434
rect 400 16214 239600 16322
rect 400 16098 239570 16214
rect 400 15990 239600 16098
rect 430 15878 239600 15990
rect 430 15874 239570 15878
rect 400 15762 239570 15874
rect 400 15542 239600 15762
rect 430 15426 239570 15542
rect 400 15206 239600 15426
rect 400 15094 239570 15206
rect 430 15090 239570 15094
rect 430 14978 239600 15090
rect 400 14870 239600 14978
rect 400 14754 239570 14870
rect 400 14646 239600 14754
rect 430 14534 239600 14646
rect 430 14530 239570 14534
rect 400 14418 239570 14530
rect 400 14198 239600 14418
rect 430 14082 239570 14198
rect 400 13862 239600 14082
rect 400 13750 239570 13862
rect 430 13746 239570 13750
rect 430 13634 239600 13746
rect 400 13526 239600 13634
rect 400 13410 239570 13526
rect 400 13302 239600 13410
rect 430 13190 239600 13302
rect 430 13186 239570 13190
rect 400 13074 239570 13186
rect 400 12854 239600 13074
rect 430 12738 239570 12854
rect 400 12518 239600 12738
rect 400 12406 239570 12518
rect 430 12402 239570 12406
rect 430 12290 239600 12402
rect 400 12182 239600 12290
rect 400 12066 239570 12182
rect 400 11958 239600 12066
rect 430 11846 239600 11958
rect 430 11842 239570 11846
rect 400 11730 239570 11842
rect 400 11510 239600 11730
rect 430 11394 239570 11510
rect 400 11174 239600 11394
rect 400 11062 239570 11174
rect 430 11058 239570 11062
rect 430 10946 239600 11058
rect 400 10838 239600 10946
rect 400 10722 239570 10838
rect 400 10614 239600 10722
rect 430 10502 239600 10614
rect 430 10498 239570 10502
rect 400 10386 239570 10498
rect 400 10166 239600 10386
rect 430 10050 239570 10166
rect 400 9830 239600 10050
rect 400 9718 239570 9830
rect 430 9714 239570 9718
rect 430 9602 239600 9714
rect 400 9494 239600 9602
rect 400 9378 239570 9494
rect 400 9270 239600 9378
rect 430 9158 239600 9270
rect 430 9154 239570 9158
rect 400 9042 239570 9154
rect 400 8822 239600 9042
rect 430 8706 239570 8822
rect 400 8486 239600 8706
rect 400 8374 239570 8486
rect 430 8370 239570 8374
rect 430 8258 239600 8370
rect 400 8150 239600 8258
rect 400 8034 239570 8150
rect 400 7926 239600 8034
rect 430 7814 239600 7926
rect 430 7810 239570 7814
rect 400 7698 239570 7810
rect 400 7478 239600 7698
rect 430 7362 239570 7478
rect 400 7142 239600 7362
rect 400 7030 239570 7142
rect 430 7026 239570 7030
rect 430 6914 239600 7026
rect 400 6806 239600 6914
rect 400 6690 239570 6806
rect 400 6582 239600 6690
rect 430 6470 239600 6582
rect 430 6466 239570 6470
rect 400 6354 239570 6466
rect 400 6134 239600 6354
rect 430 6018 239570 6134
rect 400 5798 239600 6018
rect 400 5686 239570 5798
rect 430 5682 239570 5686
rect 430 5570 239600 5682
rect 400 5462 239600 5570
rect 400 5346 239570 5462
rect 400 5238 239600 5346
rect 430 5126 239600 5238
rect 430 5122 239570 5126
rect 400 5010 239570 5122
rect 400 4790 239600 5010
rect 430 4674 239570 4790
rect 400 4454 239600 4674
rect 400 4342 239570 4454
rect 430 4338 239570 4342
rect 430 4226 239600 4338
rect 400 4118 239600 4226
rect 400 4002 239570 4118
rect 400 3894 239600 4002
rect 430 3782 239600 3894
rect 430 3778 239570 3782
rect 400 3666 239570 3778
rect 400 3446 239600 3666
rect 430 3330 239570 3446
rect 400 3110 239600 3330
rect 400 2998 239570 3110
rect 430 2994 239570 2998
rect 430 2882 239600 2994
rect 400 2774 239600 2882
rect 400 2658 239570 2774
rect 400 2550 239600 2658
rect 430 2438 239600 2550
rect 430 2434 239570 2438
rect 400 2322 239570 2434
rect 400 2102 239600 2322
rect 430 1986 239570 2102
rect 400 1766 239600 1986
rect 400 1654 239570 1766
rect 430 1650 239570 1654
rect 430 1538 239600 1650
rect 400 1430 239600 1538
rect 400 1314 239570 1430
rect 400 1206 239600 1314
rect 430 1094 239600 1206
rect 430 1090 239570 1094
rect 400 978 239570 1090
rect 400 758 239600 978
rect 430 642 239570 758
rect 400 422 239600 642
rect 400 306 239570 422
rect 400 182 239600 306
<< metal4 >>
rect 2224 1538 2384 20414
rect 9904 1538 10064 20414
rect 17584 1538 17744 20414
rect 25264 1538 25424 20414
rect 32944 1538 33104 20414
rect 40624 1538 40784 20414
rect 48304 1538 48464 20414
rect 55984 1538 56144 20414
rect 63664 1538 63824 20414
rect 71344 1538 71504 20414
rect 79024 1538 79184 20414
rect 86704 1538 86864 20414
rect 94384 1538 94544 20414
rect 102064 1538 102224 20414
rect 109744 1538 109904 20414
rect 117424 1538 117584 20414
rect 125104 1538 125264 20414
rect 132784 1538 132944 20414
rect 140464 1538 140624 20414
rect 148144 1538 148304 20414
rect 155824 1538 155984 20414
rect 163504 1538 163664 20414
rect 171184 1538 171344 20414
rect 178864 1538 179024 20414
rect 186544 1538 186704 20414
rect 194224 1538 194384 20414
rect 201904 1538 202064 20414
rect 209584 1538 209744 20414
rect 217264 1538 217424 20414
rect 224944 1538 225104 20414
rect 232624 1538 232784 20414
<< obsm4 >>
rect 40950 1801 48274 20151
rect 48494 1801 55954 20151
rect 56174 1801 63634 20151
rect 63854 1801 71314 20151
rect 71534 1801 78994 20151
rect 79214 1801 86674 20151
rect 86894 1801 94354 20151
rect 94574 1801 102034 20151
rect 102254 1801 109714 20151
rect 109934 1801 117394 20151
rect 117614 1801 125074 20151
rect 125294 1801 132754 20151
rect 132974 1801 140434 20151
rect 140654 1801 148114 20151
rect 148334 1801 155794 20151
rect 156014 1801 160034 20151
<< labels >>
rlabel metal2 s 151536 0 151592 400 6 diego_clk
port 1 nsew signal output
rlabel metal2 s 152880 0 152936 400 6 diego_ena
port 2 nsew signal output
rlabel metal2 s 196560 0 196616 400 6 diego_io_in[0]
port 3 nsew signal output
rlabel metal2 s 203280 0 203336 400 6 diego_io_in[10]
port 4 nsew signal output
rlabel metal2 s 203952 0 204008 400 6 diego_io_in[11]
port 5 nsew signal output
rlabel metal2 s 204624 0 204680 400 6 diego_io_in[12]
port 6 nsew signal output
rlabel metal2 s 205296 0 205352 400 6 diego_io_in[13]
port 7 nsew signal output
rlabel metal2 s 205968 0 206024 400 6 diego_io_in[14]
port 8 nsew signal output
rlabel metal2 s 206640 0 206696 400 6 diego_io_in[15]
port 9 nsew signal output
rlabel metal2 s 207312 0 207368 400 6 diego_io_in[16]
port 10 nsew signal output
rlabel metal2 s 207984 0 208040 400 6 diego_io_in[17]
port 11 nsew signal output
rlabel metal2 s 208656 0 208712 400 6 diego_io_in[18]
port 12 nsew signal output
rlabel metal2 s 209328 0 209384 400 6 diego_io_in[19]
port 13 nsew signal output
rlabel metal2 s 197232 0 197288 400 6 diego_io_in[1]
port 14 nsew signal output
rlabel metal2 s 210000 0 210056 400 6 diego_io_in[20]
port 15 nsew signal output
rlabel metal2 s 210672 0 210728 400 6 diego_io_in[21]
port 16 nsew signal output
rlabel metal2 s 211344 0 211400 400 6 diego_io_in[22]
port 17 nsew signal output
rlabel metal2 s 212016 0 212072 400 6 diego_io_in[23]
port 18 nsew signal output
rlabel metal2 s 212688 0 212744 400 6 diego_io_in[24]
port 19 nsew signal output
rlabel metal2 s 213360 0 213416 400 6 diego_io_in[25]
port 20 nsew signal output
rlabel metal2 s 214032 0 214088 400 6 diego_io_in[26]
port 21 nsew signal output
rlabel metal2 s 214704 0 214760 400 6 diego_io_in[27]
port 22 nsew signal output
rlabel metal2 s 215376 0 215432 400 6 diego_io_in[28]
port 23 nsew signal output
rlabel metal2 s 216048 0 216104 400 6 diego_io_in[29]
port 24 nsew signal output
rlabel metal2 s 197904 0 197960 400 6 diego_io_in[2]
port 25 nsew signal output
rlabel metal2 s 216720 0 216776 400 6 diego_io_in[30]
port 26 nsew signal output
rlabel metal2 s 217392 0 217448 400 6 diego_io_in[31]
port 27 nsew signal output
rlabel metal2 s 218064 0 218120 400 6 diego_io_in[32]
port 28 nsew signal output
rlabel metal2 s 218736 0 218792 400 6 diego_io_in[33]
port 29 nsew signal output
rlabel metal2 s 219408 0 219464 400 6 diego_io_in[34]
port 30 nsew signal output
rlabel metal2 s 220080 0 220136 400 6 diego_io_in[35]
port 31 nsew signal output
rlabel metal2 s 220752 0 220808 400 6 diego_io_in[36]
port 32 nsew signal output
rlabel metal2 s 221424 0 221480 400 6 diego_io_in[37]
port 33 nsew signal output
rlabel metal2 s 198576 0 198632 400 6 diego_io_in[3]
port 34 nsew signal output
rlabel metal2 s 199248 0 199304 400 6 diego_io_in[4]
port 35 nsew signal output
rlabel metal2 s 199920 0 199976 400 6 diego_io_in[5]
port 36 nsew signal output
rlabel metal2 s 200592 0 200648 400 6 diego_io_in[6]
port 37 nsew signal output
rlabel metal2 s 201264 0 201320 400 6 diego_io_in[7]
port 38 nsew signal output
rlabel metal2 s 201936 0 201992 400 6 diego_io_in[8]
port 39 nsew signal output
rlabel metal2 s 202608 0 202664 400 6 diego_io_in[9]
port 40 nsew signal output
rlabel metal2 s 175056 0 175112 400 6 diego_io_oeb[0]
port 41 nsew signal input
rlabel metal2 s 181776 0 181832 400 6 diego_io_oeb[10]
port 42 nsew signal input
rlabel metal2 s 182448 0 182504 400 6 diego_io_oeb[11]
port 43 nsew signal input
rlabel metal2 s 183120 0 183176 400 6 diego_io_oeb[12]
port 44 nsew signal input
rlabel metal2 s 183792 0 183848 400 6 diego_io_oeb[13]
port 45 nsew signal input
rlabel metal2 s 184464 0 184520 400 6 diego_io_oeb[14]
port 46 nsew signal input
rlabel metal2 s 185136 0 185192 400 6 diego_io_oeb[15]
port 47 nsew signal input
rlabel metal2 s 185808 0 185864 400 6 diego_io_oeb[16]
port 48 nsew signal input
rlabel metal2 s 186480 0 186536 400 6 diego_io_oeb[17]
port 49 nsew signal input
rlabel metal2 s 187152 0 187208 400 6 diego_io_oeb[18]
port 50 nsew signal input
rlabel metal2 s 187824 0 187880 400 6 diego_io_oeb[19]
port 51 nsew signal input
rlabel metal2 s 175728 0 175784 400 6 diego_io_oeb[1]
port 52 nsew signal input
rlabel metal2 s 188496 0 188552 400 6 diego_io_oeb[20]
port 53 nsew signal input
rlabel metal2 s 189168 0 189224 400 6 diego_io_oeb[21]
port 54 nsew signal input
rlabel metal2 s 189840 0 189896 400 6 diego_io_oeb[22]
port 55 nsew signal input
rlabel metal2 s 190512 0 190568 400 6 diego_io_oeb[23]
port 56 nsew signal input
rlabel metal2 s 191184 0 191240 400 6 diego_io_oeb[24]
port 57 nsew signal input
rlabel metal2 s 191856 0 191912 400 6 diego_io_oeb[25]
port 58 nsew signal input
rlabel metal2 s 192528 0 192584 400 6 diego_io_oeb[26]
port 59 nsew signal input
rlabel metal2 s 193200 0 193256 400 6 diego_io_oeb[27]
port 60 nsew signal input
rlabel metal2 s 193872 0 193928 400 6 diego_io_oeb[28]
port 61 nsew signal input
rlabel metal2 s 194544 0 194600 400 6 diego_io_oeb[29]
port 62 nsew signal input
rlabel metal2 s 176400 0 176456 400 6 diego_io_oeb[2]
port 63 nsew signal input
rlabel metal2 s 195216 0 195272 400 6 diego_io_oeb[30]
port 64 nsew signal input
rlabel metal2 s 195888 0 195944 400 6 diego_io_oeb[31]
port 65 nsew signal input
rlabel metal2 s 177072 0 177128 400 6 diego_io_oeb[3]
port 66 nsew signal input
rlabel metal2 s 177744 0 177800 400 6 diego_io_oeb[4]
port 67 nsew signal input
rlabel metal2 s 178416 0 178472 400 6 diego_io_oeb[5]
port 68 nsew signal input
rlabel metal2 s 179088 0 179144 400 6 diego_io_oeb[6]
port 69 nsew signal input
rlabel metal2 s 179760 0 179816 400 6 diego_io_oeb[7]
port 70 nsew signal input
rlabel metal2 s 180432 0 180488 400 6 diego_io_oeb[8]
port 71 nsew signal input
rlabel metal2 s 181104 0 181160 400 6 diego_io_oeb[9]
port 72 nsew signal input
rlabel metal2 s 153552 0 153608 400 6 diego_io_out[0]
port 73 nsew signal input
rlabel metal2 s 160272 0 160328 400 6 diego_io_out[10]
port 74 nsew signal input
rlabel metal2 s 160944 0 161000 400 6 diego_io_out[11]
port 75 nsew signal input
rlabel metal2 s 161616 0 161672 400 6 diego_io_out[12]
port 76 nsew signal input
rlabel metal2 s 162288 0 162344 400 6 diego_io_out[13]
port 77 nsew signal input
rlabel metal2 s 162960 0 163016 400 6 diego_io_out[14]
port 78 nsew signal input
rlabel metal2 s 163632 0 163688 400 6 diego_io_out[15]
port 79 nsew signal input
rlabel metal2 s 164304 0 164360 400 6 diego_io_out[16]
port 80 nsew signal input
rlabel metal2 s 164976 0 165032 400 6 diego_io_out[17]
port 81 nsew signal input
rlabel metal2 s 165648 0 165704 400 6 diego_io_out[18]
port 82 nsew signal input
rlabel metal2 s 166320 0 166376 400 6 diego_io_out[19]
port 83 nsew signal input
rlabel metal2 s 154224 0 154280 400 6 diego_io_out[1]
port 84 nsew signal input
rlabel metal2 s 166992 0 167048 400 6 diego_io_out[20]
port 85 nsew signal input
rlabel metal2 s 167664 0 167720 400 6 diego_io_out[21]
port 86 nsew signal input
rlabel metal2 s 168336 0 168392 400 6 diego_io_out[22]
port 87 nsew signal input
rlabel metal2 s 169008 0 169064 400 6 diego_io_out[23]
port 88 nsew signal input
rlabel metal2 s 169680 0 169736 400 6 diego_io_out[24]
port 89 nsew signal input
rlabel metal2 s 170352 0 170408 400 6 diego_io_out[25]
port 90 nsew signal input
rlabel metal2 s 171024 0 171080 400 6 diego_io_out[26]
port 91 nsew signal input
rlabel metal2 s 171696 0 171752 400 6 diego_io_out[27]
port 92 nsew signal input
rlabel metal2 s 172368 0 172424 400 6 diego_io_out[28]
port 93 nsew signal input
rlabel metal2 s 173040 0 173096 400 6 diego_io_out[29]
port 94 nsew signal input
rlabel metal2 s 154896 0 154952 400 6 diego_io_out[2]
port 95 nsew signal input
rlabel metal2 s 173712 0 173768 400 6 diego_io_out[30]
port 96 nsew signal input
rlabel metal2 s 174384 0 174440 400 6 diego_io_out[31]
port 97 nsew signal input
rlabel metal2 s 155568 0 155624 400 6 diego_io_out[3]
port 98 nsew signal input
rlabel metal2 s 156240 0 156296 400 6 diego_io_out[4]
port 99 nsew signal input
rlabel metal2 s 156912 0 156968 400 6 diego_io_out[5]
port 100 nsew signal input
rlabel metal2 s 157584 0 157640 400 6 diego_io_out[6]
port 101 nsew signal input
rlabel metal2 s 158256 0 158312 400 6 diego_io_out[7]
port 102 nsew signal input
rlabel metal2 s 158928 0 158984 400 6 diego_io_out[8]
port 103 nsew signal input
rlabel metal2 s 159600 0 159656 400 6 diego_io_out[9]
port 104 nsew signal input
rlabel metal2 s 152208 0 152264 400 6 diego_rst
port 105 nsew signal output
rlabel metal3 s 239600 2688 240000 2744 6 i_design_reset[0]
port 106 nsew signal input
rlabel metal3 s 239600 3024 240000 3080 6 i_design_reset[1]
port 107 nsew signal input
rlabel metal3 s 239600 3360 240000 3416 6 i_design_reset[2]
port 108 nsew signal input
rlabel metal3 s 239600 3696 240000 3752 6 i_design_reset[3]
port 109 nsew signal input
rlabel metal3 s 239600 4032 240000 4088 6 i_design_reset[4]
port 110 nsew signal input
rlabel metal3 s 239600 4368 240000 4424 6 i_design_reset[5]
port 111 nsew signal input
rlabel metal3 s 239600 4704 240000 4760 6 i_design_reset[6]
port 112 nsew signal input
rlabel metal3 s 239600 5040 240000 5096 6 i_design_reset[7]
port 113 nsew signal input
rlabel metal3 s 239600 2352 240000 2408 6 i_mux_auto_reset_enb
port 114 nsew signal input
rlabel metal3 s 239600 336 240000 392 6 i_mux_io5_reset_enb
port 115 nsew signal input
rlabel metal3 s 239600 672 240000 728 6 i_mux_sel[0]
port 116 nsew signal input
rlabel metal3 s 239600 1008 240000 1064 6 i_mux_sel[1]
port 117 nsew signal input
rlabel metal3 s 239600 1344 240000 1400 6 i_mux_sel[2]
port 118 nsew signal input
rlabel metal3 s 239600 1680 240000 1736 6 i_mux_sel[3]
port 119 nsew signal input
rlabel metal3 s 239600 2016 240000 2072 6 i_mux_sys_reset_enb
port 120 nsew signal input
rlabel metal3 s 239600 5712 240000 5768 6 io_in[0]
port 121 nsew signal input
rlabel metal3 s 239600 15792 240000 15848 6 io_in[10]
port 122 nsew signal input
rlabel metal3 s 239600 16800 240000 16856 6 io_in[11]
port 123 nsew signal input
rlabel metal3 s 239600 17808 240000 17864 6 io_in[12]
port 124 nsew signal input
rlabel metal3 s 239600 18816 240000 18872 6 io_in[13]
port 125 nsew signal input
rlabel metal3 s 239600 19824 240000 19880 6 io_in[14]
port 126 nsew signal input
rlabel metal3 s 239600 20832 240000 20888 6 io_in[15]
port 127 nsew signal input
rlabel metal2 s 132720 21600 132776 22000 6 io_in[16]
port 128 nsew signal input
rlabel metal2 s 130704 21600 130760 22000 6 io_in[17]
port 129 nsew signal input
rlabel metal2 s 128688 21600 128744 22000 6 io_in[18]
port 130 nsew signal input
rlabel metal2 s 66864 21600 66920 22000 6 io_in[19]
port 131 nsew signal input
rlabel metal3 s 239600 6720 240000 6776 6 io_in[1]
port 132 nsew signal input
rlabel metal2 s 64848 21600 64904 22000 6 io_in[20]
port 133 nsew signal input
rlabel metal2 s 62832 21600 62888 22000 6 io_in[21]
port 134 nsew signal input
rlabel metal2 s 60816 21600 60872 22000 6 io_in[22]
port 135 nsew signal input
rlabel metal3 s 0 21280 400 21336 6 io_in[23]
port 136 nsew signal input
rlabel metal3 s 0 19936 400 19992 6 io_in[24]
port 137 nsew signal input
rlabel metal3 s 0 18592 400 18648 6 io_in[25]
port 138 nsew signal input
rlabel metal3 s 0 17248 400 17304 6 io_in[26]
port 139 nsew signal input
rlabel metal3 s 0 15904 400 15960 6 io_in[27]
port 140 nsew signal input
rlabel metal3 s 0 14560 400 14616 6 io_in[28]
port 141 nsew signal input
rlabel metal3 s 0 13216 400 13272 6 io_in[29]
port 142 nsew signal input
rlabel metal3 s 239600 7728 240000 7784 6 io_in[2]
port 143 nsew signal input
rlabel metal3 s 0 11872 400 11928 6 io_in[30]
port 144 nsew signal input
rlabel metal3 s 0 10528 400 10584 6 io_in[31]
port 145 nsew signal input
rlabel metal3 s 0 9184 400 9240 6 io_in[32]
port 146 nsew signal input
rlabel metal3 s 0 7840 400 7896 6 io_in[33]
port 147 nsew signal input
rlabel metal3 s 0 6496 400 6552 6 io_in[34]
port 148 nsew signal input
rlabel metal3 s 0 5152 400 5208 6 io_in[35]
port 149 nsew signal input
rlabel metal3 s 0 3808 400 3864 6 io_in[36]
port 150 nsew signal input
rlabel metal3 s 0 2464 400 2520 6 io_in[37]
port 151 nsew signal input
rlabel metal3 s 239600 8736 240000 8792 6 io_in[3]
port 152 nsew signal input
rlabel metal3 s 239600 9744 240000 9800 6 io_in[4]
port 153 nsew signal input
rlabel metal3 s 239600 10752 240000 10808 6 io_in[5]
port 154 nsew signal input
rlabel metal3 s 239600 11760 240000 11816 6 io_in[6]
port 155 nsew signal input
rlabel metal3 s 239600 12768 240000 12824 6 io_in[7]
port 156 nsew signal input
rlabel metal3 s 239600 13776 240000 13832 6 io_in[8]
port 157 nsew signal input
rlabel metal3 s 239600 14784 240000 14840 6 io_in[9]
port 158 nsew signal input
rlabel metal3 s 239600 6384 240000 6440 6 io_oeb[0]
port 159 nsew signal output
rlabel metal3 s 239600 16464 240000 16520 6 io_oeb[10]
port 160 nsew signal output
rlabel metal3 s 239600 17472 240000 17528 6 io_oeb[11]
port 161 nsew signal output
rlabel metal3 s 239600 18480 240000 18536 6 io_oeb[12]
port 162 nsew signal output
rlabel metal3 s 239600 19488 240000 19544 6 io_oeb[13]
port 163 nsew signal output
rlabel metal3 s 239600 20496 240000 20552 6 io_oeb[14]
port 164 nsew signal output
rlabel metal3 s 239600 21504 240000 21560 6 io_oeb[15]
port 165 nsew signal output
rlabel metal2 s 131376 21600 131432 22000 6 io_oeb[16]
port 166 nsew signal output
rlabel metal2 s 129360 21600 129416 22000 6 io_oeb[17]
port 167 nsew signal output
rlabel metal2 s 127344 21600 127400 22000 6 io_oeb[18]
port 168 nsew signal output
rlabel metal2 s 65520 21600 65576 22000 6 io_oeb[19]
port 169 nsew signal output
rlabel metal3 s 239600 7392 240000 7448 6 io_oeb[1]
port 170 nsew signal output
rlabel metal2 s 63504 21600 63560 22000 6 io_oeb[20]
port 171 nsew signal output
rlabel metal2 s 61488 21600 61544 22000 6 io_oeb[21]
port 172 nsew signal output
rlabel metal2 s 59472 21600 59528 22000 6 io_oeb[22]
port 173 nsew signal output
rlabel metal3 s 0 20384 400 20440 6 io_oeb[23]
port 174 nsew signal output
rlabel metal3 s 0 19040 400 19096 6 io_oeb[24]
port 175 nsew signal output
rlabel metal3 s 0 17696 400 17752 6 io_oeb[25]
port 176 nsew signal output
rlabel metal3 s 0 16352 400 16408 6 io_oeb[26]
port 177 nsew signal output
rlabel metal3 s 0 15008 400 15064 6 io_oeb[27]
port 178 nsew signal output
rlabel metal3 s 0 13664 400 13720 6 io_oeb[28]
port 179 nsew signal output
rlabel metal3 s 0 12320 400 12376 6 io_oeb[29]
port 180 nsew signal output
rlabel metal3 s 239600 8400 240000 8456 6 io_oeb[2]
port 181 nsew signal output
rlabel metal3 s 0 10976 400 11032 6 io_oeb[30]
port 182 nsew signal output
rlabel metal3 s 0 9632 400 9688 6 io_oeb[31]
port 183 nsew signal output
rlabel metal3 s 0 8288 400 8344 6 io_oeb[32]
port 184 nsew signal output
rlabel metal3 s 0 6944 400 7000 6 io_oeb[33]
port 185 nsew signal output
rlabel metal3 s 0 5600 400 5656 6 io_oeb[34]
port 186 nsew signal output
rlabel metal3 s 0 4256 400 4312 6 io_oeb[35]
port 187 nsew signal output
rlabel metal3 s 0 2912 400 2968 6 io_oeb[36]
port 188 nsew signal output
rlabel metal3 s 0 1568 400 1624 6 io_oeb[37]
port 189 nsew signal output
rlabel metal3 s 239600 9408 240000 9464 6 io_oeb[3]
port 190 nsew signal output
rlabel metal3 s 239600 10416 240000 10472 6 io_oeb[4]
port 191 nsew signal output
rlabel metal3 s 239600 11424 240000 11480 6 io_oeb[5]
port 192 nsew signal output
rlabel metal3 s 239600 12432 240000 12488 6 io_oeb[6]
port 193 nsew signal output
rlabel metal3 s 239600 13440 240000 13496 6 io_oeb[7]
port 194 nsew signal output
rlabel metal3 s 239600 14448 240000 14504 6 io_oeb[8]
port 195 nsew signal output
rlabel metal3 s 239600 15456 240000 15512 6 io_oeb[9]
port 196 nsew signal output
rlabel metal3 s 239600 6048 240000 6104 6 io_out[0]
port 197 nsew signal output
rlabel metal3 s 239600 16128 240000 16184 6 io_out[10]
port 198 nsew signal output
rlabel metal3 s 239600 17136 240000 17192 6 io_out[11]
port 199 nsew signal output
rlabel metal3 s 239600 18144 240000 18200 6 io_out[12]
port 200 nsew signal output
rlabel metal3 s 239600 19152 240000 19208 6 io_out[13]
port 201 nsew signal output
rlabel metal3 s 239600 20160 240000 20216 6 io_out[14]
port 202 nsew signal output
rlabel metal3 s 239600 21168 240000 21224 6 io_out[15]
port 203 nsew signal output
rlabel metal2 s 132048 21600 132104 22000 6 io_out[16]
port 204 nsew signal output
rlabel metal2 s 130032 21600 130088 22000 6 io_out[17]
port 205 nsew signal output
rlabel metal2 s 128016 21600 128072 22000 6 io_out[18]
port 206 nsew signal output
rlabel metal2 s 66192 21600 66248 22000 6 io_out[19]
port 207 nsew signal output
rlabel metal3 s 239600 7056 240000 7112 6 io_out[1]
port 208 nsew signal output
rlabel metal2 s 64176 21600 64232 22000 6 io_out[20]
port 209 nsew signal output
rlabel metal2 s 62160 21600 62216 22000 6 io_out[21]
port 210 nsew signal output
rlabel metal2 s 60144 21600 60200 22000 6 io_out[22]
port 211 nsew signal output
rlabel metal3 s 0 20832 400 20888 6 io_out[23]
port 212 nsew signal output
rlabel metal3 s 0 19488 400 19544 6 io_out[24]
port 213 nsew signal output
rlabel metal3 s 0 18144 400 18200 6 io_out[25]
port 214 nsew signal output
rlabel metal3 s 0 16800 400 16856 6 io_out[26]
port 215 nsew signal output
rlabel metal3 s 0 15456 400 15512 6 io_out[27]
port 216 nsew signal output
rlabel metal3 s 0 14112 400 14168 6 io_out[28]
port 217 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 io_out[29]
port 218 nsew signal output
rlabel metal3 s 239600 8064 240000 8120 6 io_out[2]
port 219 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 io_out[30]
port 220 nsew signal output
rlabel metal3 s 0 10080 400 10136 6 io_out[31]
port 221 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 io_out[32]
port 222 nsew signal output
rlabel metal3 s 0 7392 400 7448 6 io_out[33]
port 223 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 io_out[34]
port 224 nsew signal output
rlabel metal3 s 0 4704 400 4760 6 io_out[35]
port 225 nsew signal output
rlabel metal3 s 0 3360 400 3416 6 io_out[36]
port 226 nsew signal output
rlabel metal3 s 0 2016 400 2072 6 io_out[37]
port 227 nsew signal output
rlabel metal3 s 239600 9072 240000 9128 6 io_out[3]
port 228 nsew signal output
rlabel metal3 s 239600 10080 240000 10136 6 io_out[4]
port 229 nsew signal output
rlabel metal3 s 239600 11088 240000 11144 6 io_out[5]
port 230 nsew signal output
rlabel metal3 s 239600 12096 240000 12152 6 io_out[6]
port 231 nsew signal output
rlabel metal3 s 239600 13104 240000 13160 6 io_out[7]
port 232 nsew signal output
rlabel metal3 s 239600 14112 240000 14168 6 io_out[8]
port 233 nsew signal output
rlabel metal3 s 239600 15120 240000 15176 6 io_out[9]
port 234 nsew signal output
rlabel metal2 s 127344 0 127400 400 6 la_in[0]
port 235 nsew signal input
rlabel metal2 s 134064 0 134120 400 6 la_in[10]
port 236 nsew signal input
rlabel metal2 s 134736 0 134792 400 6 la_in[11]
port 237 nsew signal input
rlabel metal2 s 135408 0 135464 400 6 la_in[12]
port 238 nsew signal input
rlabel metal2 s 136080 0 136136 400 6 la_in[13]
port 239 nsew signal input
rlabel metal2 s 136752 0 136808 400 6 la_in[14]
port 240 nsew signal input
rlabel metal2 s 137424 0 137480 400 6 la_in[15]
port 241 nsew signal input
rlabel metal2 s 128016 0 128072 400 6 la_in[1]
port 242 nsew signal input
rlabel metal2 s 128688 0 128744 400 6 la_in[2]
port 243 nsew signal input
rlabel metal2 s 129360 0 129416 400 6 la_in[3]
port 244 nsew signal input
rlabel metal2 s 130032 0 130088 400 6 la_in[4]
port 245 nsew signal input
rlabel metal2 s 130704 0 130760 400 6 la_in[5]
port 246 nsew signal input
rlabel metal2 s 131376 0 131432 400 6 la_in[6]
port 247 nsew signal input
rlabel metal2 s 132048 0 132104 400 6 la_in[7]
port 248 nsew signal input
rlabel metal2 s 132720 0 132776 400 6 la_in[8]
port 249 nsew signal input
rlabel metal2 s 133392 0 133448 400 6 la_in[9]
port 250 nsew signal input
rlabel metal3 s 239600 5376 240000 5432 6 mux_conf_clk
port 251 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 pawel_clk
port 252 nsew signal output
rlabel metal2 s 6384 0 6440 400 6 pawel_ena
port 253 nsew signal output
rlabel metal2 s 35280 0 35336 400 6 pawel_io_in[0]
port 254 nsew signal output
rlabel metal2 s 42000 0 42056 400 6 pawel_io_in[10]
port 255 nsew signal output
rlabel metal2 s 42672 0 42728 400 6 pawel_io_in[11]
port 256 nsew signal output
rlabel metal2 s 43344 0 43400 400 6 pawel_io_in[12]
port 257 nsew signal output
rlabel metal2 s 44016 0 44072 400 6 pawel_io_in[13]
port 258 nsew signal output
rlabel metal2 s 44688 0 44744 400 6 pawel_io_in[14]
port 259 nsew signal output
rlabel metal2 s 45360 0 45416 400 6 pawel_io_in[15]
port 260 nsew signal output
rlabel metal2 s 46032 0 46088 400 6 pawel_io_in[16]
port 261 nsew signal output
rlabel metal2 s 46704 0 46760 400 6 pawel_io_in[17]
port 262 nsew signal output
rlabel metal2 s 47376 0 47432 400 6 pawel_io_in[18]
port 263 nsew signal output
rlabel metal2 s 48048 0 48104 400 6 pawel_io_in[19]
port 264 nsew signal output
rlabel metal2 s 35952 0 36008 400 6 pawel_io_in[1]
port 265 nsew signal output
rlabel metal2 s 48720 0 48776 400 6 pawel_io_in[20]
port 266 nsew signal output
rlabel metal2 s 49392 0 49448 400 6 pawel_io_in[21]
port 267 nsew signal output
rlabel metal2 s 50064 0 50120 400 6 pawel_io_in[22]
port 268 nsew signal output
rlabel metal2 s 50736 0 50792 400 6 pawel_io_in[23]
port 269 nsew signal output
rlabel metal2 s 51408 0 51464 400 6 pawel_io_in[24]
port 270 nsew signal output
rlabel metal2 s 52080 0 52136 400 6 pawel_io_in[25]
port 271 nsew signal output
rlabel metal2 s 52752 0 52808 400 6 pawel_io_in[26]
port 272 nsew signal output
rlabel metal2 s 53424 0 53480 400 6 pawel_io_in[27]
port 273 nsew signal output
rlabel metal2 s 54096 0 54152 400 6 pawel_io_in[28]
port 274 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 pawel_io_in[29]
port 275 nsew signal output
rlabel metal2 s 36624 0 36680 400 6 pawel_io_in[2]
port 276 nsew signal output
rlabel metal2 s 55440 0 55496 400 6 pawel_io_in[30]
port 277 nsew signal output
rlabel metal2 s 56112 0 56168 400 6 pawel_io_in[31]
port 278 nsew signal output
rlabel metal2 s 56784 0 56840 400 6 pawel_io_in[32]
port 279 nsew signal output
rlabel metal2 s 57456 0 57512 400 6 pawel_io_in[33]
port 280 nsew signal output
rlabel metal2 s 58128 0 58184 400 6 pawel_io_in[34]
port 281 nsew signal output
rlabel metal2 s 58800 0 58856 400 6 pawel_io_in[35]
port 282 nsew signal output
rlabel metal2 s 59472 0 59528 400 6 pawel_io_in[36]
port 283 nsew signal output
rlabel metal2 s 60144 0 60200 400 6 pawel_io_in[37]
port 284 nsew signal output
rlabel metal2 s 37296 0 37352 400 6 pawel_io_in[3]
port 285 nsew signal output
rlabel metal2 s 37968 0 38024 400 6 pawel_io_in[4]
port 286 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 pawel_io_in[5]
port 287 nsew signal output
rlabel metal2 s 39312 0 39368 400 6 pawel_io_in[6]
port 288 nsew signal output
rlabel metal2 s 39984 0 40040 400 6 pawel_io_in[7]
port 289 nsew signal output
rlabel metal2 s 40656 0 40712 400 6 pawel_io_in[8]
port 290 nsew signal output
rlabel metal2 s 41328 0 41384 400 6 pawel_io_in[9]
port 291 nsew signal output
rlabel metal2 s 15792 0 15848 400 6 pawel_io_oeb[0]
port 292 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 pawel_io_oeb[10]
port 293 nsew signal input
rlabel metal2 s 23184 0 23240 400 6 pawel_io_oeb[11]
port 294 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 pawel_io_oeb[12]
port 295 nsew signal input
rlabel metal2 s 16464 0 16520 400 6 pawel_io_oeb[1]
port 296 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 pawel_io_oeb[2]
port 297 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 pawel_io_oeb[3]
port 298 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 pawel_io_oeb[4]
port 299 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 pawel_io_oeb[5]
port 300 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 pawel_io_oeb[6]
port 301 nsew signal input
rlabel metal2 s 20496 0 20552 400 6 pawel_io_oeb[7]
port 302 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 pawel_io_oeb[8]
port 303 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 pawel_io_oeb[9]
port 304 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 pawel_io_out[0]
port 305 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 pawel_io_out[10]
port 306 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 pawel_io_out[11]
port 307 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 pawel_io_out[12]
port 308 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 pawel_io_out[1]
port 309 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 pawel_io_out[2]
port 310 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 pawel_io_out[3]
port 311 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 pawel_io_out[4]
port 312 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 pawel_io_out[5]
port 313 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 pawel_io_out[6]
port 314 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 pawel_io_out[7]
port 315 nsew signal input
rlabel metal2 s 12432 0 12488 400 6 pawel_io_out[8]
port 316 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 pawel_io_out[9]
port 317 nsew signal input
rlabel metal2 s 24528 0 24584 400 6 pawel_la_in[0]
port 318 nsew signal output
rlabel metal2 s 31248 0 31304 400 6 pawel_la_in[10]
port 319 nsew signal output
rlabel metal2 s 31920 0 31976 400 6 pawel_la_in[11]
port 320 nsew signal output
rlabel metal2 s 32592 0 32648 400 6 pawel_la_in[12]
port 321 nsew signal output
rlabel metal2 s 33264 0 33320 400 6 pawel_la_in[13]
port 322 nsew signal output
rlabel metal2 s 33936 0 33992 400 6 pawel_la_in[14]
port 323 nsew signal output
rlabel metal2 s 34608 0 34664 400 6 pawel_la_in[15]
port 324 nsew signal output
rlabel metal2 s 25200 0 25256 400 6 pawel_la_in[1]
port 325 nsew signal output
rlabel metal2 s 25872 0 25928 400 6 pawel_la_in[2]
port 326 nsew signal output
rlabel metal2 s 26544 0 26600 400 6 pawel_la_in[3]
port 327 nsew signal output
rlabel metal2 s 27216 0 27272 400 6 pawel_la_in[4]
port 328 nsew signal output
rlabel metal2 s 27888 0 27944 400 6 pawel_la_in[5]
port 329 nsew signal output
rlabel metal2 s 28560 0 28616 400 6 pawel_la_in[6]
port 330 nsew signal output
rlabel metal2 s 29232 0 29288 400 6 pawel_la_in[7]
port 331 nsew signal output
rlabel metal2 s 29904 0 29960 400 6 pawel_la_in[8]
port 332 nsew signal output
rlabel metal2 s 30576 0 30632 400 6 pawel_la_in[9]
port 333 nsew signal output
rlabel metal2 s 5712 0 5768 400 6 pawel_rst
port 334 nsew signal output
rlabel metal2 s 190512 21600 190568 22000 6 solos_clk
port 335 nsew signal output
rlabel metal2 s 191856 21600 191912 22000 6 solos_ena
port 336 nsew signal output
rlabel metal2 s 192528 21600 192584 22000 6 solos_gpio_ready
port 337 nsew signal output
rlabel metal2 s 218064 21600 218120 22000 6 solos_io_in[0]
port 338 nsew signal output
rlabel metal2 s 211344 21600 211400 22000 6 solos_io_in[10]
port 339 nsew signal output
rlabel metal2 s 210672 21600 210728 22000 6 solos_io_in[11]
port 340 nsew signal output
rlabel metal2 s 210000 21600 210056 22000 6 solos_io_in[12]
port 341 nsew signal output
rlabel metal2 s 209328 21600 209384 22000 6 solos_io_in[13]
port 342 nsew signal output
rlabel metal2 s 208656 21600 208712 22000 6 solos_io_in[14]
port 343 nsew signal output
rlabel metal2 s 207984 21600 208040 22000 6 solos_io_in[15]
port 344 nsew signal output
rlabel metal2 s 207312 21600 207368 22000 6 solos_io_in[16]
port 345 nsew signal output
rlabel metal2 s 206640 21600 206696 22000 6 solos_io_in[17]
port 346 nsew signal output
rlabel metal2 s 205968 21600 206024 22000 6 solos_io_in[18]
port 347 nsew signal output
rlabel metal2 s 205296 21600 205352 22000 6 solos_io_in[19]
port 348 nsew signal output
rlabel metal2 s 217392 21600 217448 22000 6 solos_io_in[1]
port 349 nsew signal output
rlabel metal2 s 204624 21600 204680 22000 6 solos_io_in[20]
port 350 nsew signal output
rlabel metal2 s 203952 21600 204008 22000 6 solos_io_in[21]
port 351 nsew signal output
rlabel metal2 s 203280 21600 203336 22000 6 solos_io_in[22]
port 352 nsew signal output
rlabel metal2 s 202608 21600 202664 22000 6 solos_io_in[23]
port 353 nsew signal output
rlabel metal2 s 201936 21600 201992 22000 6 solos_io_in[24]
port 354 nsew signal output
rlabel metal2 s 201264 21600 201320 22000 6 solos_io_in[25]
port 355 nsew signal output
rlabel metal2 s 200592 21600 200648 22000 6 solos_io_in[26]
port 356 nsew signal output
rlabel metal2 s 199920 21600 199976 22000 6 solos_io_in[27]
port 357 nsew signal output
rlabel metal2 s 199248 21600 199304 22000 6 solos_io_in[28]
port 358 nsew signal output
rlabel metal2 s 198576 21600 198632 22000 6 solos_io_in[29]
port 359 nsew signal output
rlabel metal2 s 216720 21600 216776 22000 6 solos_io_in[2]
port 360 nsew signal output
rlabel metal2 s 197904 21600 197960 22000 6 solos_io_in[30]
port 361 nsew signal output
rlabel metal2 s 197232 21600 197288 22000 6 solos_io_in[31]
port 362 nsew signal output
rlabel metal2 s 196560 21600 196616 22000 6 solos_io_in[32]
port 363 nsew signal output
rlabel metal2 s 195888 21600 195944 22000 6 solos_io_in[33]
port 364 nsew signal output
rlabel metal2 s 195216 21600 195272 22000 6 solos_io_in[34]
port 365 nsew signal output
rlabel metal2 s 194544 21600 194600 22000 6 solos_io_in[35]
port 366 nsew signal output
rlabel metal2 s 193872 21600 193928 22000 6 solos_io_in[36]
port 367 nsew signal output
rlabel metal2 s 193200 21600 193256 22000 6 solos_io_in[37]
port 368 nsew signal output
rlabel metal2 s 216048 21600 216104 22000 6 solos_io_in[3]
port 369 nsew signal output
rlabel metal2 s 215376 21600 215432 22000 6 solos_io_in[4]
port 370 nsew signal output
rlabel metal2 s 214704 21600 214760 22000 6 solos_io_in[5]
port 371 nsew signal output
rlabel metal2 s 214032 21600 214088 22000 6 solos_io_in[6]
port 372 nsew signal output
rlabel metal2 s 213360 21600 213416 22000 6 solos_io_in[7]
port 373 nsew signal output
rlabel metal2 s 212688 21600 212744 22000 6 solos_io_in[8]
port 374 nsew signal output
rlabel metal2 s 212016 21600 212072 22000 6 solos_io_in[9]
port 375 nsew signal output
rlabel metal2 s 226800 21600 226856 22000 6 solos_io_out[0]
port 376 nsew signal input
rlabel metal2 s 220080 21600 220136 22000 6 solos_io_out[10]
port 377 nsew signal input
rlabel metal2 s 219408 21600 219464 22000 6 solos_io_out[11]
port 378 nsew signal input
rlabel metal2 s 218736 21600 218792 22000 6 solos_io_out[12]
port 379 nsew signal input
rlabel metal2 s 226128 21600 226184 22000 6 solos_io_out[1]
port 380 nsew signal input
rlabel metal2 s 225456 21600 225512 22000 6 solos_io_out[2]
port 381 nsew signal input
rlabel metal2 s 224784 21600 224840 22000 6 solos_io_out[3]
port 382 nsew signal input
rlabel metal2 s 224112 21600 224168 22000 6 solos_io_out[4]
port 383 nsew signal input
rlabel metal2 s 223440 21600 223496 22000 6 solos_io_out[5]
port 384 nsew signal input
rlabel metal2 s 222768 21600 222824 22000 6 solos_io_out[6]
port 385 nsew signal input
rlabel metal2 s 222096 21600 222152 22000 6 solos_io_out[7]
port 386 nsew signal input
rlabel metal2 s 221424 21600 221480 22000 6 solos_io_out[8]
port 387 nsew signal input
rlabel metal2 s 220752 21600 220808 22000 6 solos_io_out[9]
port 388 nsew signal input
rlabel metal2 s 191184 21600 191240 22000 6 solos_rst
port 389 nsew signal output
rlabel metal2 s 74928 21600 74984 22000 6 trzf2_clk
port 390 nsew signal output
rlabel metal2 s 74256 21600 74312 22000 6 trzf2_ena
port 391 nsew signal output
rlabel metal2 s 119952 21600 120008 22000 6 trzf2_io_in[0]
port 392 nsew signal output
rlabel metal2 s 113232 21600 113288 22000 6 trzf2_io_in[10]
port 393 nsew signal output
rlabel metal2 s 112560 21600 112616 22000 6 trzf2_io_in[11]
port 394 nsew signal output
rlabel metal2 s 111888 21600 111944 22000 6 trzf2_io_in[12]
port 395 nsew signal output
rlabel metal2 s 111216 21600 111272 22000 6 trzf2_io_in[13]
port 396 nsew signal output
rlabel metal2 s 110544 21600 110600 22000 6 trzf2_io_in[14]
port 397 nsew signal output
rlabel metal2 s 109872 21600 109928 22000 6 trzf2_io_in[15]
port 398 nsew signal output
rlabel metal2 s 109200 21600 109256 22000 6 trzf2_io_in[16]
port 399 nsew signal output
rlabel metal2 s 108528 21600 108584 22000 6 trzf2_io_in[17]
port 400 nsew signal output
rlabel metal2 s 107856 21600 107912 22000 6 trzf2_io_in[18]
port 401 nsew signal output
rlabel metal2 s 107184 21600 107240 22000 6 trzf2_io_in[19]
port 402 nsew signal output
rlabel metal2 s 119280 21600 119336 22000 6 trzf2_io_in[1]
port 403 nsew signal output
rlabel metal2 s 106512 21600 106568 22000 6 trzf2_io_in[20]
port 404 nsew signal output
rlabel metal2 s 105840 21600 105896 22000 6 trzf2_io_in[21]
port 405 nsew signal output
rlabel metal2 s 105168 21600 105224 22000 6 trzf2_io_in[22]
port 406 nsew signal output
rlabel metal2 s 104496 21600 104552 22000 6 trzf2_io_in[23]
port 407 nsew signal output
rlabel metal2 s 103824 21600 103880 22000 6 trzf2_io_in[24]
port 408 nsew signal output
rlabel metal2 s 103152 21600 103208 22000 6 trzf2_io_in[25]
port 409 nsew signal output
rlabel metal2 s 102480 21600 102536 22000 6 trzf2_io_in[26]
port 410 nsew signal output
rlabel metal2 s 101808 21600 101864 22000 6 trzf2_io_in[27]
port 411 nsew signal output
rlabel metal2 s 101136 21600 101192 22000 6 trzf2_io_in[28]
port 412 nsew signal output
rlabel metal2 s 100464 21600 100520 22000 6 trzf2_io_in[29]
port 413 nsew signal output
rlabel metal2 s 118608 21600 118664 22000 6 trzf2_io_in[2]
port 414 nsew signal output
rlabel metal2 s 99792 21600 99848 22000 6 trzf2_io_in[30]
port 415 nsew signal output
rlabel metal2 s 99120 21600 99176 22000 6 trzf2_io_in[31]
port 416 nsew signal output
rlabel metal2 s 98448 21600 98504 22000 6 trzf2_io_in[32]
port 417 nsew signal output
rlabel metal2 s 97776 21600 97832 22000 6 trzf2_io_in[33]
port 418 nsew signal output
rlabel metal2 s 97104 21600 97160 22000 6 trzf2_io_in[34]
port 419 nsew signal output
rlabel metal2 s 96432 21600 96488 22000 6 trzf2_io_in[35]
port 420 nsew signal output
rlabel metal2 s 95760 21600 95816 22000 6 trzf2_io_in[36]
port 421 nsew signal output
rlabel metal2 s 95088 21600 95144 22000 6 trzf2_io_in[37]
port 422 nsew signal output
rlabel metal2 s 117936 21600 117992 22000 6 trzf2_io_in[3]
port 423 nsew signal output
rlabel metal2 s 117264 21600 117320 22000 6 trzf2_io_in[4]
port 424 nsew signal output
rlabel metal2 s 116592 21600 116648 22000 6 trzf2_io_in[5]
port 425 nsew signal output
rlabel metal2 s 115920 21600 115976 22000 6 trzf2_io_in[6]
port 426 nsew signal output
rlabel metal2 s 115248 21600 115304 22000 6 trzf2_io_in[7]
port 427 nsew signal output
rlabel metal2 s 114576 21600 114632 22000 6 trzf2_io_in[8]
port 428 nsew signal output
rlabel metal2 s 113904 21600 113960 22000 6 trzf2_io_in[9]
port 429 nsew signal output
rlabel metal2 s 84336 21600 84392 22000 6 trzf2_la_in[0]
port 430 nsew signal output
rlabel metal2 s 77616 21600 77672 22000 6 trzf2_la_in[10]
port 431 nsew signal output
rlabel metal2 s 76944 21600 77000 22000 6 trzf2_la_in[11]
port 432 nsew signal output
rlabel metal2 s 76272 21600 76328 22000 6 trzf2_la_in[12]
port 433 nsew signal output
rlabel metal2 s 83664 21600 83720 22000 6 trzf2_la_in[1]
port 434 nsew signal output
rlabel metal2 s 82992 21600 83048 22000 6 trzf2_la_in[2]
port 435 nsew signal output
rlabel metal2 s 82320 21600 82376 22000 6 trzf2_la_in[3]
port 436 nsew signal output
rlabel metal2 s 81648 21600 81704 22000 6 trzf2_la_in[4]
port 437 nsew signal output
rlabel metal2 s 80976 21600 81032 22000 6 trzf2_la_in[5]
port 438 nsew signal output
rlabel metal2 s 80304 21600 80360 22000 6 trzf2_la_in[6]
port 439 nsew signal output
rlabel metal2 s 79632 21600 79688 22000 6 trzf2_la_in[7]
port 440 nsew signal output
rlabel metal2 s 78960 21600 79016 22000 6 trzf2_la_in[8]
port 441 nsew signal output
rlabel metal2 s 78288 21600 78344 22000 6 trzf2_la_in[9]
port 442 nsew signal output
rlabel metal2 s 86352 21600 86408 22000 6 trzf2_o_gpout[0]
port 443 nsew signal input
rlabel metal2 s 85680 21600 85736 22000 6 trzf2_o_gpout[1]
port 444 nsew signal input
rlabel metal2 s 85008 21600 85064 22000 6 trzf2_o_gpout[2]
port 445 nsew signal input
rlabel metal2 s 94416 21600 94472 22000 6 trzf2_o_hsync
port 446 nsew signal input
rlabel metal2 s 93072 21600 93128 22000 6 trzf2_o_rgb[0]
port 447 nsew signal input
rlabel metal2 s 92400 21600 92456 22000 6 trzf2_o_rgb[1]
port 448 nsew signal input
rlabel metal2 s 91728 21600 91784 22000 6 trzf2_o_rgb[2]
port 449 nsew signal input
rlabel metal2 s 91056 21600 91112 22000 6 trzf2_o_rgb[3]
port 450 nsew signal input
rlabel metal2 s 90384 21600 90440 22000 6 trzf2_o_rgb[4]
port 451 nsew signal input
rlabel metal2 s 89712 21600 89768 22000 6 trzf2_o_rgb[5]
port 452 nsew signal input
rlabel metal2 s 89040 21600 89096 22000 6 trzf2_o_tex_csb
port 453 nsew signal input
rlabel metal2 s 87024 21600 87080 22000 6 trzf2_o_tex_oeb0
port 454 nsew signal input
rlabel metal2 s 87696 21600 87752 22000 6 trzf2_o_tex_out0
port 455 nsew signal input
rlabel metal2 s 88368 21600 88424 22000 6 trzf2_o_tex_sclk
port 456 nsew signal input
rlabel metal2 s 93744 21600 93800 22000 6 trzf2_o_vsync
port 457 nsew signal input
rlabel metal2 s 75600 21600 75656 22000 6 trzf2_rst
port 458 nsew signal output
rlabel metal2 s 7056 21600 7112 22000 6 trzf_clk
port 459 nsew signal output
rlabel metal2 s 6384 21600 6440 22000 6 trzf_ena
port 460 nsew signal output
rlabel metal2 s 52080 21600 52136 22000 6 trzf_io_in[0]
port 461 nsew signal output
rlabel metal2 s 45360 21600 45416 22000 6 trzf_io_in[10]
port 462 nsew signal output
rlabel metal2 s 44688 21600 44744 22000 6 trzf_io_in[11]
port 463 nsew signal output
rlabel metal2 s 44016 21600 44072 22000 6 trzf_io_in[12]
port 464 nsew signal output
rlabel metal2 s 43344 21600 43400 22000 6 trzf_io_in[13]
port 465 nsew signal output
rlabel metal2 s 42672 21600 42728 22000 6 trzf_io_in[14]
port 466 nsew signal output
rlabel metal2 s 42000 21600 42056 22000 6 trzf_io_in[15]
port 467 nsew signal output
rlabel metal2 s 41328 21600 41384 22000 6 trzf_io_in[16]
port 468 nsew signal output
rlabel metal2 s 40656 21600 40712 22000 6 trzf_io_in[17]
port 469 nsew signal output
rlabel metal2 s 39984 21600 40040 22000 6 trzf_io_in[18]
port 470 nsew signal output
rlabel metal2 s 39312 21600 39368 22000 6 trzf_io_in[19]
port 471 nsew signal output
rlabel metal2 s 51408 21600 51464 22000 6 trzf_io_in[1]
port 472 nsew signal output
rlabel metal2 s 38640 21600 38696 22000 6 trzf_io_in[20]
port 473 nsew signal output
rlabel metal2 s 37968 21600 38024 22000 6 trzf_io_in[21]
port 474 nsew signal output
rlabel metal2 s 37296 21600 37352 22000 6 trzf_io_in[22]
port 475 nsew signal output
rlabel metal2 s 36624 21600 36680 22000 6 trzf_io_in[23]
port 476 nsew signal output
rlabel metal2 s 35952 21600 36008 22000 6 trzf_io_in[24]
port 477 nsew signal output
rlabel metal2 s 35280 21600 35336 22000 6 trzf_io_in[25]
port 478 nsew signal output
rlabel metal2 s 34608 21600 34664 22000 6 trzf_io_in[26]
port 479 nsew signal output
rlabel metal2 s 33936 21600 33992 22000 6 trzf_io_in[27]
port 480 nsew signal output
rlabel metal2 s 33264 21600 33320 22000 6 trzf_io_in[28]
port 481 nsew signal output
rlabel metal2 s 32592 21600 32648 22000 6 trzf_io_in[29]
port 482 nsew signal output
rlabel metal2 s 50736 21600 50792 22000 6 trzf_io_in[2]
port 483 nsew signal output
rlabel metal2 s 31920 21600 31976 22000 6 trzf_io_in[30]
port 484 nsew signal output
rlabel metal2 s 31248 21600 31304 22000 6 trzf_io_in[31]
port 485 nsew signal output
rlabel metal2 s 30576 21600 30632 22000 6 trzf_io_in[32]
port 486 nsew signal output
rlabel metal2 s 29904 21600 29960 22000 6 trzf_io_in[33]
port 487 nsew signal output
rlabel metal2 s 29232 21600 29288 22000 6 trzf_io_in[34]
port 488 nsew signal output
rlabel metal2 s 28560 21600 28616 22000 6 trzf_io_in[35]
port 489 nsew signal output
rlabel metal2 s 27888 21600 27944 22000 6 trzf_io_in[36]
port 490 nsew signal output
rlabel metal2 s 27216 21600 27272 22000 6 trzf_io_in[37]
port 491 nsew signal output
rlabel metal2 s 50064 21600 50120 22000 6 trzf_io_in[3]
port 492 nsew signal output
rlabel metal2 s 49392 21600 49448 22000 6 trzf_io_in[4]
port 493 nsew signal output
rlabel metal2 s 48720 21600 48776 22000 6 trzf_io_in[5]
port 494 nsew signal output
rlabel metal2 s 48048 21600 48104 22000 6 trzf_io_in[6]
port 495 nsew signal output
rlabel metal2 s 47376 21600 47432 22000 6 trzf_io_in[7]
port 496 nsew signal output
rlabel metal2 s 46704 21600 46760 22000 6 trzf_io_in[8]
port 497 nsew signal output
rlabel metal2 s 46032 21600 46088 22000 6 trzf_io_in[9]
port 498 nsew signal output
rlabel metal2 s 16464 21600 16520 22000 6 trzf_la_in[0]
port 499 nsew signal output
rlabel metal2 s 9744 21600 9800 22000 6 trzf_la_in[10]
port 500 nsew signal output
rlabel metal2 s 9072 21600 9128 22000 6 trzf_la_in[11]
port 501 nsew signal output
rlabel metal2 s 8400 21600 8456 22000 6 trzf_la_in[12]
port 502 nsew signal output
rlabel metal2 s 15792 21600 15848 22000 6 trzf_la_in[1]
port 503 nsew signal output
rlabel metal2 s 15120 21600 15176 22000 6 trzf_la_in[2]
port 504 nsew signal output
rlabel metal2 s 14448 21600 14504 22000 6 trzf_la_in[3]
port 505 nsew signal output
rlabel metal2 s 13776 21600 13832 22000 6 trzf_la_in[4]
port 506 nsew signal output
rlabel metal2 s 13104 21600 13160 22000 6 trzf_la_in[5]
port 507 nsew signal output
rlabel metal2 s 12432 21600 12488 22000 6 trzf_la_in[6]
port 508 nsew signal output
rlabel metal2 s 11760 21600 11816 22000 6 trzf_la_in[7]
port 509 nsew signal output
rlabel metal2 s 11088 21600 11144 22000 6 trzf_la_in[8]
port 510 nsew signal output
rlabel metal2 s 10416 21600 10472 22000 6 trzf_la_in[9]
port 511 nsew signal output
rlabel metal2 s 18480 21600 18536 22000 6 trzf_o_gpout[0]
port 512 nsew signal input
rlabel metal2 s 17808 21600 17864 22000 6 trzf_o_gpout[1]
port 513 nsew signal input
rlabel metal2 s 17136 21600 17192 22000 6 trzf_o_gpout[2]
port 514 nsew signal input
rlabel metal2 s 26544 21600 26600 22000 6 trzf_o_hsync
port 515 nsew signal input
rlabel metal2 s 25200 21600 25256 22000 6 trzf_o_rgb[0]
port 516 nsew signal input
rlabel metal2 s 24528 21600 24584 22000 6 trzf_o_rgb[1]
port 517 nsew signal input
rlabel metal2 s 23856 21600 23912 22000 6 trzf_o_rgb[2]
port 518 nsew signal input
rlabel metal2 s 23184 21600 23240 22000 6 trzf_o_rgb[3]
port 519 nsew signal input
rlabel metal2 s 22512 21600 22568 22000 6 trzf_o_rgb[4]
port 520 nsew signal input
rlabel metal2 s 21840 21600 21896 22000 6 trzf_o_rgb[5]
port 521 nsew signal input
rlabel metal2 s 21168 21600 21224 22000 6 trzf_o_tex_csb
port 522 nsew signal input
rlabel metal2 s 19152 21600 19208 22000 6 trzf_o_tex_oeb0
port 523 nsew signal input
rlabel metal2 s 19824 21600 19880 22000 6 trzf_o_tex_out0
port 524 nsew signal input
rlabel metal2 s 20496 21600 20552 22000 6 trzf_o_tex_sclk
port 525 nsew signal input
rlabel metal2 s 25872 21600 25928 22000 6 trzf_o_vsync
port 526 nsew signal input
rlabel metal2 s 7728 21600 7784 22000 6 trzf_rst
port 527 nsew signal output
rlabel metal2 s 67536 0 67592 400 6 uri_clk
port 528 nsew signal output
rlabel metal2 s 68880 0 68936 400 6 uri_ena
port 529 nsew signal output
rlabel metal2 s 95088 0 95144 400 6 uri_io_in[0]
port 530 nsew signal output
rlabel metal2 s 101808 0 101864 400 6 uri_io_in[10]
port 531 nsew signal output
rlabel metal2 s 102480 0 102536 400 6 uri_io_in[11]
port 532 nsew signal output
rlabel metal2 s 103152 0 103208 400 6 uri_io_in[12]
port 533 nsew signal output
rlabel metal2 s 103824 0 103880 400 6 uri_io_in[13]
port 534 nsew signal output
rlabel metal2 s 104496 0 104552 400 6 uri_io_in[14]
port 535 nsew signal output
rlabel metal2 s 105168 0 105224 400 6 uri_io_in[15]
port 536 nsew signal output
rlabel metal2 s 105840 0 105896 400 6 uri_io_in[16]
port 537 nsew signal output
rlabel metal2 s 106512 0 106568 400 6 uri_io_in[17]
port 538 nsew signal output
rlabel metal2 s 107184 0 107240 400 6 uri_io_in[18]
port 539 nsew signal output
rlabel metal2 s 107856 0 107912 400 6 uri_io_in[19]
port 540 nsew signal output
rlabel metal2 s 95760 0 95816 400 6 uri_io_in[1]
port 541 nsew signal output
rlabel metal2 s 108528 0 108584 400 6 uri_io_in[20]
port 542 nsew signal output
rlabel metal2 s 109200 0 109256 400 6 uri_io_in[21]
port 543 nsew signal output
rlabel metal2 s 109872 0 109928 400 6 uri_io_in[22]
port 544 nsew signal output
rlabel metal2 s 110544 0 110600 400 6 uri_io_in[23]
port 545 nsew signal output
rlabel metal2 s 111216 0 111272 400 6 uri_io_in[24]
port 546 nsew signal output
rlabel metal2 s 111888 0 111944 400 6 uri_io_in[25]
port 547 nsew signal output
rlabel metal2 s 112560 0 112616 400 6 uri_io_in[26]
port 548 nsew signal output
rlabel metal2 s 113232 0 113288 400 6 uri_io_in[27]
port 549 nsew signal output
rlabel metal2 s 113904 0 113960 400 6 uri_io_in[28]
port 550 nsew signal output
rlabel metal2 s 114576 0 114632 400 6 uri_io_in[29]
port 551 nsew signal output
rlabel metal2 s 96432 0 96488 400 6 uri_io_in[2]
port 552 nsew signal output
rlabel metal2 s 115248 0 115304 400 6 uri_io_in[30]
port 553 nsew signal output
rlabel metal2 s 115920 0 115976 400 6 uri_io_in[31]
port 554 nsew signal output
rlabel metal2 s 116592 0 116648 400 6 uri_io_in[32]
port 555 nsew signal output
rlabel metal2 s 117264 0 117320 400 6 uri_io_in[33]
port 556 nsew signal output
rlabel metal2 s 117936 0 117992 400 6 uri_io_in[34]
port 557 nsew signal output
rlabel metal2 s 118608 0 118664 400 6 uri_io_in[35]
port 558 nsew signal output
rlabel metal2 s 119280 0 119336 400 6 uri_io_in[36]
port 559 nsew signal output
rlabel metal2 s 119952 0 120008 400 6 uri_io_in[37]
port 560 nsew signal output
rlabel metal2 s 97104 0 97160 400 6 uri_io_in[3]
port 561 nsew signal output
rlabel metal2 s 97776 0 97832 400 6 uri_io_in[4]
port 562 nsew signal output
rlabel metal2 s 98448 0 98504 400 6 uri_io_in[5]
port 563 nsew signal output
rlabel metal2 s 99120 0 99176 400 6 uri_io_in[6]
port 564 nsew signal output
rlabel metal2 s 99792 0 99848 400 6 uri_io_in[7]
port 565 nsew signal output
rlabel metal2 s 100464 0 100520 400 6 uri_io_in[8]
port 566 nsew signal output
rlabel metal2 s 101136 0 101192 400 6 uri_io_in[9]
port 567 nsew signal output
rlabel metal2 s 82320 0 82376 400 6 uri_io_oeb[0]
port 568 nsew signal input
rlabel metal2 s 89040 0 89096 400 6 uri_io_oeb[10]
port 569 nsew signal input
rlabel metal2 s 89712 0 89768 400 6 uri_io_oeb[11]
port 570 nsew signal input
rlabel metal2 s 90384 0 90440 400 6 uri_io_oeb[12]
port 571 nsew signal input
rlabel metal2 s 91056 0 91112 400 6 uri_io_oeb[13]
port 572 nsew signal input
rlabel metal2 s 91728 0 91784 400 6 uri_io_oeb[14]
port 573 nsew signal input
rlabel metal2 s 92400 0 92456 400 6 uri_io_oeb[15]
port 574 nsew signal input
rlabel metal2 s 93072 0 93128 400 6 uri_io_oeb[16]
port 575 nsew signal input
rlabel metal2 s 93744 0 93800 400 6 uri_io_oeb[17]
port 576 nsew signal input
rlabel metal2 s 94416 0 94472 400 6 uri_io_oeb[18]
port 577 nsew signal input
rlabel metal2 s 82992 0 83048 400 6 uri_io_oeb[1]
port 578 nsew signal input
rlabel metal2 s 83664 0 83720 400 6 uri_io_oeb[2]
port 579 nsew signal input
rlabel metal2 s 84336 0 84392 400 6 uri_io_oeb[3]
port 580 nsew signal input
rlabel metal2 s 85008 0 85064 400 6 uri_io_oeb[4]
port 581 nsew signal input
rlabel metal2 s 85680 0 85736 400 6 uri_io_oeb[5]
port 582 nsew signal input
rlabel metal2 s 86352 0 86408 400 6 uri_io_oeb[6]
port 583 nsew signal input
rlabel metal2 s 87024 0 87080 400 6 uri_io_oeb[7]
port 584 nsew signal input
rlabel metal2 s 87696 0 87752 400 6 uri_io_oeb[8]
port 585 nsew signal input
rlabel metal2 s 88368 0 88424 400 6 uri_io_oeb[9]
port 586 nsew signal input
rlabel metal2 s 69552 0 69608 400 6 uri_io_out[0]
port 587 nsew signal input
rlabel metal2 s 76272 0 76328 400 6 uri_io_out[10]
port 588 nsew signal input
rlabel metal2 s 76944 0 77000 400 6 uri_io_out[11]
port 589 nsew signal input
rlabel metal2 s 77616 0 77672 400 6 uri_io_out[12]
port 590 nsew signal input
rlabel metal2 s 78288 0 78344 400 6 uri_io_out[13]
port 591 nsew signal input
rlabel metal2 s 78960 0 79016 400 6 uri_io_out[14]
port 592 nsew signal input
rlabel metal2 s 79632 0 79688 400 6 uri_io_out[15]
port 593 nsew signal input
rlabel metal2 s 80304 0 80360 400 6 uri_io_out[16]
port 594 nsew signal input
rlabel metal2 s 80976 0 81032 400 6 uri_io_out[17]
port 595 nsew signal input
rlabel metal2 s 81648 0 81704 400 6 uri_io_out[18]
port 596 nsew signal input
rlabel metal2 s 70224 0 70280 400 6 uri_io_out[1]
port 597 nsew signal input
rlabel metal2 s 70896 0 70952 400 6 uri_io_out[2]
port 598 nsew signal input
rlabel metal2 s 71568 0 71624 400 6 uri_io_out[3]
port 599 nsew signal input
rlabel metal2 s 72240 0 72296 400 6 uri_io_out[4]
port 600 nsew signal input
rlabel metal2 s 72912 0 72968 400 6 uri_io_out[5]
port 601 nsew signal input
rlabel metal2 s 73584 0 73640 400 6 uri_io_out[6]
port 602 nsew signal input
rlabel metal2 s 74256 0 74312 400 6 uri_io_out[7]
port 603 nsew signal input
rlabel metal2 s 74928 0 74984 400 6 uri_io_out[8]
port 604 nsew signal input
rlabel metal2 s 75600 0 75656 400 6 uri_io_out[9]
port 605 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 uri_rst
port 606 nsew signal output
rlabel metal4 s 2224 1538 2384 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 20414 6 vdd
port 607 nsew power bidirectional
rlabel metal2 s 140112 21600 140168 22000 6 vgasp_clk
port 608 nsew signal output
rlabel metal2 s 141456 21600 141512 22000 6 vgasp_ena
port 609 nsew signal output
rlabel metal2 s 183120 21600 183176 22000 6 vgasp_io_in[0]
port 610 nsew signal output
rlabel metal2 s 176400 21600 176456 22000 6 vgasp_io_in[10]
port 611 nsew signal output
rlabel metal2 s 175728 21600 175784 22000 6 vgasp_io_in[11]
port 612 nsew signal output
rlabel metal2 s 175056 21600 175112 22000 6 vgasp_io_in[12]
port 613 nsew signal output
rlabel metal2 s 174384 21600 174440 22000 6 vgasp_io_in[13]
port 614 nsew signal output
rlabel metal2 s 173712 21600 173768 22000 6 vgasp_io_in[14]
port 615 nsew signal output
rlabel metal2 s 173040 21600 173096 22000 6 vgasp_io_in[15]
port 616 nsew signal output
rlabel metal2 s 172368 21600 172424 22000 6 vgasp_io_in[16]
port 617 nsew signal output
rlabel metal2 s 171696 21600 171752 22000 6 vgasp_io_in[17]
port 618 nsew signal output
rlabel metal2 s 171024 21600 171080 22000 6 vgasp_io_in[18]
port 619 nsew signal output
rlabel metal2 s 170352 21600 170408 22000 6 vgasp_io_in[19]
port 620 nsew signal output
rlabel metal2 s 182448 21600 182504 22000 6 vgasp_io_in[1]
port 621 nsew signal output
rlabel metal2 s 169680 21600 169736 22000 6 vgasp_io_in[20]
port 622 nsew signal output
rlabel metal2 s 169008 21600 169064 22000 6 vgasp_io_in[21]
port 623 nsew signal output
rlabel metal2 s 168336 21600 168392 22000 6 vgasp_io_in[22]
port 624 nsew signal output
rlabel metal2 s 167664 21600 167720 22000 6 vgasp_io_in[23]
port 625 nsew signal output
rlabel metal2 s 166992 21600 167048 22000 6 vgasp_io_in[24]
port 626 nsew signal output
rlabel metal2 s 166320 21600 166376 22000 6 vgasp_io_in[25]
port 627 nsew signal output
rlabel metal2 s 165648 21600 165704 22000 6 vgasp_io_in[26]
port 628 nsew signal output
rlabel metal2 s 164976 21600 165032 22000 6 vgasp_io_in[27]
port 629 nsew signal output
rlabel metal2 s 164304 21600 164360 22000 6 vgasp_io_in[28]
port 630 nsew signal output
rlabel metal2 s 163632 21600 163688 22000 6 vgasp_io_in[29]
port 631 nsew signal output
rlabel metal2 s 181776 21600 181832 22000 6 vgasp_io_in[2]
port 632 nsew signal output
rlabel metal2 s 162960 21600 163016 22000 6 vgasp_io_in[30]
port 633 nsew signal output
rlabel metal2 s 162288 21600 162344 22000 6 vgasp_io_in[31]
port 634 nsew signal output
rlabel metal2 s 161616 21600 161672 22000 6 vgasp_io_in[32]
port 635 nsew signal output
rlabel metal2 s 160944 21600 161000 22000 6 vgasp_io_in[33]
port 636 nsew signal output
rlabel metal2 s 160272 21600 160328 22000 6 vgasp_io_in[34]
port 637 nsew signal output
rlabel metal2 s 159600 21600 159656 22000 6 vgasp_io_in[35]
port 638 nsew signal output
rlabel metal2 s 158928 21600 158984 22000 6 vgasp_io_in[36]
port 639 nsew signal output
rlabel metal2 s 158256 21600 158312 22000 6 vgasp_io_in[37]
port 640 nsew signal output
rlabel metal2 s 181104 21600 181160 22000 6 vgasp_io_in[3]
port 641 nsew signal output
rlabel metal2 s 180432 21600 180488 22000 6 vgasp_io_in[4]
port 642 nsew signal output
rlabel metal2 s 179760 21600 179816 22000 6 vgasp_io_in[5]
port 643 nsew signal output
rlabel metal2 s 179088 21600 179144 22000 6 vgasp_io_in[6]
port 644 nsew signal output
rlabel metal2 s 178416 21600 178472 22000 6 vgasp_io_in[7]
port 645 nsew signal output
rlabel metal2 s 177744 21600 177800 22000 6 vgasp_io_in[8]
port 646 nsew signal output
rlabel metal2 s 177072 21600 177128 22000 6 vgasp_io_in[9]
port 647 nsew signal output
rlabel metal2 s 140784 21600 140840 22000 6 vgasp_rst
port 648 nsew signal output
rlabel metal2 s 146832 21600 146888 22000 6 vgasp_uio_oe[0]
port 649 nsew signal input
rlabel metal2 s 146160 21600 146216 22000 6 vgasp_uio_oe[1]
port 650 nsew signal input
rlabel metal2 s 145488 21600 145544 22000 6 vgasp_uio_oe[2]
port 651 nsew signal input
rlabel metal2 s 144816 21600 144872 22000 6 vgasp_uio_oe[3]
port 652 nsew signal input
rlabel metal2 s 144144 21600 144200 22000 6 vgasp_uio_oe[4]
port 653 nsew signal input
rlabel metal2 s 143472 21600 143528 22000 6 vgasp_uio_oe[5]
port 654 nsew signal input
rlabel metal2 s 142800 21600 142856 22000 6 vgasp_uio_oe[6]
port 655 nsew signal input
rlabel metal2 s 142128 21600 142184 22000 6 vgasp_uio_oe[7]
port 656 nsew signal input
rlabel metal2 s 152208 21600 152264 22000 6 vgasp_uio_out[0]
port 657 nsew signal input
rlabel metal2 s 151536 21600 151592 22000 6 vgasp_uio_out[1]
port 658 nsew signal input
rlabel metal2 s 150864 21600 150920 22000 6 vgasp_uio_out[2]
port 659 nsew signal input
rlabel metal2 s 150192 21600 150248 22000 6 vgasp_uio_out[3]
port 660 nsew signal input
rlabel metal2 s 149520 21600 149576 22000 6 vgasp_uio_out[4]
port 661 nsew signal input
rlabel metal2 s 148848 21600 148904 22000 6 vgasp_uio_out[5]
port 662 nsew signal input
rlabel metal2 s 148176 21600 148232 22000 6 vgasp_uio_out[6]
port 663 nsew signal input
rlabel metal2 s 147504 21600 147560 22000 6 vgasp_uio_out[7]
port 664 nsew signal input
rlabel metal2 s 157584 21600 157640 22000 6 vgasp_uo_out[0]
port 665 nsew signal input
rlabel metal2 s 156912 21600 156968 22000 6 vgasp_uo_out[1]
port 666 nsew signal input
rlabel metal2 s 156240 21600 156296 22000 6 vgasp_uo_out[2]
port 667 nsew signal input
rlabel metal2 s 155568 21600 155624 22000 6 vgasp_uo_out[3]
port 668 nsew signal input
rlabel metal2 s 154896 21600 154952 22000 6 vgasp_uo_out[4]
port 669 nsew signal input
rlabel metal2 s 154224 21600 154280 22000 6 vgasp_uo_out[5]
port 670 nsew signal input
rlabel metal2 s 153552 21600 153608 22000 6 vgasp_uo_out[6]
port 671 nsew signal input
rlabel metal2 s 152880 21600 152936 22000 6 vgasp_uo_out[7]
port 672 nsew signal input
rlabel metal4 s 9904 1538 10064 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 20414 6 vss
port 673 nsew ground bidirectional
rlabel metal3 s 0 1120 400 1176 6 wb_clk_i
port 674 nsew signal input
rlabel metal3 s 0 672 400 728 6 wb_rst_i
port 675 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 240000 22000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4189464
string GDS_FILE /home/zerotoasic/anton/algofoogle-multi-caravel/openlane/top_design_mux/runs/23_12_11_02_08/results/signoff/top_design_mux.magic.gds
string GDS_START 274270
<< end >>

