VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 1046.490 BY 1064.410 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 991.200 4.000 991.760 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 0.000 336.560 4.000 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 530.880 4.000 531.440 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.600 4.000 538.160 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 540.960 4.000 541.520 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 591.360 4.000 591.920 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 598.080 4.000 598.640 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 618.240 4.000 618.800 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 621.600 4.000 622.160 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 608.160 4.000 608.720 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 715.680 4.000 716.240 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 722.400 4.000 722.960 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 766.080 4.000 766.640 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 745.920 4.000 746.480 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 729.120 4.000 729.680 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 742.560 4.000 743.120 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 735.840 4.000 736.400 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 732.480 4.000 733.040 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 739.200 4.000 739.760 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 725.760 4.000 726.320 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 719.040 4.000 719.600 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 712.320 4.000 712.880 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 638.400 4.000 638.960 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 641.760 4.000 642.320 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 672.000 4.000 672.560 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 698.880 4.000 699.440 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 688.800 4.000 689.360 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 682.080 4.000 682.640 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 692.160 4.000 692.720 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 678.720 4.000 679.280 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 685.440 4.000 686.000 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 661.920 4.000 662.480 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 665.280 4.000 665.840 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 668.640 4.000 669.200 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 564.480 4.000 565.040 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.920 4.000 578.480 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.120 4.000 561.680 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.400 4.000 554.960 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 594.720 4.000 595.280 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 581.280 4.000 581.840 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 0.000 282.800 4.000 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 1060.410 645.680 1064.410 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 749.280 4.000 749.840 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 702.240 4.000 702.800 ;
    END
  END i_reg_mosi
  PIN i_reg_outs_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 584.640 4.000 585.200 ;
    END
  END i_reg_outs_enb
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 762.720 4.000 763.280 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 551.040 4.000 551.600 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 571.200 4.000 571.760 ;
    END
  END i_reset_lock_b
  PIN i_spare_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END i_spare_0
  PIN i_spare_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END i_spare_1
  PIN i_test_uc2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 759.360 4.000 759.920 ;
    END
  END i_test_uc2
  PIN i_test_wci
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 756.000 4.000 756.560 ;
    END
  END i_test_wci
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 604.800 4.000 605.360 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 601.440 4.000 602.000 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 705.600 4.000 706.160 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 628.320 4.000 628.880 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 624.960 4.000 625.520 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 752.640 4.000 753.200 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.040 4.000 635.600 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.320 4.000 544.880 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 611.520 4.000 612.080 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 708.960 4.000 709.520 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 675.360 4.000 675.920 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 695.520 4.000 696.080 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 547.680 4.000 548.240 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 567.840 4.000 568.400 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 527.520 4.000 528.080 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 0.000 450.800 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 0.000 672.560 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 833.280 1060.410 833.840 1064.410 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 0.000 948.080 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 1060.410 773.360 1064.410 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.120 4.000 645.680 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 0.000 985.040 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 0.000 427.280 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 1060.410 904.400 1064.410 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 0.000 551.600 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1042.490 971.040 1046.490 971.600 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1042.490 1031.520 1046.490 1032.080 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 913.920 0.000 914.480 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 655.200 4.000 655.760 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 588.000 4.000 588.560 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1042.490 1038.240 1046.490 1038.800 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 1060.410 14.000 1064.410 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1031.520 0.000 1032.080 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 13.440 4.000 14.000 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 631.680 4.000 632.240 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.880 4.000 615.440 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 4.000 17.360 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1008.000 0.000 1008.560 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.240 4.000 534.800 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 658.560 4.000 659.120 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 648.480 4.000 649.040 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 651.840 4.000 652.400 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 557.760 4.000 558.320 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 1060.410 145.040 1064.410 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 1060.410 739.760 1064.410 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 860.160 0.000 860.720 4.000 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 977.760 0.000 978.320 4.000 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 4.000 24.080 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1042.490 1044.960 1046.490 1045.520 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 4.000 27.440 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 0.000 981.680 4.000 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 1060.410 155.120 1064.410 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 1060.410 686.000 1064.410 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1042.490 1041.600 1046.490 1042.160 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 4.000 30.800 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 0.000 507.920 4.000 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 0.000 296.240 4.000 ;
    END
  END ones[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1046.940 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1046.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1046.940 ;
    END
  END vss
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1042.490 1034.880 1046.490 1035.440 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1011.360 0.000 1011.920 4.000 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 1060.410 743.120 1064.410 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 1060.410 854.000 1064.410 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 1060.410 638.960 1064.410 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 0.000 460.880 4.000 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 887.040 1060.410 887.600 1064.410 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 1060.410 890.960 1064.410 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 1060.410 360.080 1064.410 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 0.000 319.760 4.000 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 0.000 470.960 4.000 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 806.400 1060.410 806.960 1064.410 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 1060.410 800.240 1064.410 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 1060.410 790.160 1064.410 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1014.720 0.000 1015.280 4.000 ;
    END
  END zeros[9]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1039.360 1046.940 ;
      LAYER Metal2 ;
        RECT 7.420 1060.110 13.140 1060.410 ;
        RECT 14.300 1060.110 144.180 1060.410 ;
        RECT 145.340 1060.110 154.260 1060.410 ;
        RECT 155.420 1060.110 359.220 1060.410 ;
        RECT 360.380 1060.110 638.100 1060.410 ;
        RECT 639.260 1060.110 644.820 1060.410 ;
        RECT 645.980 1060.110 685.140 1060.410 ;
        RECT 686.300 1060.110 738.900 1060.410 ;
        RECT 740.060 1060.110 742.260 1060.410 ;
        RECT 743.420 1060.110 772.500 1060.410 ;
        RECT 773.660 1060.110 789.300 1060.410 ;
        RECT 790.460 1060.110 799.380 1060.410 ;
        RECT 800.540 1060.110 806.100 1060.410 ;
        RECT 807.260 1060.110 832.980 1060.410 ;
        RECT 834.140 1060.110 853.140 1060.410 ;
        RECT 854.300 1060.110 886.740 1060.410 ;
        RECT 887.900 1060.110 890.100 1060.410 ;
        RECT 891.260 1060.110 903.540 1060.410 ;
        RECT 904.700 1060.110 1038.100 1060.410 ;
        RECT 7.420 4.300 1038.100 1060.110 ;
        RECT 7.580 4.000 164.340 4.300 ;
        RECT 165.500 4.000 255.060 4.300 ;
        RECT 256.220 4.000 281.940 4.300 ;
        RECT 283.100 4.000 285.300 4.300 ;
        RECT 286.460 4.000 295.380 4.300 ;
        RECT 296.540 4.000 318.900 4.300 ;
        RECT 320.060 4.000 335.700 4.300 ;
        RECT 336.860 4.000 426.420 4.300 ;
        RECT 427.580 4.000 449.940 4.300 ;
        RECT 451.100 4.000 460.020 4.300 ;
        RECT 461.180 4.000 470.100 4.300 ;
        RECT 471.260 4.000 507.060 4.300 ;
        RECT 508.220 4.000 550.740 4.300 ;
        RECT 551.900 4.000 671.700 4.300 ;
        RECT 672.860 4.000 859.860 4.300 ;
        RECT 861.020 4.000 913.620 4.300 ;
        RECT 914.780 4.000 947.220 4.300 ;
        RECT 948.380 4.000 977.460 4.300 ;
        RECT 978.620 4.000 980.820 4.300 ;
        RECT 981.980 4.000 984.180 4.300 ;
        RECT 985.340 4.000 1007.700 4.300 ;
        RECT 1008.860 4.000 1011.060 4.300 ;
        RECT 1012.220 4.000 1014.420 4.300 ;
        RECT 1015.580 4.000 1031.220 4.300 ;
        RECT 1032.380 4.000 1038.100 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1045.820 1042.490 1046.780 ;
        RECT 4.000 1044.660 1042.190 1045.820 ;
        RECT 4.000 1042.460 1042.490 1044.660 ;
        RECT 4.000 1041.300 1042.190 1042.460 ;
        RECT 4.000 1039.100 1042.490 1041.300 ;
        RECT 4.000 1037.940 1042.190 1039.100 ;
        RECT 4.000 1035.740 1042.490 1037.940 ;
        RECT 4.000 1034.580 1042.190 1035.740 ;
        RECT 4.000 1032.380 1042.490 1034.580 ;
        RECT 4.000 1031.220 1042.190 1032.380 ;
        RECT 4.000 992.060 1042.490 1031.220 ;
        RECT 4.300 990.900 1042.490 992.060 ;
        RECT 4.000 971.900 1042.490 990.900 ;
        RECT 4.000 970.740 1042.190 971.900 ;
        RECT 4.000 766.940 1042.490 970.740 ;
        RECT 4.300 765.780 1042.490 766.940 ;
        RECT 4.000 763.580 1042.490 765.780 ;
        RECT 4.300 762.420 1042.490 763.580 ;
        RECT 4.000 760.220 1042.490 762.420 ;
        RECT 4.300 759.060 1042.490 760.220 ;
        RECT 4.000 756.860 1042.490 759.060 ;
        RECT 4.300 755.700 1042.490 756.860 ;
        RECT 4.000 753.500 1042.490 755.700 ;
        RECT 4.300 752.340 1042.490 753.500 ;
        RECT 4.000 750.140 1042.490 752.340 ;
        RECT 4.300 748.980 1042.490 750.140 ;
        RECT 4.000 746.780 1042.490 748.980 ;
        RECT 4.300 745.620 1042.490 746.780 ;
        RECT 4.000 743.420 1042.490 745.620 ;
        RECT 4.300 742.260 1042.490 743.420 ;
        RECT 4.000 740.060 1042.490 742.260 ;
        RECT 4.300 738.900 1042.490 740.060 ;
        RECT 4.000 736.700 1042.490 738.900 ;
        RECT 4.300 735.540 1042.490 736.700 ;
        RECT 4.000 733.340 1042.490 735.540 ;
        RECT 4.300 732.180 1042.490 733.340 ;
        RECT 4.000 729.980 1042.490 732.180 ;
        RECT 4.300 728.820 1042.490 729.980 ;
        RECT 4.000 726.620 1042.490 728.820 ;
        RECT 4.300 725.460 1042.490 726.620 ;
        RECT 4.000 723.260 1042.490 725.460 ;
        RECT 4.300 722.100 1042.490 723.260 ;
        RECT 4.000 719.900 1042.490 722.100 ;
        RECT 4.300 718.740 1042.490 719.900 ;
        RECT 4.000 716.540 1042.490 718.740 ;
        RECT 4.300 715.380 1042.490 716.540 ;
        RECT 4.000 713.180 1042.490 715.380 ;
        RECT 4.300 712.020 1042.490 713.180 ;
        RECT 4.000 709.820 1042.490 712.020 ;
        RECT 4.300 708.660 1042.490 709.820 ;
        RECT 4.000 706.460 1042.490 708.660 ;
        RECT 4.300 705.300 1042.490 706.460 ;
        RECT 4.000 703.100 1042.490 705.300 ;
        RECT 4.300 701.940 1042.490 703.100 ;
        RECT 4.000 699.740 1042.490 701.940 ;
        RECT 4.300 698.580 1042.490 699.740 ;
        RECT 4.000 696.380 1042.490 698.580 ;
        RECT 4.300 695.220 1042.490 696.380 ;
        RECT 4.000 693.020 1042.490 695.220 ;
        RECT 4.300 691.860 1042.490 693.020 ;
        RECT 4.000 689.660 1042.490 691.860 ;
        RECT 4.300 688.500 1042.490 689.660 ;
        RECT 4.000 686.300 1042.490 688.500 ;
        RECT 4.300 685.140 1042.490 686.300 ;
        RECT 4.000 682.940 1042.490 685.140 ;
        RECT 4.300 681.780 1042.490 682.940 ;
        RECT 4.000 679.580 1042.490 681.780 ;
        RECT 4.300 678.420 1042.490 679.580 ;
        RECT 4.000 676.220 1042.490 678.420 ;
        RECT 4.300 675.060 1042.490 676.220 ;
        RECT 4.000 672.860 1042.490 675.060 ;
        RECT 4.300 671.700 1042.490 672.860 ;
        RECT 4.000 669.500 1042.490 671.700 ;
        RECT 4.300 668.340 1042.490 669.500 ;
        RECT 4.000 666.140 1042.490 668.340 ;
        RECT 4.300 664.980 1042.490 666.140 ;
        RECT 4.000 662.780 1042.490 664.980 ;
        RECT 4.300 661.620 1042.490 662.780 ;
        RECT 4.000 659.420 1042.490 661.620 ;
        RECT 4.300 658.260 1042.490 659.420 ;
        RECT 4.000 656.060 1042.490 658.260 ;
        RECT 4.300 654.900 1042.490 656.060 ;
        RECT 4.000 652.700 1042.490 654.900 ;
        RECT 4.300 651.540 1042.490 652.700 ;
        RECT 4.000 649.340 1042.490 651.540 ;
        RECT 4.300 648.180 1042.490 649.340 ;
        RECT 4.000 645.980 1042.490 648.180 ;
        RECT 4.300 644.820 1042.490 645.980 ;
        RECT 4.000 642.620 1042.490 644.820 ;
        RECT 4.300 641.460 1042.490 642.620 ;
        RECT 4.000 639.260 1042.490 641.460 ;
        RECT 4.300 638.100 1042.490 639.260 ;
        RECT 4.000 635.900 1042.490 638.100 ;
        RECT 4.300 634.740 1042.490 635.900 ;
        RECT 4.000 632.540 1042.490 634.740 ;
        RECT 4.300 631.380 1042.490 632.540 ;
        RECT 4.000 629.180 1042.490 631.380 ;
        RECT 4.300 628.020 1042.490 629.180 ;
        RECT 4.000 625.820 1042.490 628.020 ;
        RECT 4.300 624.660 1042.490 625.820 ;
        RECT 4.000 622.460 1042.490 624.660 ;
        RECT 4.300 621.300 1042.490 622.460 ;
        RECT 4.000 619.100 1042.490 621.300 ;
        RECT 4.300 617.940 1042.490 619.100 ;
        RECT 4.000 615.740 1042.490 617.940 ;
        RECT 4.300 614.580 1042.490 615.740 ;
        RECT 4.000 612.380 1042.490 614.580 ;
        RECT 4.300 611.220 1042.490 612.380 ;
        RECT 4.000 609.020 1042.490 611.220 ;
        RECT 4.300 607.860 1042.490 609.020 ;
        RECT 4.000 605.660 1042.490 607.860 ;
        RECT 4.300 604.500 1042.490 605.660 ;
        RECT 4.000 602.300 1042.490 604.500 ;
        RECT 4.300 601.140 1042.490 602.300 ;
        RECT 4.000 598.940 1042.490 601.140 ;
        RECT 4.300 597.780 1042.490 598.940 ;
        RECT 4.000 595.580 1042.490 597.780 ;
        RECT 4.300 594.420 1042.490 595.580 ;
        RECT 4.000 592.220 1042.490 594.420 ;
        RECT 4.300 591.060 1042.490 592.220 ;
        RECT 4.000 588.860 1042.490 591.060 ;
        RECT 4.300 587.700 1042.490 588.860 ;
        RECT 4.000 585.500 1042.490 587.700 ;
        RECT 4.300 584.340 1042.490 585.500 ;
        RECT 4.000 582.140 1042.490 584.340 ;
        RECT 4.300 580.980 1042.490 582.140 ;
        RECT 4.000 578.780 1042.490 580.980 ;
        RECT 4.300 577.620 1042.490 578.780 ;
        RECT 4.000 575.420 1042.490 577.620 ;
        RECT 4.300 574.260 1042.490 575.420 ;
        RECT 4.000 572.060 1042.490 574.260 ;
        RECT 4.300 570.900 1042.490 572.060 ;
        RECT 4.000 568.700 1042.490 570.900 ;
        RECT 4.300 567.540 1042.490 568.700 ;
        RECT 4.000 565.340 1042.490 567.540 ;
        RECT 4.300 564.180 1042.490 565.340 ;
        RECT 4.000 561.980 1042.490 564.180 ;
        RECT 4.300 560.820 1042.490 561.980 ;
        RECT 4.000 558.620 1042.490 560.820 ;
        RECT 4.300 557.460 1042.490 558.620 ;
        RECT 4.000 555.260 1042.490 557.460 ;
        RECT 4.300 554.100 1042.490 555.260 ;
        RECT 4.000 551.900 1042.490 554.100 ;
        RECT 4.300 550.740 1042.490 551.900 ;
        RECT 4.000 548.540 1042.490 550.740 ;
        RECT 4.300 547.380 1042.490 548.540 ;
        RECT 4.000 545.180 1042.490 547.380 ;
        RECT 4.300 544.020 1042.490 545.180 ;
        RECT 4.000 541.820 1042.490 544.020 ;
        RECT 4.300 540.660 1042.490 541.820 ;
        RECT 4.000 538.460 1042.490 540.660 ;
        RECT 4.300 537.300 1042.490 538.460 ;
        RECT 4.000 535.100 1042.490 537.300 ;
        RECT 4.300 533.940 1042.490 535.100 ;
        RECT 4.000 531.740 1042.490 533.940 ;
        RECT 4.300 530.580 1042.490 531.740 ;
        RECT 4.000 528.380 1042.490 530.580 ;
        RECT 4.300 527.220 1042.490 528.380 ;
        RECT 4.000 31.100 1042.490 527.220 ;
        RECT 4.300 29.940 1042.490 31.100 ;
        RECT 4.000 27.740 1042.490 29.940 ;
        RECT 4.300 26.580 1042.490 27.740 ;
        RECT 4.000 24.380 1042.490 26.580 ;
        RECT 4.300 23.220 1042.490 24.380 ;
        RECT 4.000 21.020 1042.490 23.220 ;
        RECT 4.300 19.860 1042.490 21.020 ;
        RECT 4.000 17.660 1042.490 19.860 ;
        RECT 4.300 16.500 1042.490 17.660 ;
        RECT 4.000 14.300 1042.490 16.500 ;
        RECT 4.300 13.580 1042.490 14.300 ;
      LAYER Metal4 ;
        RECT 46.060 18.010 98.740 984.950 ;
        RECT 100.940 18.010 175.540 984.950 ;
        RECT 177.740 18.010 252.340 984.950 ;
        RECT 254.540 18.010 329.140 984.950 ;
        RECT 331.340 18.010 405.940 984.950 ;
        RECT 408.140 18.010 482.740 984.950 ;
        RECT 484.940 18.010 559.540 984.950 ;
        RECT 561.740 18.010 636.340 984.950 ;
        RECT 638.540 18.010 713.140 984.950 ;
        RECT 715.340 18.010 789.940 984.950 ;
        RECT 792.140 18.010 866.740 984.950 ;
        RECT 868.940 18.010 943.540 984.950 ;
        RECT 945.740 18.010 964.740 984.950 ;
  END
END top_ew_algofoogle
END LIBRARY

