magic
tech gf180mcuD
magscale 1 10
timestamp 1702302954
<< nwell >>
rect 1258 56071 26440 56096
rect 1258 55257 58662 56071
rect 1258 55232 2541 55257
rect 1258 54503 3110 54528
rect 1258 53689 58662 54503
rect 1258 53664 2541 53689
rect 1258 52935 20237 52960
rect 1258 52121 58662 52935
rect 1258 52096 2541 52121
rect 1258 51367 6237 51392
rect 1258 50553 58662 51367
rect 1258 50528 8925 50553
rect 1258 49799 2541 49824
rect 1258 48985 58662 49799
rect 1258 48960 15374 48985
rect 1258 48231 6616 48256
rect 1258 47417 58662 48231
rect 1258 47392 3592 47417
rect 1258 46663 18911 46688
rect 1258 45849 58662 46663
rect 1258 45824 3592 45849
rect 1258 45095 6685 45120
rect 1258 44281 58662 45095
rect 1258 44256 8925 44281
rect 1258 43527 3592 43552
rect 1258 42713 58662 43527
rect 1258 42688 8925 42713
rect 1258 41959 2541 41984
rect 1258 41145 58662 41959
rect 1258 41120 9037 41145
rect 1258 40391 7400 40416
rect 1258 39577 58662 40391
rect 1258 39552 2541 39577
rect 1258 38823 20190 38848
rect 1258 38009 58662 38823
rect 1258 37984 2541 38009
rect 1258 37255 10381 37280
rect 1258 36441 58662 37255
rect 1258 36416 25992 36441
rect 1258 35687 12733 35712
rect 1258 34873 58662 35687
rect 1258 34848 16541 34873
rect 1258 34119 21176 34144
rect 1258 33305 58662 34119
rect 1258 33280 14301 33305
rect 1258 32551 13069 32576
rect 1258 31737 58662 32551
rect 1258 31712 17475 31737
rect 1258 30983 10381 31008
rect 1258 30169 58662 30983
rect 1258 30144 14301 30169
rect 1258 29415 6013 29440
rect 1258 28601 58662 29415
rect 1258 28576 9933 28601
rect 1258 27847 4221 27872
rect 1258 27033 58662 27847
rect 1258 27008 16317 27033
rect 1258 26279 4893 26304
rect 1258 25465 58662 26279
rect 1258 25440 7021 25465
rect 1258 24711 23202 24736
rect 1258 23897 58662 24711
rect 1258 23872 2989 23897
rect 1258 23143 2653 23168
rect 1258 22329 58662 23143
rect 1258 22304 31997 22329
rect 1258 21575 3101 21600
rect 1258 20761 58662 21575
rect 1258 20736 2541 20761
rect 1258 20007 29197 20032
rect 1258 19193 58662 20007
rect 1258 19168 31997 19193
rect 1258 18439 3437 18464
rect 1258 17625 58662 18439
rect 1258 17600 2541 17625
rect 1258 16871 18221 16896
rect 1258 16057 58662 16871
rect 1258 16032 9261 16057
rect 1258 15303 3549 15328
rect 1258 14489 58662 15303
rect 1258 14464 2541 14489
rect 1258 13735 14904 13760
rect 1258 12921 58662 13735
rect 1258 12896 2541 12921
rect 1258 12167 3101 12192
rect 1258 11353 58662 12167
rect 1258 11328 16429 11353
rect 1258 10599 13293 10624
rect 1258 9785 58662 10599
rect 1258 9760 9149 9785
rect 1258 9031 6461 9056
rect 1258 8217 58662 9031
rect 1258 8192 16429 8217
rect 1258 7463 20237 7488
rect 1258 6649 58662 7463
rect 1258 6624 10157 6649
rect 1258 5895 12957 5920
rect 1258 5081 58662 5895
rect 1258 5056 16429 5081
rect 1258 4327 21245 4352
rect 1258 3488 58662 4327
<< pwell >>
rect 1258 56096 58662 56534
rect 1258 54528 58662 55232
rect 1258 52960 58662 53664
rect 1258 51392 58662 52096
rect 1258 49824 58662 50528
rect 1258 48256 58662 48960
rect 1258 46688 58662 47392
rect 1258 45120 58662 45824
rect 1258 43552 58662 44256
rect 1258 41984 58662 42688
rect 1258 40416 58662 41120
rect 1258 38848 58662 39552
rect 1258 37280 58662 37984
rect 1258 35712 58662 36416
rect 1258 34144 58662 34848
rect 1258 32576 58662 33280
rect 1258 31008 58662 31712
rect 1258 29440 58662 30144
rect 1258 27872 58662 28576
rect 1258 26304 58662 27008
rect 1258 24736 58662 25440
rect 1258 23168 58662 23872
rect 1258 21600 58662 22304
rect 1258 20032 58662 20736
rect 1258 18464 58662 19168
rect 1258 16896 58662 17600
rect 1258 15328 58662 16032
rect 1258 13760 58662 14464
rect 1258 12192 58662 12896
rect 1258 10624 58662 11328
rect 1258 9056 58662 9760
rect 1258 7488 58662 8192
rect 1258 5920 58662 6624
rect 1258 4352 58662 5056
rect 1258 3050 58662 3488
<< obsm1 >>
rect 1344 3076 58576 57090
<< metal2 >>
rect 4032 59200 4144 60000
rect 4480 59200 4592 60000
rect 4928 59200 5040 60000
rect 5376 59200 5488 60000
rect 5824 59200 5936 60000
rect 6272 59200 6384 60000
rect 6720 59200 6832 60000
rect 7168 59200 7280 60000
rect 7616 59200 7728 60000
rect 8064 59200 8176 60000
rect 8512 59200 8624 60000
rect 8960 59200 9072 60000
rect 9408 59200 9520 60000
rect 9856 59200 9968 60000
rect 10304 59200 10416 60000
rect 10752 59200 10864 60000
rect 11200 59200 11312 60000
rect 11648 59200 11760 60000
rect 12096 59200 12208 60000
rect 12544 59200 12656 60000
rect 12992 59200 13104 60000
rect 13440 59200 13552 60000
rect 13888 59200 14000 60000
rect 14336 59200 14448 60000
rect 14784 59200 14896 60000
rect 15232 59200 15344 60000
rect 15680 59200 15792 60000
rect 16128 59200 16240 60000
rect 16576 59200 16688 60000
rect 17024 59200 17136 60000
rect 17472 59200 17584 60000
rect 17920 59200 18032 60000
rect 18368 59200 18480 60000
rect 18816 59200 18928 60000
rect 19264 59200 19376 60000
rect 19712 59200 19824 60000
rect 20160 59200 20272 60000
rect 20608 59200 20720 60000
rect 21056 59200 21168 60000
rect 21504 59200 21616 60000
rect 21952 59200 22064 60000
rect 22400 59200 22512 60000
rect 22848 59200 22960 60000
rect 23296 59200 23408 60000
rect 23744 59200 23856 60000
rect 24192 59200 24304 60000
rect 24640 59200 24752 60000
rect 25088 59200 25200 60000
rect 25536 59200 25648 60000
rect 25984 59200 26096 60000
rect 26432 59200 26544 60000
rect 26880 59200 26992 60000
rect 27328 59200 27440 60000
rect 27776 59200 27888 60000
rect 28224 59200 28336 60000
rect 28672 59200 28784 60000
rect 29120 59200 29232 60000
rect 29568 59200 29680 60000
rect 30016 59200 30128 60000
rect 30464 59200 30576 60000
rect 30912 59200 31024 60000
rect 31360 59200 31472 60000
rect 31808 59200 31920 60000
rect 32256 59200 32368 60000
rect 32704 59200 32816 60000
rect 33152 59200 33264 60000
rect 33600 59200 33712 60000
rect 34048 59200 34160 60000
rect 34496 59200 34608 60000
rect 34944 59200 35056 60000
rect 35392 59200 35504 60000
rect 35840 59200 35952 60000
rect 36288 59200 36400 60000
rect 36736 59200 36848 60000
rect 37184 59200 37296 60000
rect 37632 59200 37744 60000
rect 38080 59200 38192 60000
rect 38528 59200 38640 60000
rect 38976 59200 39088 60000
rect 39424 59200 39536 60000
rect 39872 59200 39984 60000
rect 40320 59200 40432 60000
rect 40768 59200 40880 60000
rect 41216 59200 41328 60000
rect 41664 59200 41776 60000
rect 42112 59200 42224 60000
rect 42560 59200 42672 60000
rect 43008 59200 43120 60000
rect 43456 59200 43568 60000
rect 43904 59200 44016 60000
rect 44352 59200 44464 60000
rect 44800 59200 44912 60000
rect 45248 59200 45360 60000
rect 45696 59200 45808 60000
rect 46144 59200 46256 60000
rect 46592 59200 46704 60000
rect 47040 59200 47152 60000
rect 47488 59200 47600 60000
rect 47936 59200 48048 60000
rect 48384 59200 48496 60000
rect 48832 59200 48944 60000
rect 49280 59200 49392 60000
rect 49728 59200 49840 60000
rect 50176 59200 50288 60000
rect 50624 59200 50736 60000
rect 51072 59200 51184 60000
rect 51520 59200 51632 60000
rect 51968 59200 52080 60000
rect 52416 59200 52528 60000
rect 52864 59200 52976 60000
rect 53312 59200 53424 60000
rect 53760 59200 53872 60000
rect 54208 59200 54320 60000
rect 54656 59200 54768 60000
rect 55104 59200 55216 60000
rect 55552 59200 55664 60000
<< obsm2 >>
rect 1596 59140 3972 59200
rect 4204 59140 4420 59200
rect 4652 59140 4868 59200
rect 5100 59140 5316 59200
rect 5548 59140 5764 59200
rect 5996 59140 6212 59200
rect 6444 59140 6660 59200
rect 6892 59140 7108 59200
rect 7340 59140 7556 59200
rect 7788 59140 8004 59200
rect 8236 59140 8452 59200
rect 8684 59140 8900 59200
rect 9132 59140 9348 59200
rect 9580 59140 9796 59200
rect 10028 59140 10244 59200
rect 10476 59140 10692 59200
rect 10924 59140 11140 59200
rect 11372 59140 11588 59200
rect 11820 59140 12036 59200
rect 12268 59140 12484 59200
rect 12716 59140 12932 59200
rect 13164 59140 13380 59200
rect 13612 59140 13828 59200
rect 14060 59140 14276 59200
rect 14508 59140 14724 59200
rect 14956 59140 15172 59200
rect 15404 59140 15620 59200
rect 15852 59140 16068 59200
rect 16300 59140 16516 59200
rect 16748 59140 16964 59200
rect 17196 59140 17412 59200
rect 17644 59140 17860 59200
rect 18092 59140 18308 59200
rect 18540 59140 18756 59200
rect 18988 59140 19204 59200
rect 19436 59140 19652 59200
rect 19884 59140 20100 59200
rect 20332 59140 20548 59200
rect 20780 59140 20996 59200
rect 21228 59140 21444 59200
rect 21676 59140 21892 59200
rect 22124 59140 22340 59200
rect 22572 59140 22788 59200
rect 23020 59140 23236 59200
rect 23468 59140 23684 59200
rect 23916 59140 24132 59200
rect 24364 59140 24580 59200
rect 24812 59140 25028 59200
rect 25260 59140 25476 59200
rect 25708 59140 25924 59200
rect 26156 59140 26372 59200
rect 26604 59140 26820 59200
rect 27052 59140 27268 59200
rect 27500 59140 27716 59200
rect 27948 59140 28164 59200
rect 28396 59140 28612 59200
rect 28844 59140 29060 59200
rect 29292 59140 29508 59200
rect 29740 59140 29956 59200
rect 30188 59140 30404 59200
rect 30636 59140 30852 59200
rect 31084 59140 31300 59200
rect 31532 59140 31748 59200
rect 31980 59140 32196 59200
rect 32428 59140 32644 59200
rect 32876 59140 33092 59200
rect 33324 59140 33540 59200
rect 33772 59140 33988 59200
rect 34220 59140 34436 59200
rect 34668 59140 34884 59200
rect 35116 59140 35332 59200
rect 35564 59140 35780 59200
rect 36012 59140 36228 59200
rect 36460 59140 36676 59200
rect 36908 59140 37124 59200
rect 37356 59140 37572 59200
rect 37804 59140 38020 59200
rect 38252 59140 38468 59200
rect 38700 59140 38916 59200
rect 39148 59140 39364 59200
rect 39596 59140 39812 59200
rect 40044 59140 40260 59200
rect 40492 59140 40708 59200
rect 40940 59140 41156 59200
rect 41388 59140 41604 59200
rect 41836 59140 42052 59200
rect 42284 59140 42500 59200
rect 42732 59140 42948 59200
rect 43180 59140 43396 59200
rect 43628 59140 43844 59200
rect 44076 59140 44292 59200
rect 44524 59140 44740 59200
rect 44972 59140 45188 59200
rect 45420 59140 45636 59200
rect 45868 59140 46084 59200
rect 46316 59140 46532 59200
rect 46764 59140 46980 59200
rect 47212 59140 47428 59200
rect 47660 59140 47876 59200
rect 48108 59140 48324 59200
rect 48556 59140 48772 59200
rect 49004 59140 49220 59200
rect 49452 59140 49668 59200
rect 49900 59140 50116 59200
rect 50348 59140 50564 59200
rect 50796 59140 51012 59200
rect 51244 59140 51460 59200
rect 51692 59140 51908 59200
rect 52140 59140 52356 59200
rect 52588 59140 52804 59200
rect 53036 59140 53252 59200
rect 53484 59140 53700 59200
rect 53932 59140 54148 59200
rect 54380 59140 54596 59200
rect 54828 59140 55044 59200
rect 55276 59140 55492 59200
rect 55724 59140 58212 59200
rect 1596 3098 58212 59140
<< obsm3 >>
rect 1586 3108 58222 57092
<< metal4 >>
rect 4448 3076 4768 56508
rect 19808 3076 20128 56508
rect 35168 3076 35488 56508
rect 50528 3076 50848 56508
<< obsm4 >>
rect 4284 7634 4388 50718
rect 4828 7634 19748 50718
rect 20188 7634 35108 50718
rect 35548 7634 48692 50718
<< labels >>
rlabel metal2 s 4928 59200 5040 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 18368 59200 18480 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 19712 59200 19824 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 21056 59200 21168 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 22400 59200 22512 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 23744 59200 23856 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 25088 59200 25200 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 26432 59200 26544 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 27776 59200 27888 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 29120 59200 29232 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 30464 59200 30576 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6272 59200 6384 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 31808 59200 31920 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 33152 59200 33264 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 34496 59200 34608 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 35840 59200 35952 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 37184 59200 37296 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 38528 59200 38640 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 39872 59200 39984 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 41216 59200 41328 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 42560 59200 42672 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 43904 59200 44016 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 7616 59200 7728 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 45248 59200 45360 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 46592 59200 46704 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 47936 59200 48048 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 49280 59200 49392 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 50624 59200 50736 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 51968 59200 52080 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 53312 59200 53424 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 54656 59200 54768 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8960 59200 9072 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10304 59200 10416 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 11648 59200 11760 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 12992 59200 13104 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 14336 59200 14448 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 15680 59200 15792 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 17024 59200 17136 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5376 59200 5488 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 18816 59200 18928 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 20160 59200 20272 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 21504 59200 21616 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 22848 59200 22960 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 24192 59200 24304 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 25536 59200 25648 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 26880 59200 26992 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 28224 59200 28336 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 29568 59200 29680 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 30912 59200 31024 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6720 59200 6832 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 32256 59200 32368 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 33600 59200 33712 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 34944 59200 35056 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 36288 59200 36400 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 37632 59200 37744 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 38976 59200 39088 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 40320 59200 40432 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 41664 59200 41776 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 43008 59200 43120 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 44352 59200 44464 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 8064 59200 8176 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 45696 59200 45808 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 47040 59200 47152 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 48384 59200 48496 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 49728 59200 49840 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 51072 59200 51184 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 52416 59200 52528 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 53760 59200 53872 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 55104 59200 55216 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9408 59200 9520 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 10752 59200 10864 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 12096 59200 12208 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 13440 59200 13552 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 14784 59200 14896 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 16128 59200 16240 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 17472 59200 17584 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5824 59200 5936 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 19264 59200 19376 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 20608 59200 20720 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 21952 59200 22064 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 23296 59200 23408 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 24640 59200 24752 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 25984 59200 26096 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 27328 59200 27440 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 28672 59200 28784 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 30016 59200 30128 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 31360 59200 31472 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7168 59200 7280 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 32704 59200 32816 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 34048 59200 34160 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 35392 59200 35504 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 36736 59200 36848 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 38080 59200 38192 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 39424 59200 39536 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 40768 59200 40880 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 42112 59200 42224 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 43456 59200 43568 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 44800 59200 44912 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8512 59200 8624 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 46144 59200 46256 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 47488 59200 47600 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 48832 59200 48944 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 50176 59200 50288 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 51520 59200 51632 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 52864 59200 52976 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 54208 59200 54320 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 55552 59200 55664 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9856 59200 9968 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 11200 59200 11312 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 12544 59200 12656 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 13888 59200 14000 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 15232 59200 15344 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 16576 59200 16688 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 17920 59200 18032 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 4448 3076 4768 56508 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 56508 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 56508 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 56508 6 vss
port 116 nsew ground bidirectional
rlabel metal2 s 4032 59200 4144 60000 6 wb_clk_i
port 117 nsew signal input
rlabel metal2 s 4480 59200 4592 60000 6 wb_rst_i
port 118 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2752652
string GDS_FILE /home/zerotoasic/anton/algofoogle-multi-caravel/openlane/urish_simon_says/runs/23_12_12_00_24/results/signoff/urish_simon_says.magic.gds
string GDS_START 371498
<< end >>

