VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO urish_simon_says
  CLASS BLOCK ;
  FOREIGN urish_simon_says ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 296.000 25.200 300.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 296.000 92.400 300.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 296.000 99.120 300.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 296.000 105.840 300.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 296.000 112.560 300.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 296.000 119.280 300.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 296.000 126.000 300.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 296.000 132.720 300.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 296.000 139.440 300.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 296.000 146.160 300.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 296.000 152.880 300.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 296.000 31.920 300.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 296.000 159.600 300.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 296.000 166.320 300.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 296.000 173.040 300.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 296.000 179.760 300.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 296.000 186.480 300.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 296.000 193.200 300.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 296.000 199.920 300.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 296.000 206.640 300.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 296.000 213.360 300.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 296.000 220.080 300.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 296.000 38.640 300.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 296.000 226.800 300.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.960 296.000 233.520 300.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 296.000 240.240 300.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 296.000 246.960 300.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 296.000 253.680 300.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 296.000 260.400 300.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 296.000 267.120 300.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 296.000 273.840 300.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 296.000 45.360 300.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 296.000 52.080 300.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 296.000 58.800 300.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 296.000 65.520 300.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 296.000 72.240 300.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 296.000 78.960 300.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 296.000 85.680 300.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 296.000 27.440 300.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 296.000 94.640 300.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 296.000 101.360 300.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 296.000 108.080 300.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 296.000 114.800 300.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 296.000 121.520 300.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 296.000 128.240 300.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 296.000 134.960 300.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 296.000 141.680 300.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 296.000 148.400 300.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 296.000 155.120 300.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 296.000 34.160 300.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 296.000 161.840 300.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 296.000 168.560 300.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 296.000 175.280 300.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 296.000 182.000 300.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 296.000 188.720 300.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 296.000 195.440 300.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 296.000 202.160 300.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 296.000 208.880 300.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 296.000 215.600 300.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 296.000 222.320 300.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 296.000 40.880 300.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 296.000 229.040 300.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 296.000 235.760 300.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 296.000 242.480 300.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 296.000 249.200 300.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 296.000 255.920 300.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 296.000 262.640 300.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 296.000 269.360 300.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 296.000 276.080 300.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 296.000 47.600 300.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 296.000 54.320 300.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 296.000 61.040 300.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 296.000 67.760 300.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 296.000 74.480 300.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 296.000 81.200 300.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 296.000 87.920 300.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 296.000 29.680 300.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 296.000 96.880 300.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 296.000 103.600 300.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 296.000 110.320 300.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 296.000 117.040 300.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 296.000 123.760 300.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 296.000 130.480 300.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 296.000 137.200 300.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 296.000 143.920 300.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 296.000 150.640 300.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 296.000 157.360 300.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 296.000 36.400 300.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 296.000 164.080 300.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 296.000 170.800 300.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 296.000 177.520 300.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 296.000 184.240 300.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 296.000 190.960 300.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 296.000 197.680 300.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 296.000 204.400 300.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 296.000 211.120 300.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 296.000 217.840 300.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 296.000 224.560 300.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 296.000 43.120 300.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 296.000 231.280 300.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 296.000 238.000 300.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 296.000 244.720 300.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 250.880 296.000 251.440 300.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 296.000 258.160 300.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 264.320 296.000 264.880 300.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 296.000 271.600 300.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 296.000 278.320 300.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 296.000 49.840 300.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 296.000 56.560 300.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 296.000 63.280 300.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 296.000 70.000 300.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 296.000 76.720 300.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 296.000 83.440 300.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 296.000 90.160 300.000 ;
    END
  END io_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 296.000 20.720 300.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 296.000 22.960 300.000 ;
    END
  END wb_rst_i
  OBS
      LAYER Pwell ;
        RECT 6.290 280.480 293.310 282.670 ;
      LAYER Nwell ;
        RECT 6.290 280.355 132.200 280.480 ;
        RECT 6.290 276.285 293.310 280.355 ;
        RECT 6.290 276.160 12.705 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 293.310 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 15.550 272.640 ;
        RECT 6.290 268.445 293.310 272.515 ;
        RECT 6.290 268.320 12.705 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 293.310 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 101.185 264.800 ;
        RECT 6.290 260.605 293.310 264.675 ;
        RECT 6.290 260.480 12.705 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 293.310 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 31.185 256.960 ;
        RECT 6.290 252.765 293.310 256.835 ;
        RECT 6.290 252.640 44.625 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 293.310 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 12.705 249.120 ;
        RECT 6.290 244.925 293.310 248.995 ;
        RECT 6.290 244.800 76.870 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 293.310 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 33.080 241.280 ;
        RECT 6.290 237.085 293.310 241.155 ;
        RECT 6.290 236.960 17.960 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 293.310 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 94.555 233.440 ;
        RECT 6.290 229.245 293.310 233.315 ;
        RECT 6.290 229.120 17.960 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 293.310 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 33.425 225.600 ;
        RECT 6.290 221.405 293.310 225.475 ;
        RECT 6.290 221.280 44.625 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 293.310 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 17.960 217.760 ;
        RECT 6.290 213.565 293.310 217.635 ;
        RECT 6.290 213.440 44.625 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 293.310 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 12.705 209.920 ;
        RECT 6.290 205.725 293.310 209.795 ;
        RECT 6.290 205.600 45.185 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 293.310 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 37.000 202.080 ;
        RECT 6.290 197.885 293.310 201.955 ;
        RECT 6.290 197.760 12.705 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 293.310 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 100.950 194.240 ;
        RECT 6.290 190.045 293.310 194.115 ;
        RECT 6.290 189.920 12.705 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 293.310 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 51.905 186.400 ;
        RECT 6.290 182.205 293.310 186.275 ;
        RECT 6.290 182.080 129.960 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 293.310 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 63.665 178.560 ;
        RECT 6.290 174.365 293.310 178.435 ;
        RECT 6.290 174.240 82.705 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 293.310 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 105.880 170.720 ;
        RECT 6.290 166.525 293.310 170.595 ;
        RECT 6.290 166.400 71.505 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 293.310 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 65.345 162.880 ;
        RECT 6.290 158.685 293.310 162.755 ;
        RECT 6.290 158.560 87.375 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 293.310 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 51.905 155.040 ;
        RECT 6.290 150.845 293.310 154.915 ;
        RECT 6.290 150.720 71.505 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 293.310 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 30.065 147.200 ;
        RECT 6.290 143.005 293.310 147.075 ;
        RECT 6.290 142.880 49.665 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 293.310 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 21.105 139.360 ;
        RECT 6.290 135.165 293.310 139.235 ;
        RECT 6.290 135.040 81.585 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 293.310 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 24.465 131.520 ;
        RECT 6.290 127.325 293.310 131.395 ;
        RECT 6.290 127.200 35.105 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 293.310 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 116.010 123.680 ;
        RECT 6.290 119.485 293.310 123.555 ;
        RECT 6.290 119.360 14.945 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 293.310 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 13.265 115.840 ;
        RECT 6.290 111.645 293.310 115.715 ;
        RECT 6.290 111.520 159.985 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 293.310 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 15.505 108.000 ;
        RECT 6.290 103.805 293.310 107.875 ;
        RECT 6.290 103.680 12.705 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 293.310 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 145.985 100.160 ;
        RECT 6.290 95.965 293.310 100.035 ;
        RECT 6.290 95.840 159.985 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 293.310 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 17.185 92.320 ;
        RECT 6.290 88.125 293.310 92.195 ;
        RECT 6.290 88.000 12.705 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 293.310 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 91.105 84.480 ;
        RECT 6.290 80.285 293.310 84.355 ;
        RECT 6.290 80.160 46.305 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 293.310 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 17.745 76.640 ;
        RECT 6.290 72.445 293.310 76.515 ;
        RECT 6.290 72.320 12.705 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 293.310 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 74.520 68.800 ;
        RECT 6.290 64.605 293.310 68.675 ;
        RECT 6.290 64.480 12.705 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 293.310 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 15.505 60.960 ;
        RECT 6.290 56.765 293.310 60.835 ;
        RECT 6.290 56.640 82.145 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 293.310 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 66.465 53.120 ;
        RECT 6.290 48.925 293.310 52.995 ;
        RECT 6.290 48.800 45.745 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 293.310 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 32.305 45.280 ;
        RECT 6.290 41.085 293.310 45.155 ;
        RECT 6.290 40.960 82.145 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 293.310 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 101.185 37.440 ;
        RECT 6.290 33.245 293.310 37.315 ;
        RECT 6.290 33.120 50.785 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 293.310 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 64.785 29.600 ;
        RECT 6.290 25.405 293.310 29.475 ;
        RECT 6.290 25.280 82.145 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 293.310 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 106.225 21.760 ;
        RECT 6.290 17.440 293.310 21.635 ;
      LAYER Pwell ;
        RECT 6.290 15.250 293.310 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 285.450 ;
      LAYER Metal2 ;
        RECT 7.980 295.700 19.860 296.000 ;
        RECT 21.020 295.700 22.100 296.000 ;
        RECT 23.260 295.700 24.340 296.000 ;
        RECT 25.500 295.700 26.580 296.000 ;
        RECT 27.740 295.700 28.820 296.000 ;
        RECT 29.980 295.700 31.060 296.000 ;
        RECT 32.220 295.700 33.300 296.000 ;
        RECT 34.460 295.700 35.540 296.000 ;
        RECT 36.700 295.700 37.780 296.000 ;
        RECT 38.940 295.700 40.020 296.000 ;
        RECT 41.180 295.700 42.260 296.000 ;
        RECT 43.420 295.700 44.500 296.000 ;
        RECT 45.660 295.700 46.740 296.000 ;
        RECT 47.900 295.700 48.980 296.000 ;
        RECT 50.140 295.700 51.220 296.000 ;
        RECT 52.380 295.700 53.460 296.000 ;
        RECT 54.620 295.700 55.700 296.000 ;
        RECT 56.860 295.700 57.940 296.000 ;
        RECT 59.100 295.700 60.180 296.000 ;
        RECT 61.340 295.700 62.420 296.000 ;
        RECT 63.580 295.700 64.660 296.000 ;
        RECT 65.820 295.700 66.900 296.000 ;
        RECT 68.060 295.700 69.140 296.000 ;
        RECT 70.300 295.700 71.380 296.000 ;
        RECT 72.540 295.700 73.620 296.000 ;
        RECT 74.780 295.700 75.860 296.000 ;
        RECT 77.020 295.700 78.100 296.000 ;
        RECT 79.260 295.700 80.340 296.000 ;
        RECT 81.500 295.700 82.580 296.000 ;
        RECT 83.740 295.700 84.820 296.000 ;
        RECT 85.980 295.700 87.060 296.000 ;
        RECT 88.220 295.700 89.300 296.000 ;
        RECT 90.460 295.700 91.540 296.000 ;
        RECT 92.700 295.700 93.780 296.000 ;
        RECT 94.940 295.700 96.020 296.000 ;
        RECT 97.180 295.700 98.260 296.000 ;
        RECT 99.420 295.700 100.500 296.000 ;
        RECT 101.660 295.700 102.740 296.000 ;
        RECT 103.900 295.700 104.980 296.000 ;
        RECT 106.140 295.700 107.220 296.000 ;
        RECT 108.380 295.700 109.460 296.000 ;
        RECT 110.620 295.700 111.700 296.000 ;
        RECT 112.860 295.700 113.940 296.000 ;
        RECT 115.100 295.700 116.180 296.000 ;
        RECT 117.340 295.700 118.420 296.000 ;
        RECT 119.580 295.700 120.660 296.000 ;
        RECT 121.820 295.700 122.900 296.000 ;
        RECT 124.060 295.700 125.140 296.000 ;
        RECT 126.300 295.700 127.380 296.000 ;
        RECT 128.540 295.700 129.620 296.000 ;
        RECT 130.780 295.700 131.860 296.000 ;
        RECT 133.020 295.700 134.100 296.000 ;
        RECT 135.260 295.700 136.340 296.000 ;
        RECT 137.500 295.700 138.580 296.000 ;
        RECT 139.740 295.700 140.820 296.000 ;
        RECT 141.980 295.700 143.060 296.000 ;
        RECT 144.220 295.700 145.300 296.000 ;
        RECT 146.460 295.700 147.540 296.000 ;
        RECT 148.700 295.700 149.780 296.000 ;
        RECT 150.940 295.700 152.020 296.000 ;
        RECT 153.180 295.700 154.260 296.000 ;
        RECT 155.420 295.700 156.500 296.000 ;
        RECT 157.660 295.700 158.740 296.000 ;
        RECT 159.900 295.700 160.980 296.000 ;
        RECT 162.140 295.700 163.220 296.000 ;
        RECT 164.380 295.700 165.460 296.000 ;
        RECT 166.620 295.700 167.700 296.000 ;
        RECT 168.860 295.700 169.940 296.000 ;
        RECT 171.100 295.700 172.180 296.000 ;
        RECT 173.340 295.700 174.420 296.000 ;
        RECT 175.580 295.700 176.660 296.000 ;
        RECT 177.820 295.700 178.900 296.000 ;
        RECT 180.060 295.700 181.140 296.000 ;
        RECT 182.300 295.700 183.380 296.000 ;
        RECT 184.540 295.700 185.620 296.000 ;
        RECT 186.780 295.700 187.860 296.000 ;
        RECT 189.020 295.700 190.100 296.000 ;
        RECT 191.260 295.700 192.340 296.000 ;
        RECT 193.500 295.700 194.580 296.000 ;
        RECT 195.740 295.700 196.820 296.000 ;
        RECT 197.980 295.700 199.060 296.000 ;
        RECT 200.220 295.700 201.300 296.000 ;
        RECT 202.460 295.700 203.540 296.000 ;
        RECT 204.700 295.700 205.780 296.000 ;
        RECT 206.940 295.700 208.020 296.000 ;
        RECT 209.180 295.700 210.260 296.000 ;
        RECT 211.420 295.700 212.500 296.000 ;
        RECT 213.660 295.700 214.740 296.000 ;
        RECT 215.900 295.700 216.980 296.000 ;
        RECT 218.140 295.700 219.220 296.000 ;
        RECT 220.380 295.700 221.460 296.000 ;
        RECT 222.620 295.700 223.700 296.000 ;
        RECT 224.860 295.700 225.940 296.000 ;
        RECT 227.100 295.700 228.180 296.000 ;
        RECT 229.340 295.700 230.420 296.000 ;
        RECT 231.580 295.700 232.660 296.000 ;
        RECT 233.820 295.700 234.900 296.000 ;
        RECT 236.060 295.700 237.140 296.000 ;
        RECT 238.300 295.700 239.380 296.000 ;
        RECT 240.540 295.700 241.620 296.000 ;
        RECT 242.780 295.700 243.860 296.000 ;
        RECT 245.020 295.700 246.100 296.000 ;
        RECT 247.260 295.700 248.340 296.000 ;
        RECT 249.500 295.700 250.580 296.000 ;
        RECT 251.740 295.700 252.820 296.000 ;
        RECT 253.980 295.700 255.060 296.000 ;
        RECT 256.220 295.700 257.300 296.000 ;
        RECT 258.460 295.700 259.540 296.000 ;
        RECT 260.700 295.700 261.780 296.000 ;
        RECT 262.940 295.700 264.020 296.000 ;
        RECT 265.180 295.700 266.260 296.000 ;
        RECT 267.420 295.700 268.500 296.000 ;
        RECT 269.660 295.700 270.740 296.000 ;
        RECT 271.900 295.700 272.980 296.000 ;
        RECT 274.140 295.700 275.220 296.000 ;
        RECT 276.380 295.700 277.460 296.000 ;
        RECT 278.620 295.700 291.060 296.000 ;
        RECT 7.980 15.490 291.060 295.700 ;
      LAYER Metal3 ;
        RECT 7.930 15.540 291.110 285.460 ;
      LAYER Metal4 ;
        RECT 21.420 38.170 21.940 253.590 ;
        RECT 24.140 38.170 98.740 253.590 ;
        RECT 100.940 38.170 175.540 253.590 ;
        RECT 177.740 38.170 243.460 253.590 ;
  END
END urish_simon_says
END LIBRARY

