magic
tech gf180mcuD
magscale 1 10
timestamp 1701411205
<< obsm1 >>
rect 1344 3076 192528 193708
<< metal2 >>
rect 2688 196755 2800 197555
rect 18144 196755 18256 197555
rect 22176 196755 22288 197555
rect 36288 196755 36400 197555
rect 121632 196755 121744 197555
rect 126336 196755 126448 197555
rect 133728 196755 133840 197555
rect 134400 196755 134512 197555
rect 137760 196755 137872 197555
rect 141120 196755 141232 197555
rect 142464 196755 142576 197555
rect 148512 196755 148624 197555
rect 153888 196755 154000 197555
rect 154560 196755 154672 197555
rect 155232 196755 155344 197555
rect 157920 196755 158032 197555
rect 166656 196755 166768 197555
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 26208 0 26320 800
rect 50400 0 50512 800
rect 51072 0 51184 800
rect 52416 0 52528 800
rect 55776 0 55888 800
rect 83328 0 83440 800
rect 92736 0 92848 800
rect 110880 0 110992 800
rect 112224 0 112336 800
rect 114912 0 115024 800
rect 134400 0 134512 800
rect 159264 0 159376 800
rect 161280 0 161392 800
rect 168672 0 168784 800
rect 170016 0 170128 800
rect 181440 0 181552 800
rect 183456 0 183568 800
rect 185472 0 185584 800
rect 186144 0 186256 800
rect 188832 0 188944 800
rect 190848 0 190960 800
<< obsm2 >>
rect 1596 196695 2628 196868
rect 2860 196695 18084 196868
rect 18316 196695 22116 196868
rect 22348 196695 36228 196868
rect 36460 196695 121572 196868
rect 121804 196695 126276 196868
rect 126508 196695 133668 196868
rect 133900 196695 134340 196868
rect 134572 196695 137700 196868
rect 137932 196695 141060 196868
rect 141292 196695 142404 196868
rect 142636 196695 148452 196868
rect 148684 196695 153828 196868
rect 154060 196695 154500 196868
rect 154732 196695 155172 196868
rect 155404 196695 157860 196868
rect 158092 196695 166596 196868
rect 166828 196695 192164 196868
rect 1596 860 192164 196695
rect 1596 800 26148 860
rect 26380 800 50340 860
rect 50572 800 51012 860
rect 51244 800 52356 860
rect 52588 800 55716 860
rect 55948 800 83268 860
rect 83500 800 92676 860
rect 92908 800 110820 860
rect 111052 800 112164 860
rect 112396 800 114852 860
rect 115084 800 134340 860
rect 134572 800 159204 860
rect 159436 800 161220 860
rect 161452 800 168612 860
rect 168844 800 169956 860
rect 170188 800 181380 860
rect 181612 800 183396 860
rect 183628 800 185412 860
rect 185644 800 186084 860
rect 186316 800 188772 860
rect 189004 800 190788 860
rect 191020 800 192164 860
<< metal3 >>
rect 193171 193536 193971 193648
rect 193171 192864 193971 192976
rect 193171 192192 193971 192304
rect 193171 191520 193971 191632
rect 193171 190848 193971 190960
rect 193171 188832 193971 188944
rect 0 184128 800 184240
rect 193171 171360 193971 171472
rect 0 144480 800 144592
rect 0 143808 800 143920
rect 0 143136 800 143248
rect 0 142464 800 142576
rect 0 141792 800 141904
rect 0 141120 800 141232
rect 0 140448 800 140560
rect 0 139776 800 139888
rect 0 139104 800 139216
rect 0 138432 800 138544
rect 0 137760 800 137872
rect 0 137088 800 137200
rect 0 136416 800 136528
rect 0 135744 800 135856
rect 0 135072 800 135184
rect 0 134400 800 134512
rect 0 133728 800 133840
rect 0 133056 800 133168
rect 0 132384 800 132496
rect 0 131712 800 131824
rect 0 131040 800 131152
rect 0 130368 800 130480
rect 0 129696 800 129808
rect 0 129024 800 129136
rect 0 128352 800 128464
rect 0 127680 800 127792
rect 0 127008 800 127120
rect 0 126336 800 126448
rect 0 125664 800 125776
rect 0 124992 800 125104
rect 0 124320 800 124432
rect 0 123648 800 123760
rect 0 122976 800 123088
rect 0 122304 800 122416
rect 0 121632 800 121744
rect 0 120960 800 121072
rect 0 120288 800 120400
rect 0 119616 800 119728
rect 0 118944 800 119056
rect 0 118272 800 118384
rect 0 117600 800 117712
rect 0 116928 800 117040
rect 0 116256 800 116368
rect 0 115584 800 115696
rect 0 114912 800 115024
rect 0 114240 800 114352
rect 0 113568 800 113680
rect 0 112896 800 113008
rect 0 112224 800 112336
rect 0 111552 800 111664
rect 0 110880 800 110992
rect 0 110208 800 110320
rect 0 109536 800 109648
rect 0 108864 800 108976
rect 0 108192 800 108304
rect 0 107520 800 107632
rect 0 106848 800 106960
rect 0 106176 800 106288
rect 0 105504 800 105616
rect 0 104832 800 104944
rect 0 104160 800 104272
rect 0 103488 800 103600
rect 0 102816 800 102928
rect 0 102144 800 102256
rect 0 101472 800 101584
rect 0 100800 800 100912
rect 0 100128 800 100240
rect 0 99456 800 99568
rect 0 98784 800 98896
rect 0 98112 800 98224
rect 0 97440 800 97552
rect 0 96768 800 96880
rect 0 96096 800 96208
rect 0 10752 800 10864
rect 0 9408 800 9520
rect 0 8736 800 8848
rect 0 6720 800 6832
rect 0 6048 800 6160
rect 0 5376 800 5488
rect 0 4704 800 4816
rect 0 4032 800 4144
<< obsm3 >>
rect 800 193476 193111 193676
rect 800 193036 193171 193476
rect 800 192804 193111 193036
rect 800 192364 193171 192804
rect 800 192132 193111 192364
rect 800 191692 193171 192132
rect 800 191460 193111 191692
rect 800 191020 193171 191460
rect 800 190788 193111 191020
rect 800 189004 193171 190788
rect 800 188772 193111 189004
rect 800 184300 193171 188772
rect 860 184068 193171 184300
rect 800 171532 193171 184068
rect 800 171300 193111 171532
rect 800 144652 193171 171300
rect 860 144420 193171 144652
rect 800 143980 193171 144420
rect 860 143748 193171 143980
rect 800 143308 193171 143748
rect 860 143076 193171 143308
rect 800 142636 193171 143076
rect 860 142404 193171 142636
rect 800 141964 193171 142404
rect 860 141732 193171 141964
rect 800 141292 193171 141732
rect 860 141060 193171 141292
rect 800 140620 193171 141060
rect 860 140388 193171 140620
rect 800 139948 193171 140388
rect 860 139716 193171 139948
rect 800 139276 193171 139716
rect 860 139044 193171 139276
rect 800 138604 193171 139044
rect 860 138372 193171 138604
rect 800 137932 193171 138372
rect 860 137700 193171 137932
rect 800 137260 193171 137700
rect 860 137028 193171 137260
rect 800 136588 193171 137028
rect 860 136356 193171 136588
rect 800 135916 193171 136356
rect 860 135684 193171 135916
rect 800 135244 193171 135684
rect 860 135012 193171 135244
rect 800 134572 193171 135012
rect 860 134340 193171 134572
rect 800 133900 193171 134340
rect 860 133668 193171 133900
rect 800 133228 193171 133668
rect 860 132996 193171 133228
rect 800 132556 193171 132996
rect 860 132324 193171 132556
rect 800 131884 193171 132324
rect 860 131652 193171 131884
rect 800 131212 193171 131652
rect 860 130980 193171 131212
rect 800 130540 193171 130980
rect 860 130308 193171 130540
rect 800 129868 193171 130308
rect 860 129636 193171 129868
rect 800 129196 193171 129636
rect 860 128964 193171 129196
rect 800 128524 193171 128964
rect 860 128292 193171 128524
rect 800 127852 193171 128292
rect 860 127620 193171 127852
rect 800 127180 193171 127620
rect 860 126948 193171 127180
rect 800 126508 193171 126948
rect 860 126276 193171 126508
rect 800 125836 193171 126276
rect 860 125604 193171 125836
rect 800 125164 193171 125604
rect 860 124932 193171 125164
rect 800 124492 193171 124932
rect 860 124260 193171 124492
rect 800 123820 193171 124260
rect 860 123588 193171 123820
rect 800 123148 193171 123588
rect 860 122916 193171 123148
rect 800 122476 193171 122916
rect 860 122244 193171 122476
rect 800 121804 193171 122244
rect 860 121572 193171 121804
rect 800 121132 193171 121572
rect 860 120900 193171 121132
rect 800 120460 193171 120900
rect 860 120228 193171 120460
rect 800 119788 193171 120228
rect 860 119556 193171 119788
rect 800 119116 193171 119556
rect 860 118884 193171 119116
rect 800 118444 193171 118884
rect 860 118212 193171 118444
rect 800 117772 193171 118212
rect 860 117540 193171 117772
rect 800 117100 193171 117540
rect 860 116868 193171 117100
rect 800 116428 193171 116868
rect 860 116196 193171 116428
rect 800 115756 193171 116196
rect 860 115524 193171 115756
rect 800 115084 193171 115524
rect 860 114852 193171 115084
rect 800 114412 193171 114852
rect 860 114180 193171 114412
rect 800 113740 193171 114180
rect 860 113508 193171 113740
rect 800 113068 193171 113508
rect 860 112836 193171 113068
rect 800 112396 193171 112836
rect 860 112164 193171 112396
rect 800 111724 193171 112164
rect 860 111492 193171 111724
rect 800 111052 193171 111492
rect 860 110820 193171 111052
rect 800 110380 193171 110820
rect 860 110148 193171 110380
rect 800 109708 193171 110148
rect 860 109476 193171 109708
rect 800 109036 193171 109476
rect 860 108804 193171 109036
rect 800 108364 193171 108804
rect 860 108132 193171 108364
rect 800 107692 193171 108132
rect 860 107460 193171 107692
rect 800 107020 193171 107460
rect 860 106788 193171 107020
rect 800 106348 193171 106788
rect 860 106116 193171 106348
rect 800 105676 193171 106116
rect 860 105444 193171 105676
rect 800 105004 193171 105444
rect 860 104772 193171 105004
rect 800 104332 193171 104772
rect 860 104100 193171 104332
rect 800 103660 193171 104100
rect 860 103428 193171 103660
rect 800 102988 193171 103428
rect 860 102756 193171 102988
rect 800 102316 193171 102756
rect 860 102084 193171 102316
rect 800 101644 193171 102084
rect 860 101412 193171 101644
rect 800 100972 193171 101412
rect 860 100740 193171 100972
rect 800 100300 193171 100740
rect 860 100068 193171 100300
rect 800 99628 193171 100068
rect 860 99396 193171 99628
rect 800 98956 193171 99396
rect 860 98724 193171 98956
rect 800 98284 193171 98724
rect 860 98052 193171 98284
rect 800 97612 193171 98052
rect 860 97380 193171 97612
rect 800 96940 193171 97380
rect 860 96708 193171 96940
rect 800 96268 193171 96708
rect 860 96036 193171 96268
rect 800 10924 193171 96036
rect 860 10692 193171 10924
rect 800 9580 193171 10692
rect 860 9348 193171 9580
rect 800 8908 193171 9348
rect 860 8676 193171 8908
rect 800 6892 193171 8676
rect 860 6660 193171 6892
rect 800 6220 193171 6660
rect 860 5988 193171 6220
rect 800 5548 193171 5988
rect 860 5316 193171 5548
rect 800 4876 193171 5316
rect 860 4644 193171 4876
rect 800 4204 193171 4644
rect 860 3972 193171 4204
rect 800 3108 193171 3972
<< metal4 >>
rect 4448 3076 4768 193708
rect 19808 3076 20128 193708
rect 35168 3076 35488 193708
rect 50528 3076 50848 193708
rect 65888 3076 66208 193708
rect 81248 3076 81568 193708
rect 96608 3076 96928 193708
rect 111968 3076 112288 193708
rect 127328 3076 127648 193708
rect 142688 3076 143008 193708
rect 158048 3076 158368 193708
rect 173408 3076 173728 193708
rect 188768 3076 189088 193708
<< obsm4 >>
rect 9660 8306 19748 186238
rect 20188 8306 35108 186238
rect 35548 8306 50468 186238
rect 50908 8306 65828 186238
rect 66268 8306 81188 186238
rect 81628 8306 96548 186238
rect 96988 8306 111908 186238
rect 112348 8306 127268 186238
rect 127708 8306 142628 186238
rect 143068 8306 157988 186238
rect 158428 8306 173348 186238
rect 173788 8306 185444 186238
<< labels >>
rlabel metal3 s 0 184128 800 184240 6 i_clk
port 1 nsew signal input
rlabel metal3 s 0 96768 800 96880 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 0 97440 800 97552 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal3 s 0 100128 800 100240 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal3 s 0 100800 800 100912 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal3 s 0 110208 800 110320 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal3 s 0 110880 800 110992 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal3 s 0 112224 800 112336 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal3 s 0 114912 800 115024 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal3 s 0 112896 800 113008 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal3 s 0 134400 800 134512 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal3 s 0 132384 800 132496 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 0 144480 800 144592 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 0 137760 800 137872 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 0 143808 800 143920 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 0 143136 800 143248 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 0 137088 800 137200 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 0 136416 800 136528 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 0 135744 800 135856 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 0 135072 800 135184 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 0 133056 800 133168 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 0 133728 800 133840 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 0 118272 800 118384 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 0 118944 800 119056 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal3 s 0 122976 800 123088 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 0 131712 800 131824 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 0 127008 800 127120 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 0 124320 800 124432 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 0 129696 800 129808 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 0 125664 800 125776 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 0 130368 800 130480 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 0 123648 800 123760 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 0 124992 800 125104 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal3 s 0 122304 800 122416 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal3 s 0 99456 800 99568 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal3 s 0 106848 800 106960 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 0 104832 800 104944 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal3 s 0 108192 800 108304 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 0 106176 800 106288 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 0 108864 800 108976 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 0 0 112 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal2 s 50400 0 50512 800 6 i_mode[0]
port 42 nsew signal input
rlabel metal2 s 51072 0 51184 800 6 i_mode[1]
port 43 nsew signal input
rlabel metal2 s 121632 196755 121744 197555 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 0 141120 800 141232 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 0 142464 800 142576 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 0 101472 800 101584 6 i_reg_outs_enb
port 47 nsew signal input
rlabel metal3 s 0 141792 800 141904 6 i_reg_sclk
port 48 nsew signal input
rlabel metal3 s 0 107520 800 107632 6 i_reset_lock_a
port 49 nsew signal input
rlabel metal3 s 0 104160 800 104272 6 i_reset_lock_b
port 50 nsew signal input
rlabel metal2 s 672 0 784 800 6 i_spare_0
port 51 nsew signal input
rlabel metal2 s 1344 0 1456 800 6 i_spare_1
port 52 nsew signal input
rlabel metal3 s 0 140448 800 140560 6 i_test_uc2
port 53 nsew signal input
rlabel metal3 s 0 139104 800 139216 6 i_test_wci
port 54 nsew signal input
rlabel metal3 s 0 98784 800 98896 6 i_tex_in[0]
port 55 nsew signal input
rlabel metal3 s 0 111552 800 111664 6 i_tex_in[1]
port 56 nsew signal input
rlabel metal3 s 0 138432 800 138544 6 i_tex_in[2]
port 57 nsew signal input
rlabel metal3 s 0 116256 800 116368 6 i_tex_in[3]
port 58 nsew signal input
rlabel metal3 s 0 115584 800 115696 6 i_vec_csb
port 59 nsew signal input
rlabel metal3 s 0 139776 800 139888 6 i_vec_mosi
port 60 nsew signal input
rlabel metal3 s 0 116928 800 117040 6 i_vec_sclk
port 61 nsew signal input
rlabel metal3 s 0 113568 800 113680 6 o_gpout[0]
port 62 nsew signal output
rlabel metal3 s 0 114240 800 114352 6 o_gpout[1]
port 63 nsew signal output
rlabel metal3 s 0 131040 800 131152 6 o_gpout[2]
port 64 nsew signal output
rlabel metal3 s 0 126336 800 126448 6 o_gpout[3]
port 65 nsew signal output
rlabel metal3 s 0 129024 800 129136 6 o_gpout[4]
port 66 nsew signal output
rlabel metal3 s 0 102144 800 102256 6 o_gpout[5]
port 67 nsew signal output
rlabel metal3 s 0 105504 800 105616 6 o_hsync
port 68 nsew signal output
rlabel metal3 s 0 96096 800 96208 6 o_reset
port 69 nsew signal output
rlabel metal2 s 55776 0 55888 800 6 o_rgb[0]
port 70 nsew signal output
rlabel metal2 s 92736 0 92848 800 6 o_rgb[10]
port 71 nsew signal output
rlabel metal2 s 154560 196755 154672 197555 6 o_rgb[11]
port 72 nsew signal output
rlabel metal2 s 168672 0 168784 800 6 o_rgb[12]
port 73 nsew signal output
rlabel metal2 s 134400 196755 134512 197555 6 o_rgb[13]
port 74 nsew signal output
rlabel metal3 s 0 109536 800 109648 6 o_rgb[14]
port 75 nsew signal output
rlabel metal3 s 0 128352 800 128464 6 o_rgb[15]
port 76 nsew signal output
rlabel metal2 s 185472 0 185584 800 6 o_rgb[16]
port 77 nsew signal output
rlabel metal2 s 112224 0 112336 800 6 o_rgb[17]
port 78 nsew signal output
rlabel metal2 s 166656 196755 166768 197555 6 o_rgb[18]
port 79 nsew signal output
rlabel metal2 s 110880 0 110992 800 6 o_rgb[19]
port 80 nsew signal output
rlabel metal3 s 193171 171360 193971 171472 6 o_rgb[1]
port 81 nsew signal output
rlabel metal3 s 193171 191520 193971 191632 6 o_rgb[20]
port 82 nsew signal output
rlabel metal2 s 159264 0 159376 800 6 o_rgb[21]
port 83 nsew signal output
rlabel metal3 s 0 127680 800 127792 6 o_rgb[22]
port 84 nsew signal output
rlabel metal3 s 0 102816 800 102928 6 o_rgb[23]
port 85 nsew signal output
rlabel metal2 s 36288 196755 36400 197555 6 o_rgb[2]
port 86 nsew signal output
rlabel metal2 s 2688 196755 2800 197555 6 o_rgb[3]
port 87 nsew signal output
rlabel metal2 s 186144 0 186256 800 6 o_rgb[4]
port 88 nsew signal output
rlabel metal3 s 0 5376 800 5488 6 o_rgb[5]
port 89 nsew signal output
rlabel metal3 s 0 120960 800 121072 6 o_rgb[6]
port 90 nsew signal output
rlabel metal3 s 0 117600 800 117712 6 o_rgb[7]
port 91 nsew signal output
rlabel metal3 s 0 6720 800 6832 6 o_rgb[8]
port 92 nsew signal output
rlabel metal2 s 183456 0 183568 800 6 o_rgb[9]
port 93 nsew signal output
rlabel metal3 s 0 98112 800 98224 6 o_tex_csb
port 94 nsew signal output
rlabel metal3 s 0 121632 800 121744 6 o_tex_oeb0
port 95 nsew signal output
rlabel metal3 s 0 119616 800 119728 6 o_tex_out0
port 96 nsew signal output
rlabel metal3 s 0 120288 800 120400 6 o_tex_sclk
port 97 nsew signal output
rlabel metal3 s 0 103488 800 103600 6 o_vsync
port 98 nsew signal output
rlabel metal2 s 18144 196755 18256 197555 6 ones[0]
port 99 nsew signal output
rlabel metal3 s 0 4704 800 4816 6 ones[10]
port 100 nsew signal output
rlabel metal2 s 141120 196755 141232 197555 6 ones[11]
port 101 nsew signal output
rlabel metal2 s 161280 0 161392 800 6 ones[12]
port 102 nsew signal output
rlabel metal2 s 190848 0 190960 800 6 ones[13]
port 103 nsew signal output
rlabel metal3 s 0 8736 800 8848 6 ones[14]
port 104 nsew signal output
rlabel metal3 s 0 9408 800 9520 6 ones[15]
port 105 nsew signal output
rlabel metal3 s 193171 193536 193971 193648 6 ones[1]
port 106 nsew signal output
rlabel metal3 s 0 4032 800 4144 6 ones[2]
port 107 nsew signal output
rlabel metal2 s 181440 0 181552 800 6 ones[3]
port 108 nsew signal output
rlabel metal2 s 22176 196755 22288 197555 6 ones[4]
port 109 nsew signal output
rlabel metal2 s 137760 196755 137872 197555 6 ones[5]
port 110 nsew signal output
rlabel metal3 s 193171 190848 193971 190960 6 ones[6]
port 111 nsew signal output
rlabel metal3 s 0 6048 800 6160 6 ones[7]
port 112 nsew signal output
rlabel metal2 s 83328 0 83440 800 6 ones[8]
port 113 nsew signal output
rlabel metal2 s 26208 0 26320 800 6 ones[9]
port 114 nsew signal output
rlabel metal4 s 4448 3076 4768 193708 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 193708 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 193708 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 193708 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 193708 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 193708 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 193708 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 193708 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 193708 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 193708 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 193708 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 193708 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 193708 6 vss
port 116 nsew ground bidirectional
rlabel metal3 s 193171 192192 193971 192304 6 zeros[0]
port 117 nsew signal output
rlabel metal2 s 170016 0 170128 800 6 zeros[10]
port 118 nsew signal output
rlabel metal2 s 142464 196755 142576 197555 6 zeros[11]
port 119 nsew signal output
rlabel metal2 s 155232 196755 155344 197555 6 zeros[12]
port 120 nsew signal output
rlabel metal2 s 126336 196755 126448 197555 6 zeros[13]
port 121 nsew signal output
rlabel metal2 s 114912 0 115024 800 6 zeros[14]
port 122 nsew signal output
rlabel metal3 s 193171 192864 193971 192976 6 zeros[15]
port 123 nsew signal output
rlabel metal2 s 148512 196755 148624 197555 6 zeros[1]
port 124 nsew signal output
rlabel metal2 s 153888 196755 154000 197555 6 zeros[2]
port 125 nsew signal output
rlabel metal2 s 52416 0 52528 800 6 zeros[3]
port 126 nsew signal output
rlabel metal2 s 134400 0 134512 800 6 zeros[4]
port 127 nsew signal output
rlabel metal2 s 133728 196755 133840 197555 6 zeros[5]
port 128 nsew signal output
rlabel metal3 s 193171 188832 193971 188944 6 zeros[6]
port 129 nsew signal output
rlabel metal2 s 157920 196755 158032 197555 6 zeros[7]
port 130 nsew signal output
rlabel metal3 s 0 10752 800 10864 6 zeros[8]
port 131 nsew signal output
rlabel metal2 s 188832 0 188944 800 6 zeros[9]
port 132 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 193971 197555
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 26733236
string GDS_FILE /home/zerotoasic/anton/algofoogle-multi-caravel/openlane/top_ew_algofoogle/runs/23_12_01_16_32/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 614794
<< end >>

