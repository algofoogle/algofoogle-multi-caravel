magic
tech gf180mcuD
magscale 1 10
timestamp 1702352917
<< nwell >>
rect 1258 232441 231142 232934
rect 1258 232416 143661 232441
rect 1258 231687 19341 231712
rect 1258 230873 231142 231687
rect 1258 230848 40509 230873
rect 1258 230119 44653 230144
rect 1258 229305 231142 230119
rect 1258 229280 17549 229305
rect 1258 228551 68552 228576
rect 1258 227737 231142 228551
rect 1258 227712 23261 227737
rect 1258 226983 27405 227008
rect 1258 226169 231142 226983
rect 1258 226144 17213 226169
rect 1258 225415 13629 225440
rect 1258 224601 231142 225415
rect 1258 224576 22141 224601
rect 1258 223847 28301 223872
rect 1258 223033 231142 223847
rect 1258 223008 34349 223033
rect 1258 222279 13965 222304
rect 1258 221467 231142 222279
rect 1258 221465 79872 221467
rect 1258 221440 23192 221465
rect 1258 220711 43421 220736
rect 1258 220709 92416 220711
rect 1258 219897 231142 220709
rect 1258 219872 26509 219897
rect 1258 219143 35469 219168
rect 1258 219141 83680 219143
rect 1258 218331 231142 219141
rect 1258 218329 89392 218331
rect 1258 218304 15645 218329
rect 1258 217575 12061 217600
rect 1258 217573 84128 217575
rect 1258 216763 231142 217573
rect 1258 216761 78864 216763
rect 1258 216736 35400 216761
rect 1258 216007 29240 216032
rect 1258 216005 90400 216007
rect 1258 215195 231142 216005
rect 1258 215193 87264 215195
rect 1258 215168 17437 215193
rect 1258 214439 13629 214464
rect 1258 214437 76848 214439
rect 1258 213625 231142 214437
rect 1258 213600 25277 213625
rect 1258 212871 29645 212896
rect 1258 212059 231142 212871
rect 1258 212057 77968 212059
rect 1258 212032 37821 212057
rect 1258 211303 13448 211328
rect 1258 211301 81888 211303
rect 1258 210489 231142 211301
rect 1258 210464 16205 210489
rect 1258 209735 29352 209760
rect 1258 209733 77856 209735
rect 1258 208921 231142 209733
rect 1258 208896 40621 208921
rect 1258 208167 14189 208192
rect 1258 208165 76960 208167
rect 1258 207353 231142 208165
rect 1258 207328 18221 207353
rect 1258 206599 27405 206624
rect 1258 205785 231142 206599
rect 1258 205760 51202 205785
rect 1258 205031 83853 205056
rect 1258 204217 231142 205031
rect 1258 204192 16765 204217
rect 1258 203463 12845 203488
rect 1258 202649 231142 203463
rect 1258 202624 47341 202649
rect 1258 201895 12216 201920
rect 1258 201081 231142 201895
rect 1258 201056 22813 201081
rect 1258 200327 14637 200352
rect 1258 199513 231142 200327
rect 1258 199488 66760 199513
rect 1258 198759 14749 198784
rect 1258 197945 231142 198759
rect 1258 197920 47901 197945
rect 1258 197191 28008 197216
rect 1258 196377 231142 197191
rect 1258 196352 16472 196377
rect 1258 195623 53949 195648
rect 1258 194809 231142 195623
rect 1258 194784 92701 194809
rect 1258 194055 19901 194080
rect 1258 193241 231142 194055
rect 1258 193216 24045 193241
rect 1258 192487 28749 192512
rect 1258 191673 231142 192487
rect 1258 191648 47117 191673
rect 1258 190919 43309 190944
rect 1258 190105 231142 190919
rect 1258 190080 23821 190105
rect 1258 189351 20237 189376
rect 1258 188537 231142 189351
rect 1258 188512 49805 188537
rect 1258 187783 57421 187808
rect 1258 186969 231142 187783
rect 1258 186944 22925 186969
rect 1258 186215 43757 186240
rect 1258 185401 231142 186215
rect 1258 185376 48392 185401
rect 1258 184647 51528 184672
rect 1258 183833 231142 184647
rect 1258 183808 38717 183833
rect 1258 183079 59325 183104
rect 1258 182265 231142 183079
rect 1258 182240 42189 182265
rect 1258 181511 74025 181536
rect 1258 180697 231142 181511
rect 1258 180672 37821 180697
rect 1258 179943 52381 179968
rect 1258 179129 231142 179943
rect 1258 179104 73913 179129
rect 1258 178375 42189 178400
rect 1258 177561 231142 178375
rect 1258 177536 39053 177561
rect 1258 176807 36072 176832
rect 1258 175993 231142 176807
rect 1258 175968 63917 175993
rect 1258 175239 45256 175264
rect 1258 174425 231142 175239
rect 1258 174400 48616 174425
rect 1258 173671 35469 173696
rect 1258 172857 231142 173671
rect 1258 172832 39949 172857
rect 1258 172103 35245 172128
rect 1258 171289 231142 172103
rect 1258 171264 48349 171289
rect 1258 170535 45704 170560
rect 1258 169721 231142 170535
rect 1258 169696 55293 169721
rect 1258 168967 35693 168992
rect 1258 168153 231142 168967
rect 1258 168128 33720 168153
rect 1258 167399 47160 167424
rect 1258 166585 231142 167399
rect 1258 166560 39837 166585
rect 1258 165831 43645 165856
rect 1258 165017 231142 165831
rect 1258 164992 40201 165017
rect 1258 164263 30429 164288
rect 1258 163449 231142 164263
rect 1258 163424 51080 163449
rect 1258 162695 38745 162720
rect 1258 161881 231142 162695
rect 1258 161856 40201 161881
rect 1258 161127 19789 161152
rect 1258 160313 231142 161127
rect 1258 160288 104728 160313
rect 1258 159559 43683 159584
rect 1258 158745 231142 159559
rect 1258 158720 23485 158745
rect 1258 157991 19229 158016
rect 1258 157177 231142 157991
rect 1258 157152 49497 157177
rect 1258 156423 53725 156448
rect 1258 155609 231142 156423
rect 1258 155584 14525 155609
rect 1258 154855 33901 154880
rect 1258 154041 231142 154855
rect 1258 154016 18557 154041
rect 1258 153287 13741 153312
rect 1258 152473 231142 153287
rect 1258 152448 8925 152473
rect 1258 151719 82397 151744
rect 1258 150905 231142 151719
rect 1258 150880 29981 150905
rect 1258 150151 4893 150176
rect 1258 149337 231142 150151
rect 1258 149312 69181 149337
rect 1258 148583 35960 148608
rect 1258 147769 231142 148583
rect 1258 147744 2541 147769
rect 1258 147015 19677 147040
rect 1258 146201 231142 147015
rect 1258 146176 62044 146201
rect 1258 145447 69784 145472
rect 1258 144633 231142 145447
rect 1258 144608 2541 144633
rect 1258 143879 21581 143904
rect 1258 143065 231142 143879
rect 1258 143040 32445 143065
rect 1258 142311 53165 142336
rect 1258 141497 231142 142311
rect 1258 141472 2541 141497
rect 1258 140743 12957 140768
rect 1258 139929 231142 140743
rect 1258 139904 46781 139929
rect 1258 139175 44696 139200
rect 1258 138361 231142 139175
rect 1258 138336 2541 138361
rect 1258 137607 36925 137632
rect 1258 136793 231142 137607
rect 1258 136768 18109 136793
rect 1258 136039 10829 136064
rect 1258 135225 231142 136039
rect 1258 135200 2541 135225
rect 1258 134471 6349 134496
rect 1258 133657 231142 134471
rect 1258 133632 10829 133657
rect 1258 132903 20125 132928
rect 1258 132089 231142 132903
rect 1258 132064 2541 132089
rect 1258 131335 36826 131360
rect 1258 130521 231142 131335
rect 1258 130496 7805 130521
rect 1258 129767 20125 129792
rect 1258 128953 231142 129767
rect 1258 128928 2541 128953
rect 1258 128199 5677 128224
rect 1258 127385 231142 128199
rect 1258 127360 10045 127385
rect 1258 126631 13293 126656
rect 1258 125817 231142 126631
rect 1258 125792 2541 125817
rect 1258 125063 6573 125088
rect 1258 124249 231142 125063
rect 1258 124224 38866 124249
rect 1258 123495 10531 123520
rect 1258 122681 231142 123495
rect 1258 122656 2541 122681
rect 1258 121927 10195 121952
rect 1258 121113 231142 121927
rect 1258 121088 8072 121113
rect 1258 120359 19901 120384
rect 1258 119545 231142 120359
rect 1258 119520 2541 119545
rect 1258 118791 12173 118816
rect 1258 117977 231142 118791
rect 1258 117952 25837 117977
rect 1258 117223 2541 117248
rect 1258 116409 231142 117223
rect 1258 116384 69181 116409
rect 1258 115655 12509 115680
rect 1258 114841 231142 115655
rect 1258 114816 56413 114841
rect 1258 114087 2541 114112
rect 1258 113273 231142 114087
rect 1258 113248 10760 113273
rect 1258 112519 12957 112544
rect 1258 111705 231142 112519
rect 1258 111680 16429 111705
rect 1258 110951 5453 110976
rect 1258 110137 231142 110951
rect 1258 110112 2541 110137
rect 1258 109383 12845 109408
rect 1258 108569 231142 109383
rect 1258 108544 19143 108569
rect 1258 107815 43128 107840
rect 1258 107001 231142 107815
rect 1258 106976 2541 107001
rect 1258 106247 10605 106272
rect 1258 105433 231142 106247
rect 1258 105408 15111 105433
rect 1258 104679 6909 104704
rect 1258 103865 231142 104679
rect 1258 103840 2541 103865
rect 1258 103111 57421 103136
rect 1258 102297 231142 103111
rect 1258 102272 14301 102297
rect 1258 101543 6909 101568
rect 1258 100729 231142 101543
rect 1258 100704 30093 100729
rect 1258 99975 2541 100000
rect 1258 99161 231142 99975
rect 1258 99136 80874 99161
rect 1258 98407 10829 98432
rect 1258 97593 231142 98407
rect 1258 97568 7021 97593
rect 1258 96839 2541 96864
rect 1258 96025 231142 96839
rect 1258 96000 26397 96025
rect 1258 95271 12621 95296
rect 1258 94457 231142 95271
rect 1258 94432 9149 94457
rect 1258 93703 4893 93728
rect 1258 92889 231142 93703
rect 1258 92864 25613 92889
rect 1258 92135 12509 92160
rect 1258 91321 231142 92135
rect 1258 91296 6685 91321
rect 1258 90567 2877 90592
rect 1258 89753 231142 90567
rect 1258 89728 15981 89753
rect 1258 88999 10381 89024
rect 1258 88185 231142 88999
rect 1258 88160 6461 88185
rect 1258 87431 34237 87456
rect 1258 86617 231142 87431
rect 1258 86592 114101 86617
rect 1258 85863 2541 85888
rect 1258 85049 231142 85863
rect 1258 85024 61677 85049
rect 1258 84295 6237 84320
rect 1258 83481 231142 84295
rect 1258 83456 14301 83481
rect 1258 82727 2541 82752
rect 1258 81913 231142 82727
rect 1258 81888 11320 81913
rect 1258 81159 49581 81184
rect 1258 80345 231142 81159
rect 1258 80320 14301 80345
rect 1258 79591 5229 79616
rect 1258 78777 231142 79591
rect 1258 78752 61789 78777
rect 1258 78023 74333 78048
rect 1258 77209 231142 78023
rect 1258 77184 9037 77209
rect 1258 76455 4781 76480
rect 1258 75641 231142 76455
rect 1258 75616 40328 75641
rect 1258 74887 6685 74912
rect 1258 74073 231142 74887
rect 1258 74048 10381 74073
rect 1258 73319 13965 73344
rect 1258 72505 231142 73319
rect 1258 72480 77693 72505
rect 1258 71751 10381 71776
rect 1258 70937 231142 71751
rect 1258 70912 25501 70937
rect 1258 70183 44765 70208
rect 1258 69369 231142 70183
rect 1258 69344 14525 69369
rect 1258 68615 100541 68640
rect 1258 67801 231142 68615
rect 1258 67776 9933 67801
rect 1258 67047 29309 67072
rect 1258 66233 231142 67047
rect 1258 66208 15533 66233
rect 1258 65479 21021 65504
rect 1258 64665 231142 65479
rect 1258 64640 10045 64665
rect 1258 63911 34797 63936
rect 1258 63097 231142 63911
rect 1258 63072 26061 63097
rect 1258 62343 11837 62368
rect 1258 61529 231142 62343
rect 1258 61504 87437 61529
rect 1258 60775 14749 60800
rect 1258 59961 231142 60775
rect 1258 59936 25613 59961
rect 1258 59207 41741 59232
rect 1258 58393 231142 59207
rect 1258 58368 22141 58393
rect 1258 57639 14637 57664
rect 1258 56825 231142 57639
rect 1258 56800 32557 56825
rect 1258 56071 27405 56096
rect 1258 55257 231142 56071
rect 1258 55232 19720 55257
rect 1258 54503 14749 54528
rect 1258 53689 231142 54503
rect 1258 53664 37821 53689
rect 1258 52935 28189 52960
rect 1258 52121 231142 52935
rect 1258 52096 24381 52121
rect 1258 51367 67837 51392
rect 1258 50553 231142 51367
rect 1258 50528 18040 50553
rect 1258 49799 20685 49824
rect 1258 48985 231142 49799
rect 1258 48960 24717 48985
rect 1258 48231 37080 48256
rect 1258 47417 231142 48231
rect 1258 47392 19048 47417
rect 1258 46663 28861 46688
rect 1258 45849 231142 46663
rect 1258 45824 33608 45849
rect 1258 45095 50632 45120
rect 1258 44281 231142 45095
rect 1258 44256 81193 44281
rect 1258 43527 69095 43552
rect 1258 42713 231142 43527
rect 1258 42688 33005 42713
rect 1258 41959 42637 41984
rect 1258 41145 231142 41959
rect 1258 41120 95320 41145
rect 1258 40391 65261 40416
rect 1258 39577 231142 40391
rect 1258 39552 32781 39577
rect 1258 38823 39320 38848
rect 1258 38009 231142 38823
rect 1258 37984 72248 38009
rect 1258 37255 59997 37280
rect 1258 36441 231142 37255
rect 1258 36416 34349 36441
rect 1258 35687 38269 35712
rect 1258 34873 231142 35687
rect 1258 34848 47677 34873
rect 1258 34119 108829 34144
rect 1258 33305 231142 34119
rect 1258 33280 78072 33305
rect 1258 32551 52045 32576
rect 1258 31737 231142 32551
rect 1258 31712 37933 31737
rect 1258 30983 45592 31008
rect 1258 30169 231142 30983
rect 1258 30144 65709 30169
rect 1258 29415 99309 29440
rect 1258 28601 231142 29415
rect 1258 28576 40845 28601
rect 1258 27847 44317 27872
rect 1258 27033 231142 27847
rect 1258 27008 47677 27033
rect 1258 26279 66829 26304
rect 1258 25465 231142 26279
rect 1258 25440 55657 25465
rect 1258 24711 42189 24736
rect 1258 23897 231142 24711
rect 1258 23872 47677 23897
rect 1258 23143 58541 23168
rect 1258 22329 231142 23143
rect 1258 22304 45661 22329
rect 1258 21575 52045 21600
rect 1258 20761 231142 21575
rect 1258 20736 48573 20761
rect 1258 20007 108200 20032
rect 1258 19193 231142 20007
rect 1258 19168 65261 19193
rect 1258 18439 53501 18464
rect 1258 17625 231142 18439
rect 1258 17600 89229 17625
rect 1258 16871 137165 16896
rect 1258 16057 231142 16871
rect 1258 16032 85309 16057
rect 1258 15303 67949 15328
rect 1258 14489 231142 15303
rect 1258 14464 71421 14489
rect 1258 13735 85785 13760
rect 1258 12921 231142 13735
rect 1258 12896 141900 12921
rect 1258 12167 75901 12192
rect 1258 11353 231142 12167
rect 1258 11328 72093 11353
rect 1258 10599 82957 10624
rect 1258 9785 231142 10599
rect 1258 9760 97896 9785
rect 1258 9031 114093 9056
rect 1258 8217 231142 9031
rect 1258 8192 72989 8217
rect 1258 7463 91469 7488
rect 1258 6649 231142 7463
rect 1258 6624 84861 6649
rect 1258 5895 161848 5920
rect 1258 5081 231142 5895
rect 1258 5056 87032 5081
rect 1258 4327 82061 4352
rect 1258 3513 231142 4327
rect 1258 3488 155197 3513
<< pwell >>
rect 1258 231712 231142 232416
rect 1258 230144 231142 230848
rect 1258 228576 231142 229280
rect 1258 227008 231142 227712
rect 1258 225440 231142 226144
rect 1258 223872 231142 224576
rect 1258 222304 231142 223008
rect 1258 220736 231142 221440
rect 1258 219168 231142 219872
rect 1258 217600 231142 218304
rect 1258 216032 231142 216736
rect 1258 214464 231142 215168
rect 1258 212896 231142 213600
rect 1258 211328 231142 212032
rect 1258 209760 231142 210464
rect 1258 208192 231142 208896
rect 1258 206624 231142 207328
rect 1258 205056 231142 205760
rect 1258 203488 231142 204192
rect 1258 201920 231142 202624
rect 1258 200352 231142 201056
rect 1258 198784 231142 199488
rect 1258 197216 231142 197920
rect 1258 195648 231142 196352
rect 1258 194080 231142 194784
rect 1258 192512 231142 193216
rect 1258 190944 231142 191648
rect 1258 189376 231142 190080
rect 1258 187808 231142 188512
rect 1258 186240 231142 186944
rect 1258 184672 231142 185376
rect 1258 183104 231142 183808
rect 1258 181536 231142 182240
rect 1258 179968 231142 180672
rect 1258 178400 231142 179104
rect 1258 176832 231142 177536
rect 1258 175264 231142 175968
rect 1258 173696 231142 174400
rect 1258 172128 231142 172832
rect 1258 170560 231142 171264
rect 1258 168992 231142 169696
rect 1258 167424 231142 168128
rect 1258 165856 231142 166560
rect 1258 164288 231142 164992
rect 1258 162720 231142 163424
rect 1258 161152 231142 161856
rect 1258 159584 231142 160288
rect 1258 158016 231142 158720
rect 1258 156448 231142 157152
rect 1258 154880 231142 155584
rect 1258 153312 231142 154016
rect 1258 151744 231142 152448
rect 1258 150176 231142 150880
rect 1258 148608 231142 149312
rect 1258 147040 231142 147744
rect 1258 145472 231142 146176
rect 1258 143904 231142 144608
rect 1258 142336 231142 143040
rect 1258 140768 231142 141472
rect 1258 139200 231142 139904
rect 1258 137632 231142 138336
rect 1258 136064 231142 136768
rect 1258 134496 231142 135200
rect 1258 132928 231142 133632
rect 1258 131360 231142 132064
rect 1258 129792 231142 130496
rect 1258 128224 231142 128928
rect 1258 126656 231142 127360
rect 1258 125088 231142 125792
rect 1258 123520 231142 124224
rect 1258 121952 231142 122656
rect 1258 120384 231142 121088
rect 1258 118816 231142 119520
rect 1258 117248 231142 117952
rect 1258 115680 231142 116384
rect 1258 114112 231142 114816
rect 1258 112544 231142 113248
rect 1258 110976 231142 111680
rect 1258 109408 231142 110112
rect 1258 107840 231142 108544
rect 1258 106272 231142 106976
rect 1258 104704 231142 105408
rect 1258 103136 231142 103840
rect 1258 101568 231142 102272
rect 1258 100000 231142 100704
rect 1258 98432 231142 99136
rect 1258 96864 231142 97568
rect 1258 95296 231142 96000
rect 1258 93728 231142 94432
rect 1258 92160 231142 92864
rect 1258 90592 231142 91296
rect 1258 89024 231142 89728
rect 1258 87456 231142 88160
rect 1258 85888 231142 86592
rect 1258 84320 231142 85024
rect 1258 82752 231142 83456
rect 1258 81184 231142 81888
rect 1258 79616 231142 80320
rect 1258 78048 231142 78752
rect 1258 76480 231142 77184
rect 1258 74912 231142 75616
rect 1258 73344 231142 74048
rect 1258 71776 231142 72480
rect 1258 70208 231142 70912
rect 1258 68640 231142 69344
rect 1258 67072 231142 67776
rect 1258 65504 231142 66208
rect 1258 63936 231142 64640
rect 1258 62368 231142 63072
rect 1258 60800 231142 61504
rect 1258 59232 231142 59936
rect 1258 57664 231142 58368
rect 1258 56096 231142 56800
rect 1258 54528 231142 55232
rect 1258 52960 231142 53664
rect 1258 51392 231142 52096
rect 1258 49824 231142 50528
rect 1258 48256 231142 48960
rect 1258 46688 231142 47392
rect 1258 45120 231142 45824
rect 1258 43552 231142 44256
rect 1258 41984 231142 42688
rect 1258 40416 231142 41120
rect 1258 38848 231142 39552
rect 1258 37280 231142 37984
rect 1258 35712 231142 36416
rect 1258 34144 231142 34848
rect 1258 32576 231142 33280
rect 1258 31008 231142 31712
rect 1258 29440 231142 30144
rect 1258 27872 231142 28576
rect 1258 26304 231142 27008
rect 1258 24736 231142 25440
rect 1258 23168 231142 23872
rect 1258 21600 231142 22304
rect 1258 20032 231142 20736
rect 1258 18464 231142 19168
rect 1258 16896 231142 17600
rect 1258 15328 231142 16032
rect 1258 13760 231142 14464
rect 1258 12192 231142 12896
rect 1258 10624 231142 11328
rect 1258 9056 231142 9760
rect 1258 7488 231142 8192
rect 1258 5920 231142 6624
rect 1258 4352 231142 5056
rect 1258 3050 231142 3488
<< obsm1 >>
rect 1344 3076 231056 233490
<< metal2 >>
rect 6272 235248 6384 236048
rect 12992 235248 13104 236048
rect 15232 235248 15344 236048
rect 17472 235248 17584 236048
rect 19712 235248 19824 236048
rect 21952 235248 22064 236048
rect 24192 235248 24304 236048
rect 26432 235248 26544 236048
rect 28672 235248 28784 236048
rect 30912 235248 31024 236048
rect 33152 235248 33264 236048
rect 35392 235248 35504 236048
rect 37632 235248 37744 236048
rect 39872 235248 39984 236048
rect 42112 235248 42224 236048
rect 44352 235248 44464 236048
rect 46592 235248 46704 236048
rect 48832 235248 48944 236048
rect 51072 235248 51184 236048
rect 53312 235248 53424 236048
rect 55552 235248 55664 236048
rect 57792 235248 57904 236048
rect 60032 235248 60144 236048
rect 62272 235248 62384 236048
rect 64512 235248 64624 236048
rect 66752 235248 66864 236048
rect 68992 235248 69104 236048
rect 71232 235248 71344 236048
rect 73472 235248 73584 236048
rect 75712 235248 75824 236048
rect 77952 235248 78064 236048
rect 80192 235248 80304 236048
rect 82432 235248 82544 236048
rect 84672 235248 84784 236048
rect 86912 235248 87024 236048
rect 89152 235248 89264 236048
rect 91392 235248 91504 236048
rect 93632 235248 93744 236048
rect 95872 235248 95984 236048
rect 98112 235248 98224 236048
rect 100352 235248 100464 236048
rect 102592 235248 102704 236048
rect 104832 235248 104944 236048
rect 107072 235248 107184 236048
rect 109312 235248 109424 236048
rect 111552 235248 111664 236048
rect 113792 235248 113904 236048
rect 116032 235248 116144 236048
rect 118272 235248 118384 236048
rect 120512 235248 120624 236048
rect 122752 235248 122864 236048
rect 124992 235248 125104 236048
rect 127232 235248 127344 236048
rect 129472 235248 129584 236048
rect 131712 235248 131824 236048
rect 133952 235248 134064 236048
rect 136192 235248 136304 236048
rect 138432 235248 138544 236048
rect 140672 235248 140784 236048
rect 142912 235248 143024 236048
rect 145152 235248 145264 236048
rect 147392 235248 147504 236048
rect 149632 235248 149744 236048
rect 151872 235248 151984 236048
rect 154112 235248 154224 236048
rect 156352 235248 156464 236048
rect 158592 235248 158704 236048
rect 160832 235248 160944 236048
rect 163072 235248 163184 236048
rect 165312 235248 165424 236048
rect 167552 235248 167664 236048
rect 169792 235248 169904 236048
rect 172032 235248 172144 236048
rect 174272 235248 174384 236048
rect 176512 235248 176624 236048
rect 178752 235248 178864 236048
rect 180992 235248 181104 236048
rect 183232 235248 183344 236048
rect 185472 235248 185584 236048
rect 187712 235248 187824 236048
rect 189952 235248 190064 236048
rect 192192 235248 192304 236048
rect 194432 235248 194544 236048
rect 196672 235248 196784 236048
rect 198912 235248 199024 236048
rect 201152 235248 201264 236048
rect 203392 235248 203504 236048
rect 205632 235248 205744 236048
rect 207872 235248 207984 236048
rect 210112 235248 210224 236048
rect 212352 235248 212464 236048
rect 214592 235248 214704 236048
rect 216832 235248 216944 236048
rect 219072 235248 219184 236048
rect 221312 235248 221424 236048
rect 223552 235248 223664 236048
rect 225792 235248 225904 236048
<< obsm2 >>
rect 1596 235188 6212 235396
rect 6444 235188 12932 235396
rect 13164 235188 15172 235396
rect 15404 235188 17412 235396
rect 17644 235188 19652 235396
rect 19884 235188 21892 235396
rect 22124 235188 24132 235396
rect 24364 235188 26372 235396
rect 26604 235188 28612 235396
rect 28844 235188 30852 235396
rect 31084 235188 33092 235396
rect 33324 235188 35332 235396
rect 35564 235188 37572 235396
rect 37804 235188 39812 235396
rect 40044 235188 42052 235396
rect 42284 235188 44292 235396
rect 44524 235188 46532 235396
rect 46764 235188 48772 235396
rect 49004 235188 51012 235396
rect 51244 235188 53252 235396
rect 53484 235188 55492 235396
rect 55724 235188 57732 235396
rect 57964 235188 59972 235396
rect 60204 235188 62212 235396
rect 62444 235188 64452 235396
rect 64684 235188 66692 235396
rect 66924 235188 68932 235396
rect 69164 235188 71172 235396
rect 71404 235188 73412 235396
rect 73644 235188 75652 235396
rect 75884 235188 77892 235396
rect 78124 235188 80132 235396
rect 80364 235188 82372 235396
rect 82604 235188 84612 235396
rect 84844 235188 86852 235396
rect 87084 235188 89092 235396
rect 89324 235188 91332 235396
rect 91564 235188 93572 235396
rect 93804 235188 95812 235396
rect 96044 235188 98052 235396
rect 98284 235188 100292 235396
rect 100524 235188 102532 235396
rect 102764 235188 104772 235396
rect 105004 235188 107012 235396
rect 107244 235188 109252 235396
rect 109484 235188 111492 235396
rect 111724 235188 113732 235396
rect 113964 235188 115972 235396
rect 116204 235188 118212 235396
rect 118444 235188 120452 235396
rect 120684 235188 122692 235396
rect 122924 235188 124932 235396
rect 125164 235188 127172 235396
rect 127404 235188 129412 235396
rect 129644 235188 131652 235396
rect 131884 235188 133892 235396
rect 134124 235188 136132 235396
rect 136364 235188 138372 235396
rect 138604 235188 140612 235396
rect 140844 235188 142852 235396
rect 143084 235188 145092 235396
rect 145324 235188 147332 235396
rect 147564 235188 149572 235396
rect 149804 235188 151812 235396
rect 152044 235188 154052 235396
rect 154284 235188 156292 235396
rect 156524 235188 158532 235396
rect 158764 235188 160772 235396
rect 161004 235188 163012 235396
rect 163244 235188 165252 235396
rect 165484 235188 167492 235396
rect 167724 235188 169732 235396
rect 169964 235188 171972 235396
rect 172204 235188 174212 235396
rect 174444 235188 176452 235396
rect 176684 235188 178692 235396
rect 178924 235188 180932 235396
rect 181164 235188 183172 235396
rect 183404 235188 185412 235396
rect 185644 235188 187652 235396
rect 187884 235188 189892 235396
rect 190124 235188 192132 235396
rect 192364 235188 194372 235396
rect 194604 235188 196612 235396
rect 196844 235188 198852 235396
rect 199084 235188 201092 235396
rect 201324 235188 203332 235396
rect 203564 235188 205572 235396
rect 205804 235188 207812 235396
rect 208044 235188 210052 235396
rect 210284 235188 212292 235396
rect 212524 235188 214532 235396
rect 214764 235188 216772 235396
rect 217004 235188 219012 235396
rect 219244 235188 221252 235396
rect 221484 235188 223492 235396
rect 223724 235188 225732 235396
rect 225964 235188 230692 235396
rect 1596 802 230692 235188
<< obsm3 >>
rect 1586 812 230702 235060
<< metal4 >>
rect 4448 3076 4768 232908
rect 19808 3076 20128 232908
rect 35168 3076 35488 232908
rect 50528 3076 50848 232908
rect 65888 3076 66208 232908
rect 81248 3076 81568 232908
rect 96608 3076 96928 232908
rect 111968 3076 112288 232908
rect 127328 3076 127648 232908
rect 142688 3076 143008 232908
rect 158048 3076 158368 232908
rect 173408 3076 173728 232908
rect 188768 3076 189088 232908
rect 204128 3076 204448 232908
rect 219488 3076 219808 232908
<< obsm4 >>
rect 24220 232968 225764 234622
rect 24220 3016 35108 232968
rect 35548 3016 50468 232968
rect 50908 3016 65828 232968
rect 66268 3016 81188 232968
rect 81628 3016 96548 232968
rect 96988 3016 111908 232968
rect 112348 3016 127268 232968
rect 127708 3016 142628 232968
rect 143068 3016 157988 232968
rect 158428 3016 173348 232968
rect 173788 3016 188708 232968
rect 189148 3016 204068 232968
rect 204508 3016 219428 232968
rect 219868 3016 225764 232968
rect 24220 914 225764 3016
<< labels >>
rlabel metal2 s 156352 235248 156464 236048 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 178752 235248 178864 236048 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 180992 235248 181104 236048 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 183232 235248 183344 236048 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 185472 235248 185584 236048 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 187712 235248 187824 236048 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 189952 235248 190064 236048 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 192192 235248 192304 236048 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 194432 235248 194544 236048 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 196672 235248 196784 236048 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 198912 235248 199024 236048 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 158592 235248 158704 236048 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 201152 235248 201264 236048 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 203392 235248 203504 236048 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 205632 235248 205744 236048 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 207872 235248 207984 236048 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 210112 235248 210224 236048 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 212352 235248 212464 236048 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 214592 235248 214704 236048 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 216832 235248 216944 236048 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 219072 235248 219184 236048 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 221312 235248 221424 236048 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 160832 235248 160944 236048 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 223552 235248 223664 236048 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 225792 235248 225904 236048 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 163072 235248 163184 236048 6 io_in[3]
port 26 nsew signal input
rlabel metal2 s 165312 235248 165424 236048 6 io_in[4]
port 27 nsew signal input
rlabel metal2 s 167552 235248 167664 236048 6 io_in[5]
port 28 nsew signal input
rlabel metal2 s 169792 235248 169904 236048 6 io_in[6]
port 29 nsew signal input
rlabel metal2 s 172032 235248 172144 236048 6 io_in[7]
port 30 nsew signal input
rlabel metal2 s 174272 235248 174384 236048 6 io_in[8]
port 31 nsew signal input
rlabel metal2 s 176512 235248 176624 236048 6 io_in[9]
port 32 nsew signal input
rlabel metal2 s 84672 235248 84784 236048 6 io_oeb[0]
port 33 nsew signal output
rlabel metal2 s 107072 235248 107184 236048 6 io_oeb[10]
port 34 nsew signal output
rlabel metal2 s 109312 235248 109424 236048 6 io_oeb[11]
port 35 nsew signal output
rlabel metal2 s 111552 235248 111664 236048 6 io_oeb[12]
port 36 nsew signal output
rlabel metal2 s 113792 235248 113904 236048 6 io_oeb[13]
port 37 nsew signal output
rlabel metal2 s 116032 235248 116144 236048 6 io_oeb[14]
port 38 nsew signal output
rlabel metal2 s 118272 235248 118384 236048 6 io_oeb[15]
port 39 nsew signal output
rlabel metal2 s 120512 235248 120624 236048 6 io_oeb[16]
port 40 nsew signal output
rlabel metal2 s 122752 235248 122864 236048 6 io_oeb[17]
port 41 nsew signal output
rlabel metal2 s 124992 235248 125104 236048 6 io_oeb[18]
port 42 nsew signal output
rlabel metal2 s 127232 235248 127344 236048 6 io_oeb[19]
port 43 nsew signal output
rlabel metal2 s 86912 235248 87024 236048 6 io_oeb[1]
port 44 nsew signal output
rlabel metal2 s 129472 235248 129584 236048 6 io_oeb[20]
port 45 nsew signal output
rlabel metal2 s 131712 235248 131824 236048 6 io_oeb[21]
port 46 nsew signal output
rlabel metal2 s 133952 235248 134064 236048 6 io_oeb[22]
port 47 nsew signal output
rlabel metal2 s 136192 235248 136304 236048 6 io_oeb[23]
port 48 nsew signal output
rlabel metal2 s 138432 235248 138544 236048 6 io_oeb[24]
port 49 nsew signal output
rlabel metal2 s 140672 235248 140784 236048 6 io_oeb[25]
port 50 nsew signal output
rlabel metal2 s 142912 235248 143024 236048 6 io_oeb[26]
port 51 nsew signal output
rlabel metal2 s 145152 235248 145264 236048 6 io_oeb[27]
port 52 nsew signal output
rlabel metal2 s 147392 235248 147504 236048 6 io_oeb[28]
port 53 nsew signal output
rlabel metal2 s 149632 235248 149744 236048 6 io_oeb[29]
port 54 nsew signal output
rlabel metal2 s 89152 235248 89264 236048 6 io_oeb[2]
port 55 nsew signal output
rlabel metal2 s 151872 235248 151984 236048 6 io_oeb[30]
port 56 nsew signal output
rlabel metal2 s 154112 235248 154224 236048 6 io_oeb[31]
port 57 nsew signal output
rlabel metal2 s 91392 235248 91504 236048 6 io_oeb[3]
port 58 nsew signal output
rlabel metal2 s 93632 235248 93744 236048 6 io_oeb[4]
port 59 nsew signal output
rlabel metal2 s 95872 235248 95984 236048 6 io_oeb[5]
port 60 nsew signal output
rlabel metal2 s 98112 235248 98224 236048 6 io_oeb[6]
port 61 nsew signal output
rlabel metal2 s 100352 235248 100464 236048 6 io_oeb[7]
port 62 nsew signal output
rlabel metal2 s 102592 235248 102704 236048 6 io_oeb[8]
port 63 nsew signal output
rlabel metal2 s 104832 235248 104944 236048 6 io_oeb[9]
port 64 nsew signal output
rlabel metal2 s 12992 235248 13104 236048 6 io_out[0]
port 65 nsew signal output
rlabel metal2 s 35392 235248 35504 236048 6 io_out[10]
port 66 nsew signal output
rlabel metal2 s 37632 235248 37744 236048 6 io_out[11]
port 67 nsew signal output
rlabel metal2 s 39872 235248 39984 236048 6 io_out[12]
port 68 nsew signal output
rlabel metal2 s 42112 235248 42224 236048 6 io_out[13]
port 69 nsew signal output
rlabel metal2 s 44352 235248 44464 236048 6 io_out[14]
port 70 nsew signal output
rlabel metal2 s 46592 235248 46704 236048 6 io_out[15]
port 71 nsew signal output
rlabel metal2 s 48832 235248 48944 236048 6 io_out[16]
port 72 nsew signal output
rlabel metal2 s 51072 235248 51184 236048 6 io_out[17]
port 73 nsew signal output
rlabel metal2 s 53312 235248 53424 236048 6 io_out[18]
port 74 nsew signal output
rlabel metal2 s 55552 235248 55664 236048 6 io_out[19]
port 75 nsew signal output
rlabel metal2 s 15232 235248 15344 236048 6 io_out[1]
port 76 nsew signal output
rlabel metal2 s 57792 235248 57904 236048 6 io_out[20]
port 77 nsew signal output
rlabel metal2 s 60032 235248 60144 236048 6 io_out[21]
port 78 nsew signal output
rlabel metal2 s 62272 235248 62384 236048 6 io_out[22]
port 79 nsew signal output
rlabel metal2 s 64512 235248 64624 236048 6 io_out[23]
port 80 nsew signal output
rlabel metal2 s 66752 235248 66864 236048 6 io_out[24]
port 81 nsew signal output
rlabel metal2 s 68992 235248 69104 236048 6 io_out[25]
port 82 nsew signal output
rlabel metal2 s 71232 235248 71344 236048 6 io_out[26]
port 83 nsew signal output
rlabel metal2 s 73472 235248 73584 236048 6 io_out[27]
port 84 nsew signal output
rlabel metal2 s 75712 235248 75824 236048 6 io_out[28]
port 85 nsew signal output
rlabel metal2 s 77952 235248 78064 236048 6 io_out[29]
port 86 nsew signal output
rlabel metal2 s 17472 235248 17584 236048 6 io_out[2]
port 87 nsew signal output
rlabel metal2 s 80192 235248 80304 236048 6 io_out[30]
port 88 nsew signal output
rlabel metal2 s 82432 235248 82544 236048 6 io_out[31]
port 89 nsew signal output
rlabel metal2 s 19712 235248 19824 236048 6 io_out[3]
port 90 nsew signal output
rlabel metal2 s 21952 235248 22064 236048 6 io_out[4]
port 91 nsew signal output
rlabel metal2 s 24192 235248 24304 236048 6 io_out[5]
port 92 nsew signal output
rlabel metal2 s 26432 235248 26544 236048 6 io_out[6]
port 93 nsew signal output
rlabel metal2 s 28672 235248 28784 236048 6 io_out[7]
port 94 nsew signal output
rlabel metal2 s 30912 235248 31024 236048 6 io_out[8]
port 95 nsew signal output
rlabel metal2 s 33152 235248 33264 236048 6 io_out[9]
port 96 nsew signal output
rlabel metal4 s 4448 3076 4768 232908 6 vdd
port 97 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 232908 6 vdd
port 97 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 232908 6 vdd
port 97 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 232908 6 vdd
port 97 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 232908 6 vdd
port 97 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 232908 6 vdd
port 97 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 232908 6 vdd
port 97 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 232908 6 vdd
port 97 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 232908 6 vss
port 98 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 232908 6 vss
port 98 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 232908 6 vss
port 98 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 232908 6 vss
port 98 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 232908 6 vss
port 98 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 232908 6 vss
port 98 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 232908 6 vss
port 98 nsew ground bidirectional
rlabel metal2 s 6272 235248 6384 236048 6 wb_clk_i
port 99 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 232464 236048
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 33687368
string GDS_FILE /home/zerotoasic/anton/algofoogle-multi-caravel/openlane/user_proj_cpu/runs/23_12_12_14_00/results/signoff/user_proj_cpu.magic.gds
string GDS_START 519820
<< end >>

