VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO asic_hat_logo
  CLASS BLOCK ;
  FOREIGN asic_hat_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 310.500 BY 310.500 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 167.400 296.100 172.800 297.000 ;
        RECT 159.300 295.200 173.700 296.100 ;
        RECT 153.000 294.300 175.500 295.200 ;
        RECT 147.600 293.400 178.200 294.300 ;
        RECT 142.200 292.500 181.800 293.400 ;
        RECT 137.700 291.600 182.700 292.500 ;
        RECT 133.200 290.700 176.400 291.600 ;
        RECT 130.500 289.800 171.900 290.700 ;
        RECT 126.900 288.900 168.300 289.800 ;
        RECT 123.300 288.000 163.800 288.900 ;
        RECT 120.600 287.100 162.000 288.000 ;
        RECT 118.800 286.200 159.300 287.100 ;
        RECT 116.100 285.300 156.600 286.200 ;
        RECT 114.300 284.400 153.900 285.300 ;
        RECT 111.600 283.500 151.200 284.400 ;
        RECT 109.800 282.600 148.500 283.500 ;
        RECT 204.300 282.600 211.500 283.500 ;
        RECT 108.000 281.700 144.900 282.600 ;
        RECT 205.200 281.700 215.100 282.600 ;
        RECT 107.100 280.800 143.100 281.700 ;
        RECT 207.000 280.800 217.800 281.700 ;
        RECT 105.300 279.900 141.300 280.800 ;
        RECT 207.900 279.900 218.700 280.800 ;
        RECT 104.400 279.000 139.500 279.900 ;
        RECT 209.700 279.000 220.500 279.900 ;
        RECT 102.600 278.100 135.900 279.000 ;
        RECT 211.500 278.100 221.400 279.000 ;
        RECT 100.800 277.200 132.300 278.100 ;
        RECT 213.300 277.200 222.300 278.100 ;
        RECT 99.900 276.300 129.600 277.200 ;
        RECT 214.200 276.300 223.200 277.200 ;
        RECT 99.000 275.400 126.900 276.300 ;
        RECT 216.000 275.400 224.100 276.300 ;
        RECT 97.200 274.500 124.200 275.400 ;
        RECT 216.900 274.500 225.000 275.400 ;
        RECT 96.300 273.600 121.500 274.500 ;
        RECT 217.800 273.600 225.900 274.500 ;
        RECT 95.400 272.700 119.700 273.600 ;
        RECT 219.600 272.700 226.800 273.600 ;
        RECT 94.500 271.800 117.900 272.700 ;
        RECT 220.500 271.800 227.700 272.700 ;
        RECT 93.600 270.900 116.100 271.800 ;
        RECT 221.400 270.900 228.600 271.800 ;
        RECT 92.700 270.000 114.300 270.900 ;
        RECT 222.300 270.000 228.600 270.900 ;
        RECT 91.800 269.100 111.600 270.000 ;
        RECT 222.300 269.100 229.500 270.000 ;
        RECT 90.900 268.200 110.700 269.100 ;
        RECT 223.200 268.200 230.400 269.100 ;
        RECT 90.000 267.300 108.900 268.200 ;
        RECT 224.100 267.300 230.400 268.200 ;
        RECT 89.100 266.400 108.000 267.300 ;
        RECT 88.200 265.500 106.200 266.400 ;
        RECT 225.000 265.500 231.300 267.300 ;
        RECT 88.200 264.600 105.300 265.500 ;
        RECT 87.300 263.700 104.400 264.600 ;
        RECT 225.900 263.700 232.200 265.500 ;
        RECT 86.400 262.800 103.500 263.700 ;
        RECT 226.800 262.800 232.200 263.700 ;
        RECT 86.400 261.900 102.600 262.800 ;
        RECT 227.700 261.900 233.100 262.800 ;
        RECT 85.500 261.000 101.700 261.900 ;
        RECT 85.500 260.100 100.800 261.000 ;
        RECT 227.700 260.100 234.000 261.900 ;
        RECT 84.600 259.200 99.900 260.100 ;
        RECT 228.600 259.200 234.000 260.100 ;
        RECT 84.600 258.300 99.000 259.200 ;
        RECT 228.600 258.300 234.900 259.200 ;
        RECT 83.700 257.400 99.000 258.300 ;
        RECT 83.700 256.500 98.100 257.400 ;
        RECT 229.500 256.500 234.900 258.300 ;
        RECT 82.800 254.700 97.200 256.500 ;
        RECT 229.500 254.700 235.800 256.500 ;
        RECT 82.800 253.800 96.300 254.700 ;
        RECT 81.900 252.900 96.300 253.800 ;
        RECT 81.900 252.000 95.400 252.900 ;
        RECT 81.000 251.100 95.400 252.000 ;
        RECT 230.400 252.000 235.800 254.700 ;
        RECT 81.000 250.200 94.500 251.100 ;
        RECT 230.400 250.200 236.700 252.000 ;
        RECT 81.000 248.400 93.600 250.200 ;
        RECT 80.100 247.500 93.600 248.400 ;
        RECT 80.100 245.700 92.700 247.500 ;
        RECT 79.200 243.900 92.700 245.700 ;
        RECT 231.300 244.800 236.700 250.200 ;
        RECT 79.200 242.100 91.800 243.900 ;
        RECT 231.300 243.000 237.600 244.800 ;
        RECT 78.300 241.200 91.800 242.100 ;
        RECT 78.300 237.600 90.900 241.200 ;
        RECT 77.400 236.700 90.900 237.600 ;
        RECT 77.400 234.000 90.000 236.700 ;
        RECT 76.500 230.400 90.000 234.000 ;
        RECT 76.500 226.800 89.100 230.400 ;
        RECT 75.600 224.100 89.100 226.800 ;
        RECT 75.600 215.100 88.200 224.100 ;
        RECT 232.200 223.200 237.600 243.000 ;
        RECT 74.700 213.300 88.200 215.100 ;
        RECT 231.300 220.500 237.600 223.200 ;
        RECT 74.700 176.400 87.300 213.300 ;
        RECT 231.300 210.600 236.700 220.500 ;
        RECT 230.400 208.800 236.700 210.600 ;
        RECT 230.400 201.600 235.800 208.800 ;
        RECT 229.500 199.800 235.800 201.600 ;
        RECT 229.500 193.500 234.900 199.800 ;
        RECT 228.600 191.700 234.900 193.500 ;
        RECT 228.600 185.400 234.000 191.700 ;
        RECT 227.700 183.600 234.000 185.400 ;
        RECT 227.700 178.200 233.100 183.600 ;
        RECT 227.700 176.400 232.200 178.200 ;
        RECT 75.600 173.700 87.300 176.400 ;
        RECT 76.500 171.000 87.300 173.700 ;
        RECT 77.400 168.300 87.300 171.000 ;
        RECT 226.800 168.300 232.200 176.400 ;
        RECT 78.300 165.600 88.200 168.300 ;
        RECT 226.800 167.400 231.300 168.300 ;
        RECT 78.300 164.700 89.100 165.600 ;
        RECT 79.200 163.800 90.000 164.700 ;
        RECT 80.100 162.900 90.000 163.800 ;
        RECT 80.100 162.000 90.900 162.900 ;
        RECT 81.000 161.100 90.900 162.000 ;
        RECT 81.000 160.200 91.800 161.100 ;
        RECT 81.000 159.300 93.600 160.200 ;
        RECT 81.900 158.400 95.400 159.300 ;
        RECT 225.900 158.400 231.300 167.400 ;
        RECT 81.900 157.500 96.300 158.400 ;
        RECT 82.800 156.600 97.200 157.500 ;
        RECT 84.600 155.700 99.900 156.600 ;
        RECT 225.900 155.700 230.400 158.400 ;
        RECT 86.400 154.800 102.600 155.700 ;
        RECT 88.200 153.900 106.200 154.800 ;
        RECT 90.900 153.000 108.900 153.900 ;
        RECT 92.700 152.100 111.600 153.000 ;
        RECT 95.400 151.200 116.100 152.100 ;
        RECT 98.100 150.300 119.700 151.200 ;
        RECT 100.800 149.400 124.200 150.300 ;
        RECT 104.400 148.500 128.700 149.400 ;
        RECT 108.000 147.600 134.100 148.500 ;
        RECT 111.600 146.700 138.600 147.600 ;
        RECT 115.200 145.800 143.100 146.700 ;
        RECT 119.700 144.900 148.500 145.800 ;
        RECT 123.300 144.000 153.900 144.900 ;
        RECT 127.800 143.100 159.300 144.000 ;
        RECT 133.200 142.200 165.600 143.100 ;
        RECT 137.700 141.300 171.900 142.200 ;
        RECT 142.200 140.400 178.200 141.300 ;
        RECT 147.600 139.500 185.400 140.400 ;
        RECT 153.000 138.600 194.400 139.500 ;
        RECT 225.000 138.600 230.400 155.700 ;
        RECT 158.400 137.700 204.300 138.600 ;
        RECT 224.100 137.700 230.400 138.600 ;
        RECT 239.400 137.700 244.800 138.600 ;
        RECT 164.700 136.800 251.100 137.700 ;
        RECT 168.300 135.900 252.000 136.800 ;
        RECT 175.500 135.000 250.200 135.900 ;
        RECT 182.700 134.100 248.400 135.000 ;
        RECT 190.800 133.200 247.500 134.100 ;
        RECT 199.800 132.300 240.300 133.200 ;
        RECT 243.000 132.300 245.700 133.200 ;
        RECT 212.400 131.400 225.900 132.300 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 221.400 294.300 228.600 295.200 ;
        RECT 216.000 293.400 233.100 294.300 ;
        RECT 211.500 292.500 236.700 293.400 ;
        RECT 207.000 291.600 240.300 292.500 ;
        RECT 200.700 290.700 243.000 291.600 ;
        RECT 194.400 289.800 245.700 290.700 ;
        RECT 187.200 288.900 248.400 289.800 ;
        RECT 183.600 288.000 251.100 288.900 ;
        RECT 178.200 287.100 253.800 288.000 ;
        RECT 172.800 286.200 256.500 287.100 ;
        RECT 169.200 285.300 202.500 286.200 ;
        RECT 214.200 285.300 258.300 286.200 ;
        RECT 165.600 284.400 182.700 285.300 ;
        RECT 217.800 284.400 260.100 285.300 ;
        RECT 163.800 283.500 175.500 284.400 ;
        RECT 221.400 283.500 261.900 284.400 ;
        RECT 161.100 282.600 170.100 283.500 ;
        RECT 224.100 282.600 263.700 283.500 ;
        RECT 158.400 281.700 166.500 282.600 ;
        RECT 228.600 281.700 265.500 282.600 ;
        RECT 155.700 280.800 163.800 281.700 ;
        RECT 231.300 280.800 266.400 281.700 ;
        RECT 153.000 279.900 161.100 280.800 ;
        RECT 234.900 279.900 269.100 280.800 ;
        RECT 149.400 279.000 158.400 279.900 ;
        RECT 237.600 279.000 270.000 279.900 ;
        RECT 146.700 278.100 155.700 279.000 ;
        RECT 241.200 278.100 271.800 279.000 ;
        RECT 144.900 277.200 153.000 278.100 ;
        RECT 243.900 277.200 273.600 278.100 ;
        RECT 144.000 276.300 151.200 277.200 ;
        RECT 246.600 276.300 274.500 277.200 ;
        RECT 142.200 275.400 149.400 276.300 ;
        RECT 248.400 275.400 275.400 276.300 ;
        RECT 141.300 274.500 147.600 275.400 ;
        RECT 251.100 274.500 277.200 275.400 ;
        RECT 139.500 273.600 145.800 274.500 ;
        RECT 252.900 273.600 278.100 274.500 ;
        RECT 138.600 272.700 144.000 273.600 ;
        RECT 255.600 272.700 279.900 273.600 ;
        RECT 137.700 271.800 142.200 272.700 ;
        RECT 257.400 271.800 280.800 272.700 ;
        RECT 136.800 270.900 141.300 271.800 ;
        RECT 259.200 270.900 281.700 271.800 ;
        RECT 135.000 270.000 139.500 270.900 ;
        RECT 261.000 270.000 282.600 270.900 ;
        RECT 134.100 269.100 138.600 270.000 ;
        RECT 261.900 269.100 283.500 270.000 ;
        RECT 133.200 268.200 136.800 269.100 ;
        RECT 263.700 268.200 285.300 269.100 ;
        RECT 132.300 267.300 135.900 268.200 ;
        RECT 265.500 267.300 286.200 268.200 ;
        RECT 131.400 266.400 135.000 267.300 ;
        RECT 266.400 266.400 287.100 267.300 ;
        RECT 130.500 265.500 134.100 266.400 ;
        RECT 268.200 265.500 288.000 266.400 ;
        RECT 129.600 264.600 133.200 265.500 ;
        RECT 269.100 264.600 288.900 265.500 ;
        RECT 128.700 263.700 132.300 264.600 ;
        RECT 270.900 263.700 289.800 264.600 ;
        RECT 127.800 262.800 131.400 263.700 ;
        RECT 271.800 262.800 290.700 263.700 ;
        RECT 126.900 261.900 130.500 262.800 ;
        RECT 272.700 261.900 290.700 262.800 ;
        RECT 126.900 261.000 128.700 261.900 ;
        RECT 273.600 261.000 291.600 261.900 ;
        RECT 126.000 260.100 128.700 261.000 ;
        RECT 275.400 260.100 292.500 261.000 ;
        RECT 125.100 259.200 127.800 260.100 ;
        RECT 276.300 259.200 293.400 260.100 ;
        RECT 124.200 258.300 126.900 259.200 ;
        RECT 277.200 258.300 294.300 259.200 ;
        RECT 124.200 257.400 126.000 258.300 ;
        RECT 278.100 257.400 295.200 258.300 ;
        RECT 123.300 256.500 125.100 257.400 ;
        RECT 279.000 256.500 295.200 257.400 ;
        RECT 122.400 255.600 125.100 256.500 ;
        RECT 279.900 255.600 296.100 256.500 ;
        RECT 122.400 254.700 124.200 255.600 ;
        RECT 280.800 254.700 297.000 255.600 ;
        RECT 121.500 253.800 123.300 254.700 ;
        RECT 281.700 253.800 297.000 254.700 ;
        RECT 120.600 252.900 123.300 253.800 ;
        RECT 282.600 252.900 297.900 253.800 ;
        RECT 120.600 252.000 122.400 252.900 ;
        RECT 283.500 252.000 297.900 252.900 ;
        RECT 119.700 250.200 121.500 252.000 ;
        RECT 283.500 251.100 298.800 252.000 ;
        RECT 284.400 250.200 298.800 251.100 ;
        RECT 119.700 249.300 120.600 250.200 ;
        RECT 285.300 249.300 299.700 250.200 ;
        RECT 118.800 248.400 120.600 249.300 ;
        RECT 286.200 248.400 299.700 249.300 ;
        RECT 118.800 247.500 119.700 248.400 ;
        RECT 286.200 247.500 300.600 248.400 ;
        RECT 117.900 246.600 119.700 247.500 ;
        RECT 287.100 246.600 300.600 247.500 ;
        RECT 117.900 244.800 118.800 246.600 ;
        RECT 117.000 243.900 118.800 244.800 ;
        RECT 288.000 245.700 300.600 246.600 ;
        RECT 288.000 243.900 301.500 245.700 ;
        RECT 117.000 242.100 117.900 243.900 ;
        RECT 288.900 242.100 302.400 243.900 ;
        RECT 289.800 241.200 302.400 242.100 ;
        RECT 289.800 239.400 303.300 241.200 ;
        RECT 290.700 236.700 303.300 239.400 ;
        RECT 290.700 235.800 304.200 236.700 ;
        RECT 291.600 232.200 304.200 235.800 ;
        RECT 291.600 231.300 305.100 232.200 ;
        RECT 292.500 225.900 305.100 231.300 ;
        RECT 293.400 216.000 306.000 225.900 ;
        RECT 294.300 214.200 306.000 216.000 ;
        RECT 294.300 186.300 306.900 214.200 ;
        RECT 293.400 175.500 306.000 186.300 ;
        RECT 292.500 174.600 306.000 175.500 ;
        RECT 70.200 172.800 72.000 173.700 ;
        RECT 68.400 171.900 72.000 172.800 ;
        RECT 66.600 171.000 72.900 171.900 ;
        RECT 64.800 170.100 72.900 171.000 ;
        RECT 62.100 169.200 72.900 170.100 ;
        RECT 61.200 168.300 73.800 169.200 ;
        RECT 58.500 167.400 73.800 168.300 ;
        RECT 292.500 167.400 305.100 174.600 ;
        RECT 56.700 166.500 73.800 167.400 ;
        RECT 54.900 165.600 74.700 166.500 ;
        RECT 52.200 164.700 74.700 165.600 ;
        RECT 50.400 163.800 74.700 164.700 ;
        RECT 48.600 162.900 75.600 163.800 ;
        RECT 46.800 162.000 75.600 162.900 ;
        RECT 291.600 162.000 304.200 167.400 ;
        RECT 44.100 161.100 74.700 162.000 ;
        RECT 290.700 161.100 304.200 162.000 ;
        RECT 42.300 160.200 72.900 161.100 ;
        RECT 40.500 159.300 70.200 160.200 ;
        RECT 37.800 158.400 68.400 159.300 ;
        RECT 36.000 157.500 66.600 158.400 ;
        RECT 290.700 157.500 303.300 161.100 ;
        RECT 34.200 156.600 64.800 157.500 ;
        RECT 289.800 156.600 303.300 157.500 ;
        RECT 32.400 155.700 62.100 156.600 ;
        RECT 30.600 154.800 60.300 155.700 ;
        RECT 28.800 153.900 58.500 154.800 ;
        RECT 289.800 153.900 302.400 156.600 ;
        RECT 27.000 153.000 55.800 153.900 ;
        RECT 288.900 153.000 302.400 153.900 ;
        RECT 25.200 152.100 54.900 153.000 ;
        RECT 23.400 151.200 53.100 152.100 ;
        RECT 21.600 150.300 51.300 151.200 ;
        RECT 288.900 150.300 301.500 153.000 ;
        RECT 19.800 149.400 48.600 150.300 ;
        RECT 18.000 148.500 46.800 149.400 ;
        RECT 288.000 148.500 300.600 150.300 ;
        RECT 16.200 147.600 45.000 148.500 ;
        RECT 287.100 147.600 300.600 148.500 ;
        RECT 15.300 146.700 43.200 147.600 ;
        RECT 287.100 146.700 299.700 147.600 ;
        RECT 13.500 145.800 40.500 146.700 ;
        RECT 11.700 144.900 38.700 145.800 ;
        RECT 286.200 144.900 299.700 146.700 ;
        RECT 10.800 144.000 36.900 144.900 ;
        RECT 285.300 144.000 298.800 144.900 ;
        RECT 9.900 143.100 35.100 144.000 ;
        RECT 283.500 143.100 298.800 144.000 ;
        RECT 8.100 142.200 33.300 143.100 ;
        RECT 281.700 142.200 298.800 143.100 ;
        RECT 8.100 141.300 31.500 142.200 ;
        RECT 280.800 141.300 297.900 142.200 ;
        RECT 7.200 140.400 29.700 141.300 ;
        RECT 279.000 140.400 297.900 141.300 ;
        RECT 6.300 139.500 27.900 140.400 ;
        RECT 276.300 139.500 297.000 140.400 ;
        RECT 5.400 138.600 26.100 139.500 ;
        RECT 274.500 138.600 296.100 139.500 ;
        RECT 5.400 137.700 24.300 138.600 ;
        RECT 271.800 137.700 296.100 138.600 ;
        RECT 4.500 136.800 22.500 137.700 ;
        RECT 269.100 136.800 295.200 137.700 ;
        RECT 4.500 135.900 21.600 136.800 ;
        RECT 266.400 135.900 294.300 136.800 ;
        RECT 4.500 135.000 19.800 135.900 ;
        RECT 261.900 135.000 293.400 135.900 ;
        RECT 3.600 134.100 18.900 135.000 ;
        RECT 259.200 134.100 292.500 135.000 ;
        RECT 3.600 132.300 17.100 134.100 ;
        RECT 255.600 133.200 291.600 134.100 ;
        RECT 253.800 132.300 289.800 133.200 ;
        RECT 3.600 128.700 16.200 132.300 ;
        RECT 252.000 131.400 288.900 132.300 ;
        RECT 250.200 130.500 287.100 131.400 ;
        RECT 249.300 129.600 285.300 130.500 ;
        RECT 247.500 128.700 283.500 129.600 ;
        RECT 3.600 126.900 17.100 128.700 ;
        RECT 245.700 127.800 281.700 128.700 ;
        RECT 243.900 126.900 279.000 127.800 ;
        RECT 3.600 126.000 18.900 126.900 ;
        RECT 243.000 126.000 276.300 126.900 ;
        RECT 4.500 125.100 19.800 126.000 ;
        RECT 242.100 125.100 273.600 126.000 ;
        RECT 4.500 124.200 21.600 125.100 ;
        RECT 241.200 124.200 270.000 125.100 ;
        RECT 4.500 123.300 23.400 124.200 ;
        RECT 240.300 123.300 266.400 124.200 ;
        RECT 5.400 122.400 26.100 123.300 ;
        RECT 238.500 122.400 261.900 123.300 ;
        RECT 6.300 121.500 28.800 122.400 ;
        RECT 237.600 121.500 258.300 122.400 ;
        RECT 6.300 120.600 32.400 121.500 ;
        RECT 236.700 120.600 256.500 121.500 ;
        RECT 7.200 119.700 34.200 120.600 ;
        RECT 235.800 119.700 255.600 120.600 ;
        RECT 7.200 118.800 36.900 119.700 ;
        RECT 234.900 118.800 254.700 119.700 ;
        RECT 8.100 117.900 40.500 118.800 ;
        RECT 233.100 117.900 253.800 118.800 ;
        RECT 9.900 117.000 43.200 117.900 ;
        RECT 232.200 117.000 252.000 117.900 ;
        RECT 10.800 116.100 46.800 117.000 ;
        RECT 230.400 116.100 251.100 117.000 ;
        RECT 11.700 115.200 49.500 116.100 ;
        RECT 229.500 115.200 250.200 116.100 ;
        RECT 13.500 114.300 53.100 115.200 ;
        RECT 227.700 114.300 248.400 115.200 ;
        RECT 14.400 113.400 55.800 114.300 ;
        RECT 226.800 113.400 247.500 114.300 ;
        RECT 16.200 112.500 59.400 113.400 ;
        RECT 225.000 112.500 246.600 113.400 ;
        RECT 18.900 111.600 63.000 112.500 ;
        RECT 223.200 111.600 245.700 112.500 ;
        RECT 21.600 110.700 65.700 111.600 ;
        RECT 221.400 110.700 244.800 111.600 ;
        RECT 24.300 109.800 69.300 110.700 ;
        RECT 219.600 109.800 243.000 110.700 ;
        RECT 27.000 108.900 72.000 109.800 ;
        RECT 216.900 108.900 242.100 109.800 ;
        RECT 29.700 108.000 75.600 108.900 ;
        RECT 215.100 108.000 241.200 108.900 ;
        RECT 32.400 107.100 79.200 108.000 ;
        RECT 213.300 107.100 239.400 108.000 ;
        RECT 36.000 106.200 82.800 107.100 ;
        RECT 210.600 106.200 238.500 107.100 ;
        RECT 38.700 105.300 86.400 106.200 ;
        RECT 208.800 105.300 236.700 106.200 ;
        RECT 41.400 104.400 90.000 105.300 ;
        RECT 206.100 104.400 235.800 105.300 ;
        RECT 44.100 103.500 92.700 104.400 ;
        RECT 204.300 103.500 234.000 104.400 ;
        RECT 46.800 102.600 96.300 103.500 ;
        RECT 201.600 102.600 232.200 103.500 ;
        RECT 50.400 101.700 100.800 102.600 ;
        RECT 198.900 101.700 231.300 102.600 ;
        RECT 54.000 100.800 104.400 101.700 ;
        RECT 195.300 100.800 229.500 101.700 ;
        RECT 56.700 99.900 108.900 100.800 ;
        RECT 192.600 99.900 227.700 100.800 ;
        RECT 60.300 99.000 113.400 99.900 ;
        RECT 189.000 99.000 225.900 99.900 ;
        RECT 63.900 98.100 118.800 99.000 ;
        RECT 185.400 98.100 224.100 99.000 ;
        RECT 67.500 97.200 124.200 98.100 ;
        RECT 180.000 97.200 222.300 98.100 ;
        RECT 71.100 96.300 129.600 97.200 ;
        RECT 175.500 96.300 220.500 97.200 ;
        RECT 73.800 95.400 135.900 96.300 ;
        RECT 168.300 95.400 217.800 96.300 ;
        RECT 78.300 94.500 145.800 95.400 ;
        RECT 156.600 94.500 215.100 95.400 ;
        RECT 81.900 93.600 213.300 94.500 ;
        RECT 85.500 92.700 210.600 93.600 ;
        RECT 89.100 91.800 207.900 92.700 ;
        RECT 92.700 90.900 205.200 91.800 ;
        RECT 97.200 90.000 202.500 90.900 ;
        RECT 100.800 89.100 199.800 90.000 ;
        RECT 105.300 88.200 196.200 89.100 ;
        RECT 108.000 87.300 193.500 88.200 ;
        RECT 112.500 86.400 189.900 87.300 ;
        RECT 117.900 85.500 186.300 86.400 ;
        RECT 122.400 84.600 180.900 85.500 ;
        RECT 128.700 83.700 175.500 84.600 ;
        RECT 135.900 82.800 168.300 83.700 ;
        RECT 145.800 81.900 158.400 82.800 ;
    END
  END vdd
  OBS
      LAYER Metal2 ;
        RECT 0.000 0.000 310.500 310.500 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 310.500 310.500 ;
      LAYER Metal4 ;
        RECT 195.300 304.200 198.900 305.100 ;
        RECT 188.100 303.300 206.100 304.200 ;
        RECT 184.500 302.400 208.800 303.300 ;
        RECT 182.700 301.500 210.600 302.400 ;
        RECT 181.800 300.600 212.400 301.500 ;
        RECT 180.000 299.700 213.300 300.600 ;
        RECT 179.100 298.800 214.200 299.700 ;
        RECT 178.200 297.900 215.100 298.800 ;
        RECT 179.100 297.000 214.200 297.900 ;
        RECT 183.600 296.100 209.700 297.000 ;
        RECT 188.100 295.200 205.200 296.100 ;
        RECT 245.700 273.600 248.400 274.500 ;
        RECT 245.700 272.700 250.200 273.600 ;
        RECT 245.700 271.800 252.000 272.700 ;
        RECT 246.600 270.900 251.100 271.800 ;
        RECT 248.400 270.000 249.300 270.900 ;
        RECT 255.600 269.100 256.500 270.000 ;
        RECT 253.800 268.200 258.300 269.100 ;
        RECT 253.800 267.300 259.200 268.200 ;
        RECT 252.900 265.500 260.100 267.300 ;
        RECT 253.800 264.600 260.100 265.500 ;
        RECT 253.800 263.700 259.200 264.600 ;
        RECT 254.700 262.800 258.300 263.700 ;
        RECT 246.600 261.000 251.100 261.900 ;
        RECT 262.800 261.000 266.400 261.900 ;
        RECT 246.600 260.100 252.000 261.000 ;
        RECT 261.000 260.100 267.300 261.000 ;
        RECT 246.600 257.400 252.900 260.100 ;
        RECT 261.000 257.400 268.200 260.100 ;
        RECT 246.600 256.500 252.000 257.400 ;
        RECT 261.000 256.500 267.300 257.400 ;
        RECT 247.500 255.600 251.100 256.500 ;
        RECT 261.900 255.600 266.400 256.500 ;
        RECT 248.400 254.700 249.300 255.600 ;
        RECT 263.700 254.700 264.600 255.600 ;
        RECT 255.600 253.800 257.400 254.700 ;
        RECT 270.900 253.800 273.600 254.700 ;
        RECT 253.800 252.900 259.200 253.800 ;
        RECT 270.000 252.900 274.500 253.800 ;
        RECT 253.800 252.000 260.100 252.900 ;
        RECT 252.900 250.200 260.100 252.000 ;
        RECT 253.800 249.300 260.100 250.200 ;
        RECT 253.800 248.400 259.200 249.300 ;
        RECT 269.100 248.400 275.400 252.900 ;
        RECT 254.700 247.500 259.200 248.400 ;
        RECT 270.000 247.500 274.500 248.400 ;
        RECT 262.800 245.700 265.500 246.600 ;
        RECT 278.100 245.700 281.700 246.600 ;
        RECT 261.900 244.800 267.300 245.700 ;
        RECT 277.200 244.800 282.600 245.700 ;
        RECT 261.000 242.100 268.200 244.800 ;
        RECT 276.300 243.900 282.600 244.800 ;
        RECT 276.300 242.100 283.500 243.900 ;
        RECT 261.000 241.200 267.300 242.100 ;
        RECT 276.300 241.200 282.600 242.100 ;
        RECT 261.900 240.300 266.400 241.200 ;
        RECT 277.200 240.300 281.700 241.200 ;
        RECT 262.800 239.400 265.500 240.300 ;
        RECT 279.000 239.400 280.800 240.300 ;
        RECT 255.600 238.500 257.400 239.400 ;
        RECT 270.900 238.500 272.700 239.400 ;
        RECT 254.700 237.600 259.200 238.500 ;
        RECT 270.000 237.600 274.500 238.500 ;
        RECT 282.600 237.600 286.200 238.500 ;
        RECT 253.800 236.700 260.100 237.600 ;
        RECT 252.900 234.900 260.100 236.700 ;
        RECT 253.800 234.000 260.100 234.900 ;
        RECT 269.100 234.000 275.400 237.600 ;
        RECT 281.700 234.000 287.100 237.600 ;
        RECT 253.800 233.100 259.200 234.000 ;
        RECT 269.100 233.100 274.500 234.000 ;
        RECT 278.100 233.100 288.000 234.000 ;
        RECT 254.700 232.200 259.200 233.100 ;
        RECT 270.000 232.200 274.500 233.100 ;
        RECT 277.200 231.300 288.000 233.100 ;
        RECT 262.800 230.400 265.500 231.300 ;
        RECT 276.300 230.400 287.100 231.300 ;
        RECT 261.900 229.500 267.300 230.400 ;
        RECT 276.300 229.500 286.200 230.400 ;
        RECT 261.000 228.600 267.300 229.500 ;
        RECT 261.000 226.800 268.200 228.600 ;
        RECT 275.400 226.800 285.300 229.500 ;
        RECT 102.600 225.900 110.700 226.800 ;
        RECT 261.000 225.900 267.300 226.800 ;
        RECT 102.600 225.000 117.900 225.900 ;
        RECT 137.700 225.000 141.300 225.900 ;
        RECT 261.900 225.000 267.300 225.900 ;
        RECT 274.500 225.900 286.200 226.800 ;
        RECT 274.500 225.000 288.900 225.900 ;
        RECT 102.600 224.100 118.800 225.000 ;
        RECT 133.200 224.100 145.800 225.000 ;
        RECT 262.800 224.100 265.500 225.000 ;
        RECT 273.600 224.100 288.900 225.000 ;
        RECT 101.700 216.900 119.700 224.100 ;
        RECT 130.500 223.200 147.600 224.100 ;
        RECT 271.800 223.200 289.800 224.100 ;
        RECT 129.600 222.300 149.400 223.200 ;
        RECT 254.700 222.300 259.200 223.200 ;
        RECT 270.000 222.300 289.800 223.200 ;
        RECT 128.700 221.400 150.300 222.300 ;
        RECT 159.300 221.400 171.900 222.300 ;
        RECT 187.200 221.400 195.300 222.300 ;
        RECT 253.800 221.400 260.100 222.300 ;
        RECT 127.800 220.500 152.100 221.400 ;
        RECT 126.900 219.600 152.100 220.500 ;
        RECT 126.900 218.700 153.000 219.600 ;
        RECT 100.800 210.600 120.600 216.900 ;
        RECT 126.000 215.100 153.900 218.700 ;
        RECT 126.000 214.200 138.600 215.100 ;
        RECT 140.400 214.200 154.800 215.100 ;
        RECT 99.900 208.800 120.600 210.600 ;
        RECT 125.100 208.800 137.700 214.200 ;
        RECT 99.900 205.200 121.500 208.800 ;
        RECT 125.100 207.000 138.600 208.800 ;
        RECT 141.300 207.000 154.800 214.200 ;
        RECT 125.100 206.100 139.500 207.000 ;
        RECT 145.800 206.100 154.800 207.000 ;
        RECT 99.900 203.400 109.800 205.200 ;
        RECT 110.700 204.300 121.500 205.200 ;
        RECT 99.000 197.100 109.800 203.400 ;
        RECT 98.100 196.200 109.800 197.100 ;
        RECT 111.600 200.700 121.500 204.300 ;
        RECT 126.000 205.200 140.400 206.100 ;
        RECT 126.000 204.300 141.300 205.200 ;
        RECT 126.000 203.400 142.200 204.300 ;
        RECT 126.000 202.500 144.000 203.400 ;
        RECT 126.900 201.600 144.900 202.500 ;
        RECT 126.900 200.700 145.800 201.600 ;
        RECT 98.100 193.500 108.900 196.200 ;
        RECT 111.600 193.500 122.400 200.700 ;
        RECT 127.800 199.800 146.700 200.700 ;
        RECT 127.800 198.900 147.600 199.800 ;
        RECT 128.700 198.000 149.400 198.900 ;
        RECT 129.600 197.100 150.300 198.000 ;
        RECT 130.500 196.200 151.200 197.100 ;
        RECT 131.400 195.300 152.100 196.200 ;
        RECT 132.300 194.400 153.000 195.300 ;
        RECT 134.100 193.500 153.000 194.400 ;
        RECT 98.100 192.600 109.800 193.500 ;
        RECT 111.600 192.600 123.300 193.500 ;
        RECT 135.000 192.600 153.900 193.500 ;
        RECT 98.100 190.800 123.300 192.600 ;
        RECT 135.900 191.700 153.900 192.600 ;
        RECT 136.800 190.800 154.800 191.700 ;
        RECT 97.200 187.200 123.300 190.800 ;
        RECT 137.700 189.900 154.800 190.800 ;
        RECT 126.000 189.000 135.000 189.900 ;
        RECT 138.600 189.000 154.800 189.900 ;
        RECT 97.200 183.600 124.200 187.200 ;
        RECT 96.300 182.700 124.200 183.600 ;
        RECT 96.300 181.800 109.800 182.700 ;
        RECT 111.600 181.800 124.200 182.700 ;
        RECT 96.300 177.300 108.900 181.800 ;
        RECT 112.500 180.900 124.200 181.800 ;
        RECT 126.000 186.300 137.700 189.000 ;
        RECT 140.400 188.100 154.800 189.000 ;
        RECT 140.400 187.200 155.700 188.100 ;
        RECT 112.500 180.000 125.100 180.900 ;
        RECT 126.000 180.000 138.600 186.300 ;
        RECT 141.300 185.400 155.700 187.200 ;
        RECT 97.200 176.400 108.900 177.300 ;
        RECT 100.800 175.500 108.900 176.400 ;
        RECT 105.300 174.600 108.900 175.500 ;
        RECT 113.400 175.500 125.100 180.000 ;
        RECT 126.900 178.200 138.600 180.000 ;
        RECT 142.200 179.100 155.700 185.400 ;
        RECT 159.300 186.300 172.800 221.400 ;
        RECT 184.500 220.500 198.000 221.400 ;
        RECT 182.700 219.600 199.800 220.500 ;
        RECT 252.900 219.600 260.100 221.400 ;
        RECT 181.800 218.700 201.600 219.600 ;
        RECT 253.800 218.700 260.100 219.600 ;
        RECT 269.100 218.700 277.200 222.300 ;
        RECT 180.000 217.800 202.500 218.700 ;
        RECT 253.800 217.800 259.200 218.700 ;
        RECT 270.000 217.800 277.200 218.700 ;
        RECT 281.700 217.800 289.800 222.300 ;
        RECT 179.100 216.000 203.400 217.800 ;
        RECT 254.700 216.900 258.300 217.800 ;
        RECT 256.500 216.000 257.400 216.900 ;
        RECT 178.200 215.100 204.300 216.000 ;
        RECT 262.800 215.100 265.500 216.000 ;
        RECT 270.900 215.100 289.800 217.800 ;
        RECT 178.200 214.200 205.200 215.100 ;
        RECT 250.200 214.200 252.000 215.100 ;
        RECT 261.900 214.200 266.400 215.100 ;
        RECT 271.800 214.200 288.900 215.100 ;
        RECT 177.300 212.400 205.200 214.200 ;
        RECT 249.300 213.300 252.000 214.200 ;
        RECT 261.000 213.300 267.300 214.200 ;
        RECT 273.600 213.300 285.300 214.200 ;
        RECT 177.300 211.500 206.100 212.400 ;
        RECT 176.400 210.600 190.800 211.500 ;
        RECT 192.600 210.600 206.100 211.500 ;
        RECT 176.400 186.300 189.900 210.600 ;
        RECT 193.500 196.200 206.100 210.600 ;
        RECT 249.300 211.500 252.900 213.300 ;
        RECT 249.300 209.700 252.000 211.500 ;
        RECT 261.000 210.600 268.200 213.300 ;
        RECT 274.500 211.500 285.300 213.300 ;
        RECT 273.600 210.600 285.300 211.500 ;
        RECT 261.900 209.700 267.300 210.600 ;
        RECT 270.900 209.700 289.800 210.600 ;
        RECT 249.300 208.800 251.100 209.700 ;
        RECT 262.800 208.800 265.500 209.700 ;
        RECT 270.000 208.800 289.800 209.700 ;
        RECT 254.700 207.000 259.200 207.900 ;
        RECT 253.800 206.100 259.200 207.000 ;
        RECT 269.100 207.000 290.700 208.800 ;
        RECT 269.100 206.100 277.200 207.000 ;
        RECT 253.800 205.200 260.100 206.100 ;
        RECT 252.900 204.300 260.100 205.200 ;
        RECT 253.800 203.400 260.100 204.300 ;
        RECT 253.800 202.500 259.200 203.400 ;
        RECT 268.200 202.500 277.200 206.100 ;
        RECT 281.700 202.500 290.700 207.000 ;
        RECT 254.700 201.600 259.200 202.500 ;
        RECT 267.300 200.700 290.700 202.500 ;
        RECT 248.400 199.800 249.300 200.700 ;
        RECT 266.400 199.800 290.700 200.700 ;
        RECT 246.600 198.900 251.100 199.800 ;
        RECT 261.900 198.900 289.800 199.800 ;
        RECT 246.600 198.000 252.000 198.900 ;
        RECT 198.900 195.300 206.100 196.200 ;
        RECT 245.700 196.200 252.900 198.000 ;
        RECT 245.700 194.400 252.000 196.200 ;
        RECT 261.000 195.300 270.000 198.900 ;
        RECT 261.900 194.400 270.000 195.300 ;
        RECT 274.500 195.300 285.300 198.900 ;
        RECT 274.500 194.400 288.900 195.300 ;
        RECT 246.600 193.500 251.100 194.400 ;
        RECT 262.800 193.500 289.800 194.400 ;
        RECT 264.600 192.600 290.700 193.500 ;
        RECT 254.700 191.700 258.300 192.600 ;
        RECT 265.500 191.700 290.700 192.600 ;
        RECT 253.800 190.800 259.200 191.700 ;
        RECT 253.800 189.900 260.100 190.800 ;
        RECT 252.900 188.100 260.100 189.900 ;
        RECT 266.400 188.100 277.200 191.700 ;
        RECT 193.500 187.200 197.100 188.100 ;
        RECT 253.800 187.200 260.100 188.100 ;
        RECT 265.500 187.200 277.200 188.100 ;
        RECT 281.700 187.200 290.700 191.700 ;
        RECT 193.500 186.300 206.100 187.200 ;
        RECT 254.700 186.300 259.200 187.200 ;
        RECT 264.600 186.300 289.800 187.200 ;
        RECT 159.300 182.700 171.900 186.300 ;
        RECT 141.300 178.200 155.700 179.100 ;
        RECT 126.900 177.300 155.700 178.200 ;
        RECT 127.800 175.500 155.700 177.300 ;
        RECT 113.400 173.700 126.000 175.500 ;
        RECT 127.800 174.600 154.800 175.500 ;
        RECT 128.700 173.700 154.800 174.600 ;
        RECT 114.300 172.800 126.000 173.700 ;
        RECT 129.600 172.800 154.800 173.700 ;
        RECT 118.800 171.900 126.000 172.800 ;
        RECT 130.500 171.900 153.900 172.800 ;
        RECT 123.300 171.000 126.000 171.900 ;
        RECT 132.300 171.000 153.900 171.900 ;
        RECT 133.200 170.100 153.000 171.000 ;
        RECT 158.400 170.100 171.900 182.700 ;
        RECT 176.400 175.500 189.000 186.300 ;
        RECT 192.600 178.200 206.100 186.300 ;
        RECT 263.700 185.400 289.800 186.300 ;
        RECT 247.500 184.500 250.200 185.400 ;
        RECT 262.800 184.500 289.800 185.400 ;
        RECT 246.600 183.600 251.100 184.500 ;
        RECT 261.900 183.600 288.900 184.500 ;
        RECT 245.700 182.700 252.000 183.600 ;
        RECT 245.700 180.900 252.900 182.700 ;
        RECT 245.700 179.100 252.000 180.900 ;
        RECT 261.000 179.100 270.000 183.600 ;
        RECT 274.500 182.700 286.200 183.600 ;
        RECT 274.500 180.000 285.300 182.700 ;
        RECT 274.500 179.100 286.200 180.000 ;
        RECT 246.600 178.200 251.100 179.100 ;
        RECT 261.000 178.200 288.900 179.100 ;
        RECT 176.400 174.600 189.900 175.500 ;
        RECT 192.600 174.600 205.200 178.200 ;
        RECT 239.400 176.400 243.000 177.300 ;
        RECT 255.600 176.400 257.400 177.300 ;
        RECT 260.100 176.400 288.900 178.200 ;
        RECT 239.400 175.500 243.900 176.400 ;
        RECT 176.400 173.700 190.800 174.600 ;
        RECT 191.700 173.700 205.200 174.600 ;
        RECT 177.300 172.800 205.200 173.700 ;
        RECT 177.300 171.000 204.300 172.800 ;
        RECT 238.500 171.900 244.800 175.500 ;
        RECT 253.800 174.600 261.900 176.400 ;
        RECT 252.900 172.800 261.900 174.600 ;
        RECT 253.800 171.900 261.900 172.800 ;
        RECT 266.400 171.900 277.200 176.400 ;
        RECT 281.700 173.700 289.800 176.400 ;
        RECT 281.700 171.900 288.900 173.700 ;
        RECT 238.500 171.000 243.900 171.900 ;
        RECT 254.700 171.000 288.900 171.900 ;
        RECT 178.200 170.100 203.400 171.000 ;
        RECT 240.300 170.100 242.100 171.000 ;
        RECT 135.000 169.200 151.200 170.100 ;
        RECT 135.900 168.300 150.300 169.200 ;
        RECT 139.500 167.400 147.600 168.300 ;
        RECT 159.300 166.500 171.900 170.100 ;
        RECT 179.100 169.200 203.400 170.100 ;
        RECT 247.500 169.200 250.200 170.100 ;
        RECT 255.600 169.200 288.000 171.000 ;
        RECT 179.100 168.300 202.500 169.200 ;
        RECT 246.600 168.300 251.100 169.200 ;
        RECT 256.500 168.300 287.100 169.200 ;
        RECT 180.000 167.400 201.600 168.300 ;
        RECT 245.700 167.400 252.000 168.300 ;
        RECT 257.400 167.400 270.000 168.300 ;
        RECT 180.900 166.500 200.700 167.400 ;
        RECT 170.100 165.600 171.900 166.500 ;
        RECT 182.700 165.600 199.800 166.500 ;
        RECT 245.700 165.600 252.900 167.400 ;
        RECT 184.500 164.700 198.000 165.600 ;
        RECT 186.300 163.800 195.300 164.700 ;
        RECT 245.700 163.800 252.000 165.600 ;
        RECT 258.300 163.800 270.000 167.400 ;
        RECT 274.500 167.400 286.200 168.300 ;
        RECT 274.500 163.800 285.300 167.400 ;
        RECT 246.600 162.900 251.100 163.800 ;
        RECT 253.800 162.900 286.200 163.800 ;
        RECT 252.900 162.000 286.200 162.900 ;
        RECT 239.400 161.100 243.000 162.000 ;
        RECT 252.000 161.100 286.200 162.000 ;
        RECT 238.500 160.200 243.900 161.100 ;
        RECT 252.000 160.200 261.900 161.100 ;
        RECT 237.600 157.500 244.800 160.200 ;
        RECT 238.500 156.600 244.800 157.500 ;
        RECT 251.100 156.600 261.900 160.200 ;
        RECT 238.500 155.700 243.900 156.600 ;
        RECT 250.200 155.700 261.900 156.600 ;
        RECT 263.700 155.700 265.500 156.600 ;
        RECT 266.400 155.700 277.200 161.100 ;
        RECT 281.700 158.400 287.100 161.100 ;
        RECT 281.700 156.600 286.200 158.400 ;
        RECT 279.000 155.700 280.800 156.600 ;
        RECT 281.700 155.700 283.500 156.600 ;
        RECT 240.300 154.800 242.100 155.700 ;
        RECT 249.300 154.800 283.500 155.700 ;
        RECT 248.400 153.900 282.600 154.800 ;
        RECT 246.600 153.000 282.600 153.900 ;
        RECT 246.600 152.100 254.700 153.000 ;
        RECT 245.700 148.500 254.700 152.100 ;
        RECT 259.200 148.500 270.000 153.000 ;
        RECT 274.500 148.500 282.600 153.000 ;
        RECT 246.600 147.600 281.700 148.500 ;
        RECT 247.500 146.700 279.900 147.600 ;
        RECT 240.300 145.800 243.000 146.700 ;
        RECT 248.400 145.800 275.400 146.700 ;
        RECT 238.500 144.900 243.900 145.800 ;
        RECT 249.300 144.900 275.400 145.800 ;
        RECT 237.600 143.100 244.800 144.900 ;
        RECT 251.100 143.100 261.900 144.900 ;
        RECT 265.500 144.000 275.400 144.900 ;
        RECT 237.600 142.200 243.900 143.100 ;
        RECT 252.000 142.200 261.900 143.100 ;
        RECT 266.400 143.100 275.400 144.000 ;
        RECT 266.400 142.200 274.500 143.100 ;
        RECT 252.900 141.300 261.900 142.200 ;
        RECT 269.100 141.300 273.600 142.200 ;
        RECT 253.800 140.400 260.100 141.300 ;
        RECT 270.000 140.400 271.800 141.300 ;
        RECT 254.700 139.500 258.300 140.400 ;
        RECT 140.400 132.300 157.500 133.200 ;
        RECT 133.200 131.400 164.700 132.300 ;
        RECT 128.700 130.500 170.100 131.400 ;
        RECT 125.100 129.600 173.700 130.500 ;
        RECT 120.600 128.700 177.300 129.600 ;
        RECT 117.900 127.800 180.000 128.700 ;
        RECT 115.200 126.900 181.800 127.800 ;
        RECT 113.400 126.000 184.500 126.900 ;
        RECT 111.600 125.100 186.300 126.000 ;
        RECT 109.800 124.200 187.200 125.100 ;
        RECT 108.900 123.300 189.000 124.200 ;
        RECT 107.100 122.400 189.900 123.300 ;
        RECT 107.100 121.500 190.800 122.400 ;
        RECT 106.200 120.600 191.700 121.500 ;
        RECT 105.300 119.700 191.700 120.600 ;
        RECT 105.300 116.100 192.600 119.700 ;
        RECT 105.300 114.300 191.700 116.100 ;
        RECT 106.200 113.400 190.800 114.300 ;
        RECT 107.100 112.500 190.800 113.400 ;
        RECT 108.000 111.600 189.900 112.500 ;
        RECT 108.900 110.700 188.100 111.600 ;
        RECT 110.700 109.800 187.200 110.700 ;
        RECT 112.500 108.900 185.400 109.800 ;
        RECT 114.300 108.000 183.600 108.900 ;
        RECT 117.000 107.100 180.900 108.000 ;
        RECT 118.800 106.200 179.100 107.100 ;
        RECT 121.500 105.300 176.400 106.200 ;
        RECT 125.100 104.400 172.800 105.300 ;
        RECT 128.700 103.500 169.200 104.400 ;
        RECT 133.200 102.600 164.700 103.500 ;
        RECT 140.400 101.700 157.500 102.600 ;
        RECT 65.700 71.100 70.200 72.900 ;
        RECT 64.800 70.200 70.200 71.100 ;
        RECT 90.000 70.200 91.800 71.100 ;
        RECT 64.800 69.300 71.100 70.200 ;
        RECT 64.800 68.400 67.500 69.300 ;
        RECT 63.900 67.500 67.500 68.400 ;
        RECT 68.400 67.500 71.100 69.300 ;
        RECT 89.100 68.400 91.800 70.200 ;
        RECT 76.500 67.500 79.200 68.400 ;
        RECT 81.000 67.500 84.600 68.400 ;
        RECT 63.900 65.700 66.600 67.500 ;
        RECT 63.000 64.800 66.600 65.700 ;
        RECT 69.300 65.700 72.000 67.500 ;
        RECT 76.500 66.600 85.500 67.500 ;
        RECT 88.200 66.600 94.500 68.400 ;
        RECT 99.000 67.500 102.600 68.400 ;
        RECT 108.900 67.500 111.600 68.400 ;
        RECT 112.500 67.500 117.000 68.400 ;
        RECT 97.200 66.600 104.400 67.500 ;
        RECT 108.900 66.600 117.900 67.500 ;
        RECT 69.300 64.800 72.900 65.700 ;
        RECT 63.000 63.900 65.700 64.800 ;
        RECT 70.200 63.900 72.900 64.800 ;
        RECT 63.000 63.000 72.900 63.900 ;
        RECT 76.500 64.800 80.100 66.600 ;
        RECT 82.800 65.700 86.400 66.600 ;
        RECT 62.100 61.200 73.800 63.000 ;
        RECT 62.100 60.300 64.800 61.200 ;
        RECT 61.200 59.400 64.800 60.300 ;
        RECT 71.100 60.300 73.800 61.200 ;
        RECT 71.100 59.400 74.700 60.300 ;
        RECT 61.200 57.600 63.900 59.400 ;
        RECT 72.000 57.600 74.700 59.400 ;
        RECT 76.500 57.600 79.200 64.800 ;
        RECT 83.700 57.600 86.400 65.700 ;
        RECT 89.100 60.300 91.800 66.600 ;
        RECT 96.300 65.700 99.900 66.600 ;
        RECT 102.600 65.700 105.300 66.600 ;
        RECT 108.900 65.700 112.500 66.600 ;
        RECT 95.400 64.800 99.000 65.700 ;
        RECT 102.600 64.800 106.200 65.700 ;
        RECT 95.400 61.200 98.100 64.800 ;
        RECT 103.500 61.200 106.200 64.800 ;
        RECT 95.400 60.300 99.000 61.200 ;
        RECT 102.600 60.300 106.200 61.200 ;
        RECT 89.100 59.400 92.700 60.300 ;
        RECT 96.300 59.400 99.900 60.300 ;
        RECT 102.600 59.400 105.300 60.300 ;
        RECT 90.000 58.500 94.500 59.400 ;
        RECT 97.200 58.500 104.400 59.400 ;
        RECT 90.900 57.600 94.500 58.500 ;
        RECT 99.000 57.600 102.600 58.500 ;
        RECT 108.900 57.600 111.600 65.700 ;
        RECT 115.200 57.600 117.900 66.600 ;
        RECT 126.000 64.800 128.700 68.400 ;
        RECT 132.300 67.500 135.000 68.400 ;
        RECT 131.400 65.700 135.000 67.500 ;
        RECT 138.600 66.600 141.300 68.400 ;
        RECT 145.800 67.500 149.400 68.400 ;
        RECT 144.000 66.600 151.200 67.500 ;
        RECT 126.900 62.100 129.600 64.800 ;
        RECT 131.400 63.900 135.900 65.700 ;
        RECT 137.700 63.900 140.400 66.600 ;
        RECT 143.100 65.700 146.700 66.600 ;
        RECT 149.400 65.700 152.100 66.600 ;
        RECT 142.200 64.800 145.800 65.700 ;
        RECT 149.400 64.800 153.000 65.700 ;
        RECT 130.500 62.100 133.200 63.900 ;
        RECT 134.100 62.100 135.900 63.900 ;
        RECT 136.800 62.100 139.500 63.900 ;
        RECT 127.800 59.400 132.300 62.100 ;
        RECT 134.100 61.200 139.500 62.100 ;
        RECT 142.200 61.200 144.900 64.800 ;
        RECT 150.300 61.200 153.000 64.800 ;
        RECT 134.100 60.300 138.600 61.200 ;
        RECT 142.200 60.300 145.800 61.200 ;
        RECT 149.400 60.300 153.000 61.200 ;
        RECT 128.700 58.500 132.300 59.400 ;
        RECT 135.000 58.500 138.600 60.300 ;
        RECT 143.100 59.400 146.700 60.300 ;
        RECT 149.400 59.400 152.100 60.300 ;
        RECT 155.700 59.400 158.400 68.400 ;
        RECT 162.000 60.300 164.700 68.400 ;
        RECT 161.100 59.400 164.700 60.300 ;
        RECT 144.000 58.500 151.200 59.400 ;
        RECT 155.700 58.500 164.700 59.400 ;
        RECT 128.700 57.600 131.400 58.500 ;
        RECT 135.000 57.600 137.700 58.500 ;
        RECT 145.800 57.600 149.400 58.500 ;
        RECT 157.500 57.600 161.100 58.500 ;
        RECT 162.900 57.600 164.700 58.500 ;
        RECT 168.300 57.600 171.000 72.900 ;
        RECT 175.500 67.500 179.100 68.400 ;
        RECT 180.900 67.500 183.600 72.900 ;
        RECT 174.600 66.600 183.600 67.500 ;
        RECT 173.700 65.700 177.300 66.600 ;
        RECT 179.100 65.700 183.600 66.600 ;
        RECT 173.700 64.800 176.400 65.700 ;
        RECT 180.000 64.800 183.600 65.700 ;
        RECT 172.800 63.900 176.400 64.800 ;
        RECT 172.800 62.100 175.500 63.900 ;
        RECT 172.800 61.200 176.400 62.100 ;
        RECT 180.900 61.200 183.600 64.800 ;
        RECT 173.700 60.300 176.400 61.200 ;
        RECT 180.000 60.300 183.600 61.200 ;
        RECT 173.700 59.400 177.300 60.300 ;
        RECT 179.100 59.400 183.600 60.300 ;
        RECT 174.600 58.500 183.600 59.400 ;
        RECT 175.500 57.600 179.100 58.500 ;
        RECT 180.900 57.600 183.600 58.500 ;
        RECT 191.700 57.600 194.400 72.900 ;
        RECT 197.100 70.200 199.800 72.900 ;
        RECT 197.100 57.600 199.800 68.400 ;
        RECT 203.400 64.800 206.100 72.900 ;
        RECT 232.200 68.400 234.900 71.100 ;
        RECT 208.800 67.500 212.400 68.400 ;
        RECT 216.900 67.500 220.500 68.400 ;
        RECT 207.900 66.600 211.500 67.500 ;
        RECT 215.100 66.600 222.300 67.500 ;
        RECT 230.400 66.600 236.700 68.400 ;
        RECT 241.200 67.500 245.700 68.400 ;
        RECT 239.400 66.600 247.500 67.500 ;
        RECT 207.900 65.700 210.600 66.600 ;
        RECT 214.200 65.700 217.800 66.600 ;
        RECT 219.600 65.700 223.200 66.600 ;
        RECT 207.000 64.800 209.700 65.700 ;
        RECT 203.400 63.000 209.700 64.800 ;
        RECT 214.200 63.900 216.900 65.700 ;
        RECT 220.500 63.900 223.200 65.700 ;
        RECT 203.400 62.100 210.600 63.000 ;
        RECT 203.400 57.600 206.100 62.100 ;
        RECT 207.900 61.200 210.600 62.100 ;
        RECT 214.200 62.100 224.100 63.900 ;
        RECT 208.800 59.400 211.500 61.200 ;
        RECT 214.200 60.300 216.900 62.100 ;
        RECT 220.500 60.300 223.200 61.200 ;
        RECT 214.200 59.400 217.800 60.300 ;
        RECT 219.600 59.400 223.200 60.300 ;
        RECT 232.200 59.400 234.900 66.600 ;
        RECT 238.500 65.700 242.100 66.600 ;
        RECT 244.800 65.700 248.400 66.600 ;
        RECT 238.500 63.900 241.200 65.700 ;
        RECT 237.600 62.100 241.200 63.900 ;
        RECT 238.500 60.300 241.200 62.100 ;
        RECT 245.700 64.800 248.400 65.700 ;
        RECT 245.700 61.200 249.300 64.800 ;
        RECT 245.700 60.300 248.400 61.200 ;
        RECT 238.500 59.400 242.100 60.300 ;
        RECT 244.800 59.400 248.400 60.300 ;
        RECT 209.700 57.600 212.400 59.400 ;
        RECT 215.100 58.500 222.300 59.400 ;
        RECT 232.200 58.500 236.700 59.400 ;
        RECT 239.400 58.500 247.500 59.400 ;
        RECT 216.900 57.600 220.500 58.500 ;
        RECT 233.100 57.600 236.700 58.500 ;
        RECT 241.200 57.600 245.700 58.500 ;
        RECT 15.300 45.900 17.100 46.800 ;
        RECT 14.400 44.100 17.100 45.900 ;
        RECT 13.500 42.300 19.800 44.100 ;
        RECT 21.600 43.200 24.300 48.600 ;
        RECT 25.200 43.200 28.800 44.100 ;
        RECT 36.000 43.200 40.500 44.100 ;
        RECT 45.000 43.200 47.700 44.100 ;
        RECT 49.500 43.200 53.100 44.100 ;
        RECT 21.600 42.300 30.600 43.200 ;
        RECT 14.400 36.000 17.100 42.300 ;
        RECT 21.600 41.400 25.200 42.300 ;
        RECT 14.400 35.100 18.000 36.000 ;
        RECT 15.300 34.200 19.800 35.100 ;
        RECT 16.200 33.300 19.800 34.200 ;
        RECT 21.600 33.300 24.300 41.400 ;
        RECT 27.900 33.300 30.600 42.300 ;
        RECT 34.200 42.300 42.300 43.200 ;
        RECT 34.200 41.400 36.900 42.300 ;
        RECT 33.300 40.500 36.000 41.400 ;
        RECT 39.600 40.500 42.300 42.300 ;
        RECT 38.700 39.600 42.300 40.500 ;
        RECT 35.100 38.700 42.300 39.600 ;
        RECT 33.300 37.800 37.800 38.700 ;
        RECT 33.300 36.000 36.000 37.800 ;
        RECT 39.600 36.000 42.300 38.700 ;
        RECT 33.300 35.100 36.900 36.000 ;
        RECT 38.700 35.100 42.300 36.000 ;
        RECT 45.000 42.300 54.000 43.200 ;
        RECT 45.000 40.500 48.600 42.300 ;
        RECT 51.300 41.400 54.900 42.300 ;
        RECT 33.300 34.200 43.200 35.100 ;
        RECT 35.100 33.300 38.700 34.200 ;
        RECT 40.500 33.300 43.200 34.200 ;
        RECT 45.000 33.300 47.700 40.500 ;
        RECT 52.200 33.300 54.900 41.400 ;
        RECT 57.600 40.500 60.300 48.600 ;
        RECT 74.700 46.800 79.200 48.600 ;
        RECT 84.600 46.800 89.100 48.600 ;
        RECT 105.300 46.800 106.200 47.700 ;
        RECT 63.900 43.200 66.600 44.100 ;
        RECT 74.700 43.200 80.100 46.800 ;
        RECT 83.700 44.100 89.100 46.800 ;
        RECT 104.400 45.900 106.200 46.800 ;
        RECT 103.500 44.100 106.200 45.900 ;
        RECT 110.700 44.100 113.400 46.800 ;
        RECT 83.700 43.200 85.500 44.100 ;
        RECT 63.000 42.300 65.700 43.200 ;
        RECT 62.100 41.400 64.800 42.300 ;
        RECT 61.200 40.500 63.900 41.400 ;
        RECT 57.600 38.700 63.900 40.500 ;
        RECT 57.600 37.800 64.800 38.700 ;
        RECT 57.600 36.900 61.200 37.800 ;
        RECT 62.100 36.900 64.800 37.800 ;
        RECT 57.600 33.300 60.300 36.900 ;
        RECT 63.000 36.000 65.700 36.900 ;
        RECT 63.000 35.100 66.600 36.000 ;
        RECT 63.900 34.200 66.600 35.100 ;
        RECT 64.800 33.300 67.500 34.200 ;
        RECT 74.700 33.300 77.400 43.200 ;
        RECT 78.300 41.400 81.000 43.200 ;
        RECT 79.200 40.500 81.000 41.400 ;
        RECT 82.800 41.400 85.500 43.200 ;
        RECT 79.200 39.600 81.900 40.500 ;
        RECT 82.800 39.600 84.600 41.400 ;
        RECT 79.200 37.800 84.600 39.600 ;
        RECT 80.100 36.900 84.600 37.800 ;
        RECT 80.100 33.300 83.700 36.900 ;
        RECT 86.400 33.300 89.100 44.100 ;
        RECT 93.600 43.200 99.000 44.100 ;
        RECT 92.700 42.300 99.900 43.200 ;
        RECT 102.600 42.300 108.000 44.100 ;
        RECT 108.900 42.300 115.200 44.100 ;
        RECT 91.800 40.500 94.500 42.300 ;
        RECT 97.200 41.400 100.800 42.300 ;
        RECT 98.100 40.500 100.800 41.400 ;
        RECT 96.300 39.600 100.800 40.500 ;
        RECT 92.700 38.700 100.800 39.600 ;
        RECT 91.800 37.800 95.400 38.700 ;
        RECT 90.900 35.100 94.500 37.800 ;
        RECT 98.100 36.900 100.800 38.700 ;
        RECT 97.200 35.100 100.800 36.900 ;
        RECT 91.800 34.200 100.800 35.100 ;
        RECT 103.500 35.100 106.200 42.300 ;
        RECT 110.700 35.100 113.400 42.300 ;
        RECT 128.700 36.900 131.400 48.600 ;
        RECT 137.700 38.700 140.400 48.600 ;
        RECT 151.200 45.900 153.900 48.600 ;
        RECT 166.500 47.700 174.600 48.600 ;
        RECT 166.500 45.900 176.400 47.700 ;
        RECT 136.800 36.900 140.400 38.700 ;
        RECT 143.100 43.200 145.800 44.100 ;
        RECT 146.700 43.200 149.400 44.100 ;
        RECT 143.100 42.300 149.400 43.200 ;
        RECT 143.100 40.500 146.700 42.300 ;
        RECT 128.700 36.000 132.300 36.900 ;
        RECT 135.900 36.000 139.500 36.900 ;
        RECT 103.500 34.200 108.000 35.100 ;
        RECT 110.700 34.200 115.200 35.100 ;
        RECT 92.700 33.300 96.300 34.200 ;
        RECT 98.100 33.300 100.800 34.200 ;
        RECT 104.400 33.300 108.000 34.200 ;
        RECT 111.600 33.300 115.200 34.200 ;
        RECT 117.000 33.300 119.700 36.000 ;
        RECT 129.600 35.100 139.500 36.000 ;
        RECT 129.600 34.200 138.600 35.100 ;
        RECT 131.400 33.300 136.800 34.200 ;
        RECT 143.100 33.300 145.800 40.500 ;
        RECT 151.200 33.300 153.900 44.100 ;
        RECT 166.500 41.400 169.200 45.900 ;
        RECT 173.700 45.000 177.300 45.900 ;
        RECT 174.600 42.300 177.300 45.000 ;
        RECT 181.800 43.200 187.200 44.100 ;
        RECT 189.900 43.200 192.600 44.100 ;
        RECT 180.900 42.300 188.100 43.200 ;
        RECT 173.700 41.400 177.300 42.300 ;
        RECT 166.500 39.600 176.400 41.400 ;
        RECT 180.000 40.500 182.700 42.300 ;
        RECT 185.400 40.500 189.000 42.300 ;
        RECT 190.800 40.500 193.500 43.200 ;
        RECT 196.200 40.500 199.800 44.100 ;
        RECT 203.400 43.200 206.100 44.100 ;
        RECT 209.700 43.200 213.300 44.100 ;
        RECT 202.500 40.500 205.200 43.200 ;
        RECT 207.900 42.300 215.100 43.200 ;
        RECT 207.000 41.400 210.600 42.300 ;
        RECT 212.400 41.400 216.000 42.300 ;
        RECT 184.500 39.600 189.000 40.500 ;
        RECT 166.500 38.700 174.600 39.600 ;
        RECT 180.900 38.700 189.000 39.600 ;
        RECT 156.600 33.300 159.300 36.000 ;
        RECT 166.500 33.300 169.200 38.700 ;
        RECT 180.000 37.800 183.600 38.700 ;
        RECT 179.100 36.900 182.700 37.800 ;
        RECT 179.100 36.000 181.800 36.900 ;
        RECT 185.400 36.000 189.000 38.700 ;
        RECT 191.700 39.600 193.500 40.500 ;
        RECT 191.700 37.800 194.400 39.600 ;
        RECT 195.300 38.700 200.700 40.500 ;
        RECT 202.500 39.600 204.300 40.500 ;
        RECT 195.300 37.800 197.100 38.700 ;
        RECT 191.700 36.900 197.100 37.800 ;
        RECT 179.100 35.100 182.700 36.000 ;
        RECT 184.500 35.100 189.000 36.000 ;
        RECT 180.000 34.200 189.000 35.100 ;
        RECT 192.600 35.100 197.100 36.900 ;
        RECT 198.900 37.800 200.700 38.700 ;
        RECT 201.600 37.800 204.300 39.600 ;
        RECT 207.000 39.600 209.700 41.400 ;
        RECT 213.300 39.600 216.000 41.400 ;
        RECT 207.000 37.800 216.900 39.600 ;
        RECT 198.900 35.100 203.400 37.800 ;
        RECT 207.000 36.000 209.700 37.800 ;
        RECT 213.300 36.000 216.000 36.900 ;
        RECT 207.000 35.100 210.600 36.000 ;
        RECT 212.400 35.100 216.000 36.000 ;
        RECT 192.600 34.200 196.200 35.100 ;
        RECT 180.900 33.300 184.500 34.200 ;
        RECT 186.300 33.300 189.000 34.200 ;
        RECT 193.500 33.300 196.200 34.200 ;
        RECT 199.800 34.200 203.400 35.100 ;
        RECT 207.900 34.200 215.100 35.100 ;
        RECT 199.800 33.300 202.500 34.200 ;
        RECT 209.700 33.300 213.300 34.200 ;
        RECT 218.700 33.300 221.400 48.600 ;
        RECT 235.800 47.700 244.800 48.600 ;
        RECT 235.800 46.800 245.700 47.700 ;
        RECT 235.800 45.900 246.600 46.800 ;
        RECT 250.200 45.900 252.900 48.600 ;
        RECT 235.800 36.000 238.500 45.900 ;
        RECT 243.900 45.000 247.500 45.900 ;
        RECT 244.800 44.100 247.500 45.000 ;
        RECT 244.800 42.300 248.400 44.100 ;
        RECT 245.700 39.600 248.400 42.300 ;
        RECT 244.800 37.800 248.400 39.600 ;
        RECT 244.800 36.900 247.500 37.800 ;
        RECT 243.900 36.000 247.500 36.900 ;
        RECT 224.100 33.300 226.800 36.000 ;
        RECT 235.800 35.100 246.600 36.000 ;
        RECT 235.800 34.200 245.700 35.100 ;
        RECT 235.800 33.300 243.900 34.200 ;
        RECT 250.200 33.300 252.900 44.100 ;
        RECT 258.300 43.200 262.800 44.100 ;
        RECT 270.000 43.200 273.600 44.100 ;
        RECT 274.500 43.200 278.100 44.100 ;
        RECT 282.600 43.200 287.100 44.100 ;
        RECT 257.400 42.300 263.700 43.200 ;
        RECT 268.200 42.300 278.100 43.200 ;
        RECT 281.700 42.300 288.900 43.200 ;
        RECT 256.500 41.400 259.200 42.300 ;
        RECT 261.900 41.400 264.600 42.300 ;
        RECT 268.200 41.400 270.900 42.300 ;
        RECT 273.600 41.400 278.100 42.300 ;
        RECT 280.800 41.400 283.500 42.300 ;
        RECT 286.200 41.400 289.800 42.300 ;
        RECT 255.600 40.500 259.200 41.400 ;
        RECT 255.600 39.600 258.300 40.500 ;
        RECT 262.800 39.600 265.500 41.400 ;
        RECT 255.600 37.800 265.500 39.600 ;
        RECT 267.300 40.500 270.900 41.400 ;
        RECT 255.600 36.000 258.300 37.800 ;
        RECT 267.300 36.900 270.000 40.500 ;
        RECT 274.500 39.600 278.100 41.400 ;
        RECT 275.400 37.800 278.100 39.600 ;
        RECT 262.800 36.000 265.500 36.900 ;
        RECT 267.300 36.000 270.900 36.900 ;
        RECT 274.500 36.000 278.100 37.800 ;
        RECT 279.900 36.000 282.600 41.400 ;
        RECT 287.100 40.500 289.800 41.400 ;
        RECT 288.000 36.900 290.700 40.500 ;
        RECT 287.100 36.000 289.800 36.900 ;
        RECT 256.500 35.100 259.200 36.000 ;
        RECT 261.900 35.100 264.600 36.000 ;
        RECT 268.200 35.100 270.900 36.000 ;
        RECT 273.600 35.100 278.100 36.000 ;
        RECT 280.800 35.100 283.500 36.000 ;
        RECT 286.200 35.100 289.800 36.000 ;
        RECT 257.400 34.200 263.700 35.100 ;
        RECT 268.200 34.200 278.100 35.100 ;
        RECT 281.700 34.200 288.900 35.100 ;
        RECT 258.300 33.300 262.800 34.200 ;
        RECT 270.000 33.300 273.600 34.200 ;
        RECT 117.900 31.500 119.700 33.300 ;
        RECT 157.500 31.500 159.300 33.300 ;
        RECT 225.000 31.500 226.800 33.300 ;
        RECT 274.500 32.400 278.100 34.200 ;
        RECT 282.600 33.300 287.100 34.200 ;
        RECT 292.500 33.300 295.200 36.000 ;
        RECT 117.900 30.600 118.800 31.500 ;
        RECT 157.500 30.600 158.400 31.500 ;
        RECT 225.000 30.600 225.900 31.500 ;
        RECT 267.300 30.600 270.900 31.500 ;
        RECT 274.500 30.600 277.200 32.400 ;
        RECT 293.400 31.500 295.200 33.300 ;
        RECT 293.400 30.600 294.300 31.500 ;
        RECT 268.200 29.700 276.300 30.600 ;
        RECT 270.000 28.800 275.400 29.700 ;
        RECT 84.600 21.600 89.100 23.400 ;
        RECT 94.500 21.600 99.000 23.400 ;
        RECT 84.600 18.000 90.000 21.600 ;
        RECT 93.600 18.900 99.000 21.600 ;
        RECT 93.600 18.000 95.400 18.900 ;
        RECT 84.600 8.100 87.300 18.000 ;
        RECT 88.200 16.200 90.900 18.000 ;
        RECT 89.100 15.300 90.900 16.200 ;
        RECT 92.700 16.200 95.400 18.000 ;
        RECT 89.100 14.400 91.800 15.300 ;
        RECT 92.700 14.400 94.500 16.200 ;
        RECT 89.100 12.600 94.500 14.400 ;
        RECT 90.000 11.700 94.500 12.600 ;
        RECT 90.000 8.100 93.600 11.700 ;
        RECT 96.300 8.100 99.000 18.900 ;
        RECT 103.500 18.000 108.900 18.900 ;
        RECT 113.400 18.000 115.200 18.900 ;
        RECT 116.100 18.000 119.700 18.900 ;
        RECT 123.300 18.000 126.900 18.900 ;
        RECT 127.800 18.000 131.400 23.400 ;
        RECT 134.100 20.700 136.800 23.400 ;
        RECT 102.600 17.100 109.800 18.000 ;
        RECT 113.400 17.100 118.800 18.000 ;
        RECT 121.500 17.100 131.400 18.000 ;
        RECT 101.700 15.300 104.400 17.100 ;
        RECT 107.100 16.200 110.700 17.100 ;
        RECT 108.000 15.300 110.700 16.200 ;
        RECT 106.200 14.400 110.700 15.300 ;
        RECT 102.600 13.500 110.700 14.400 ;
        RECT 101.700 12.600 105.300 13.500 ;
        RECT 100.800 9.900 104.400 12.600 ;
        RECT 108.000 11.700 110.700 13.500 ;
        RECT 107.100 9.900 110.700 11.700 ;
        RECT 101.700 9.000 110.700 9.900 ;
        RECT 102.600 8.100 106.200 9.000 ;
        RECT 108.000 8.100 110.700 9.000 ;
        RECT 113.400 16.200 117.000 17.100 ;
        RECT 121.500 16.200 124.200 17.100 ;
        RECT 126.900 16.200 131.400 17.100 ;
        RECT 113.400 8.100 116.100 16.200 ;
        RECT 120.600 15.300 124.200 16.200 ;
        RECT 120.600 11.700 123.300 15.300 ;
        RECT 120.600 10.800 124.200 11.700 ;
        RECT 127.800 10.800 131.400 16.200 ;
        RECT 121.500 9.900 124.200 10.800 ;
        RECT 126.900 9.900 131.400 10.800 ;
        RECT 122.400 9.000 131.400 9.900 ;
        RECT 123.300 8.100 126.900 9.000 ;
        RECT 128.700 8.100 131.400 9.000 ;
        RECT 134.100 8.100 136.800 18.900 ;
        RECT 153.000 18.000 157.500 18.900 ;
        RECT 162.000 18.000 164.700 18.900 ;
        RECT 166.500 18.000 170.100 18.900 ;
        RECT 176.400 18.000 180.000 18.900 ;
        RECT 181.800 18.000 184.500 23.400 ;
        RECT 151.200 17.100 159.300 18.000 ;
        RECT 151.200 16.200 153.900 17.100 ;
        RECT 150.300 15.300 153.000 16.200 ;
        RECT 156.600 15.300 159.300 17.100 ;
        RECT 155.700 14.400 159.300 15.300 ;
        RECT 152.100 13.500 159.300 14.400 ;
        RECT 150.300 12.600 154.800 13.500 ;
        RECT 150.300 10.800 153.000 12.600 ;
        RECT 156.600 10.800 159.300 13.500 ;
        RECT 139.500 8.100 142.200 10.800 ;
        RECT 150.300 9.900 153.900 10.800 ;
        RECT 155.700 9.900 159.300 10.800 ;
        RECT 162.000 17.100 171.000 18.000 ;
        RECT 175.500 17.100 184.500 18.000 ;
        RECT 162.000 15.300 165.600 17.100 ;
        RECT 168.300 16.200 171.900 17.100 ;
        RECT 150.300 9.000 160.200 9.900 ;
        RECT 152.100 8.100 155.700 9.000 ;
        RECT 157.500 8.100 160.200 9.000 ;
        RECT 162.000 8.100 164.700 15.300 ;
        RECT 169.200 8.100 171.900 16.200 ;
        RECT 174.600 16.200 178.200 17.100 ;
        RECT 180.900 16.200 184.500 17.100 ;
        RECT 174.600 10.800 177.300 16.200 ;
        RECT 181.800 10.800 184.500 16.200 ;
        RECT 174.600 9.900 178.200 10.800 ;
        RECT 180.900 9.900 184.500 10.800 ;
        RECT 175.500 9.000 184.500 9.900 ;
        RECT 176.400 8.100 180.900 9.000 ;
        RECT 181.800 8.100 184.500 9.000 ;
        RECT 193.500 10.800 196.200 23.400 ;
        RECT 205.200 20.700 207.900 23.400 ;
        RECT 193.500 8.100 203.400 10.800 ;
        RECT 205.200 8.100 207.900 18.900 ;
        RECT 211.500 8.100 214.200 23.400 ;
        RECT 216.000 17.100 218.700 18.900 ;
        RECT 224.100 18.000 226.800 18.900 ;
        RECT 216.000 16.200 219.600 17.100 ;
        RECT 216.900 14.400 219.600 16.200 ;
        RECT 223.200 15.300 225.900 18.000 ;
        RECT 217.800 11.700 220.500 14.400 ;
        RECT 222.300 13.500 225.000 15.300 ;
        RECT 221.400 12.600 225.000 13.500 ;
        RECT 221.400 11.700 224.100 12.600 ;
        RECT 218.700 10.800 224.100 11.700 ;
        RECT 218.700 9.900 223.200 10.800 ;
        RECT 219.600 8.100 223.200 9.900 ;
        RECT 140.400 6.300 142.200 8.100 ;
        RECT 219.600 6.300 222.300 8.100 ;
        RECT 140.400 5.400 141.300 6.300 ;
        RECT 218.700 5.400 222.300 6.300 ;
        RECT 216.900 4.500 221.400 5.400 ;
        RECT 216.900 3.600 220.500 4.500 ;
  END
END asic_hat_logo
END LIBRARY

