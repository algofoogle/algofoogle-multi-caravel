VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 969.855 BY 987.775 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 920.640 4.000 921.200 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 483.840 4.000 484.400 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.200 4.000 487.760 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 500.640 4.000 501.200 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 504.000 4.000 504.560 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 551.040 4.000 551.600 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.400 4.000 554.960 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.120 4.000 561.680 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 564.480 4.000 565.040 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 672.000 4.000 672.560 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 661.920 4.000 662.480 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 722.400 4.000 722.960 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 688.800 4.000 689.360 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 719.040 4.000 719.600 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 715.680 4.000 716.240 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 685.440 4.000 686.000 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 682.080 4.000 682.640 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 678.720 4.000 679.280 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 675.360 4.000 675.920 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 665.280 4.000 665.840 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 668.640 4.000 669.200 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 591.360 4.000 591.920 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 594.720 4.000 595.280 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.880 4.000 615.440 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 658.560 4.000 659.120 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.040 4.000 635.600 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 621.600 4.000 622.160 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 648.480 4.000 649.040 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 628.320 4.000 628.880 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 651.840 4.000 652.400 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 618.240 4.000 618.800 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 624.960 4.000 625.520 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 611.520 4.000 612.080 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 497.280 4.000 497.840 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.240 4.000 534.800 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 524.160 4.000 524.720 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 540.960 4.000 541.520 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 530.880 4.000 531.440 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.320 4.000 544.880 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 4.000 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 983.775 608.720 987.775 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 705.600 4.000 706.160 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 712.320 4.000 712.880 ;
    END
  END i_reg_mosi
  PIN i_reg_outs_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 507.360 4.000 507.920 ;
    END
  END i_reg_outs_enb
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 708.960 4.000 709.520 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.600 4.000 538.160 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 520.800 4.000 521.360 ;
    END
  END i_reset_lock_b
  PIN i_spare_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END i_spare_0
  PIN i_spare_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END i_spare_1
  PIN i_test_uc2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 702.240 4.000 702.800 ;
    END
  END i_test_uc2
  PIN i_test_wci
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 695.520 4.000 696.080 ;
    END
  END i_test_wci
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 493.920 4.000 494.480 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 557.760 4.000 558.320 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 692.160 4.000 692.720 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 581.280 4.000 581.840 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.920 4.000 578.480 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 698.880 4.000 699.440 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 584.640 4.000 585.200 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 567.840 4.000 568.400 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 571.200 4.000 571.760 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 655.200 4.000 655.760 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 631.680 4.000 632.240 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.120 4.000 645.680 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 510.720 4.000 511.280 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 527.520 4.000 528.080 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 480.480 4.000 481.040 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 0.000 464.240 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 983.775 773.360 987.775 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 0.000 843.920 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 983.775 672.560 987.775 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 547.680 4.000 548.240 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 641.760 4.000 642.320 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 0.000 927.920 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 0.000 561.680 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 833.280 983.775 833.840 987.775 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 0.000 554.960 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 965.855 856.800 969.855 857.360 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 965.855 957.600 969.855 958.160 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 0.000 796.880 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 638.400 4.000 638.960 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.080 4.000 514.640 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 983.775 182.000 987.775 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 983.775 14.000 987.775 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 930.720 0.000 931.280 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 4.000 27.440 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 604.800 4.000 605.360 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 588.000 4.000 588.560 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 0.000 917.840 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 490.560 4.000 491.120 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 608.160 4.000 608.720 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 598.080 4.000 598.640 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 601.440 4.000 602.000 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 517.440 4.000 518.000 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 983.775 91.280 987.775 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 4.000 24.080 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 983.775 706.160 987.775 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 806.400 0.000 806.960 4.000 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 0.000 954.800 4.000 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 4.000 47.600 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 965.855 967.680 969.855 968.240 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 0.000 907.760 4.000 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 983.775 111.440 987.775 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 983.775 689.360 987.775 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 965.855 954.240 969.855 954.800 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 4.000 30.800 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 0.000 417.200 4.000 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END ones[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 968.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 968.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 968.540 ;
    END
  END vss
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 965.855 960.960 969.855 961.520 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 0.000 850.640 4.000 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 983.775 712.880 987.775 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 983.775 776.720 987.775 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 983.775 632.240 987.775 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 0.000 575.120 4.000 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 965.855 964.320 969.855 964.880 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 983.775 743.120 987.775 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 983.775 770.000 987.775 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 0.000 672.560 4.000 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 983.775 669.200 987.775 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 965.855 944.160 969.855 944.720 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 983.775 790.160 987.775 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 0.000 944.720 4.000 ;
    END
  END zeros[9]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 962.640 968.540 ;
      LAYER Metal2 ;
        RECT 7.980 983.475 13.140 984.340 ;
        RECT 14.300 983.475 90.420 984.340 ;
        RECT 91.580 983.475 110.580 984.340 ;
        RECT 111.740 983.475 181.140 984.340 ;
        RECT 182.300 983.475 607.860 984.340 ;
        RECT 609.020 983.475 631.380 984.340 ;
        RECT 632.540 983.475 668.340 984.340 ;
        RECT 669.500 983.475 671.700 984.340 ;
        RECT 672.860 983.475 688.500 984.340 ;
        RECT 689.660 983.475 705.300 984.340 ;
        RECT 706.460 983.475 712.020 984.340 ;
        RECT 713.180 983.475 742.260 984.340 ;
        RECT 743.420 983.475 769.140 984.340 ;
        RECT 770.300 983.475 772.500 984.340 ;
        RECT 773.660 983.475 775.860 984.340 ;
        RECT 777.020 983.475 789.300 984.340 ;
        RECT 790.460 983.475 832.980 984.340 ;
        RECT 834.140 983.475 960.820 984.340 ;
        RECT 7.980 4.300 960.820 983.475 ;
        RECT 7.980 4.000 130.740 4.300 ;
        RECT 131.900 4.000 251.700 4.300 ;
        RECT 252.860 4.000 255.060 4.300 ;
        RECT 256.220 4.000 261.780 4.300 ;
        RECT 262.940 4.000 278.580 4.300 ;
        RECT 279.740 4.000 416.340 4.300 ;
        RECT 417.500 4.000 463.380 4.300 ;
        RECT 464.540 4.000 554.100 4.300 ;
        RECT 555.260 4.000 560.820 4.300 ;
        RECT 561.980 4.000 574.260 4.300 ;
        RECT 575.420 4.000 671.700 4.300 ;
        RECT 672.860 4.000 796.020 4.300 ;
        RECT 797.180 4.000 806.100 4.300 ;
        RECT 807.260 4.000 843.060 4.300 ;
        RECT 844.220 4.000 849.780 4.300 ;
        RECT 850.940 4.000 906.900 4.300 ;
        RECT 908.060 4.000 916.980 4.300 ;
        RECT 918.140 4.000 927.060 4.300 ;
        RECT 928.220 4.000 930.420 4.300 ;
        RECT 931.580 4.000 943.860 4.300 ;
        RECT 945.020 4.000 953.940 4.300 ;
        RECT 955.100 4.000 960.820 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 967.380 965.555 968.380 ;
        RECT 4.000 965.180 965.855 967.380 ;
        RECT 4.000 964.020 965.555 965.180 ;
        RECT 4.000 961.820 965.855 964.020 ;
        RECT 4.000 960.660 965.555 961.820 ;
        RECT 4.000 958.460 965.855 960.660 ;
        RECT 4.000 957.300 965.555 958.460 ;
        RECT 4.000 955.100 965.855 957.300 ;
        RECT 4.000 953.940 965.555 955.100 ;
        RECT 4.000 945.020 965.855 953.940 ;
        RECT 4.000 943.860 965.555 945.020 ;
        RECT 4.000 921.500 965.855 943.860 ;
        RECT 4.300 920.340 965.855 921.500 ;
        RECT 4.000 857.660 965.855 920.340 ;
        RECT 4.000 856.500 965.555 857.660 ;
        RECT 4.000 723.260 965.855 856.500 ;
        RECT 4.300 722.100 965.855 723.260 ;
        RECT 4.000 719.900 965.855 722.100 ;
        RECT 4.300 718.740 965.855 719.900 ;
        RECT 4.000 716.540 965.855 718.740 ;
        RECT 4.300 715.380 965.855 716.540 ;
        RECT 4.000 713.180 965.855 715.380 ;
        RECT 4.300 712.020 965.855 713.180 ;
        RECT 4.000 709.820 965.855 712.020 ;
        RECT 4.300 708.660 965.855 709.820 ;
        RECT 4.000 706.460 965.855 708.660 ;
        RECT 4.300 705.300 965.855 706.460 ;
        RECT 4.000 703.100 965.855 705.300 ;
        RECT 4.300 701.940 965.855 703.100 ;
        RECT 4.000 699.740 965.855 701.940 ;
        RECT 4.300 698.580 965.855 699.740 ;
        RECT 4.000 696.380 965.855 698.580 ;
        RECT 4.300 695.220 965.855 696.380 ;
        RECT 4.000 693.020 965.855 695.220 ;
        RECT 4.300 691.860 965.855 693.020 ;
        RECT 4.000 689.660 965.855 691.860 ;
        RECT 4.300 688.500 965.855 689.660 ;
        RECT 4.000 686.300 965.855 688.500 ;
        RECT 4.300 685.140 965.855 686.300 ;
        RECT 4.000 682.940 965.855 685.140 ;
        RECT 4.300 681.780 965.855 682.940 ;
        RECT 4.000 679.580 965.855 681.780 ;
        RECT 4.300 678.420 965.855 679.580 ;
        RECT 4.000 676.220 965.855 678.420 ;
        RECT 4.300 675.060 965.855 676.220 ;
        RECT 4.000 672.860 965.855 675.060 ;
        RECT 4.300 671.700 965.855 672.860 ;
        RECT 4.000 669.500 965.855 671.700 ;
        RECT 4.300 668.340 965.855 669.500 ;
        RECT 4.000 666.140 965.855 668.340 ;
        RECT 4.300 664.980 965.855 666.140 ;
        RECT 4.000 662.780 965.855 664.980 ;
        RECT 4.300 661.620 965.855 662.780 ;
        RECT 4.000 659.420 965.855 661.620 ;
        RECT 4.300 658.260 965.855 659.420 ;
        RECT 4.000 656.060 965.855 658.260 ;
        RECT 4.300 654.900 965.855 656.060 ;
        RECT 4.000 652.700 965.855 654.900 ;
        RECT 4.300 651.540 965.855 652.700 ;
        RECT 4.000 649.340 965.855 651.540 ;
        RECT 4.300 648.180 965.855 649.340 ;
        RECT 4.000 645.980 965.855 648.180 ;
        RECT 4.300 644.820 965.855 645.980 ;
        RECT 4.000 642.620 965.855 644.820 ;
        RECT 4.300 641.460 965.855 642.620 ;
        RECT 4.000 639.260 965.855 641.460 ;
        RECT 4.300 638.100 965.855 639.260 ;
        RECT 4.000 635.900 965.855 638.100 ;
        RECT 4.300 634.740 965.855 635.900 ;
        RECT 4.000 632.540 965.855 634.740 ;
        RECT 4.300 631.380 965.855 632.540 ;
        RECT 4.000 629.180 965.855 631.380 ;
        RECT 4.300 628.020 965.855 629.180 ;
        RECT 4.000 625.820 965.855 628.020 ;
        RECT 4.300 624.660 965.855 625.820 ;
        RECT 4.000 622.460 965.855 624.660 ;
        RECT 4.300 621.300 965.855 622.460 ;
        RECT 4.000 619.100 965.855 621.300 ;
        RECT 4.300 617.940 965.855 619.100 ;
        RECT 4.000 615.740 965.855 617.940 ;
        RECT 4.300 614.580 965.855 615.740 ;
        RECT 4.000 612.380 965.855 614.580 ;
        RECT 4.300 611.220 965.855 612.380 ;
        RECT 4.000 609.020 965.855 611.220 ;
        RECT 4.300 607.860 965.855 609.020 ;
        RECT 4.000 605.660 965.855 607.860 ;
        RECT 4.300 604.500 965.855 605.660 ;
        RECT 4.000 602.300 965.855 604.500 ;
        RECT 4.300 601.140 965.855 602.300 ;
        RECT 4.000 598.940 965.855 601.140 ;
        RECT 4.300 597.780 965.855 598.940 ;
        RECT 4.000 595.580 965.855 597.780 ;
        RECT 4.300 594.420 965.855 595.580 ;
        RECT 4.000 592.220 965.855 594.420 ;
        RECT 4.300 591.060 965.855 592.220 ;
        RECT 4.000 588.860 965.855 591.060 ;
        RECT 4.300 587.700 965.855 588.860 ;
        RECT 4.000 585.500 965.855 587.700 ;
        RECT 4.300 584.340 965.855 585.500 ;
        RECT 4.000 582.140 965.855 584.340 ;
        RECT 4.300 580.980 965.855 582.140 ;
        RECT 4.000 578.780 965.855 580.980 ;
        RECT 4.300 577.620 965.855 578.780 ;
        RECT 4.000 575.420 965.855 577.620 ;
        RECT 4.300 574.260 965.855 575.420 ;
        RECT 4.000 572.060 965.855 574.260 ;
        RECT 4.300 570.900 965.855 572.060 ;
        RECT 4.000 568.700 965.855 570.900 ;
        RECT 4.300 567.540 965.855 568.700 ;
        RECT 4.000 565.340 965.855 567.540 ;
        RECT 4.300 564.180 965.855 565.340 ;
        RECT 4.000 561.980 965.855 564.180 ;
        RECT 4.300 560.820 965.855 561.980 ;
        RECT 4.000 558.620 965.855 560.820 ;
        RECT 4.300 557.460 965.855 558.620 ;
        RECT 4.000 555.260 965.855 557.460 ;
        RECT 4.300 554.100 965.855 555.260 ;
        RECT 4.000 551.900 965.855 554.100 ;
        RECT 4.300 550.740 965.855 551.900 ;
        RECT 4.000 548.540 965.855 550.740 ;
        RECT 4.300 547.380 965.855 548.540 ;
        RECT 4.000 545.180 965.855 547.380 ;
        RECT 4.300 544.020 965.855 545.180 ;
        RECT 4.000 541.820 965.855 544.020 ;
        RECT 4.300 540.660 965.855 541.820 ;
        RECT 4.000 538.460 965.855 540.660 ;
        RECT 4.300 537.300 965.855 538.460 ;
        RECT 4.000 535.100 965.855 537.300 ;
        RECT 4.300 533.940 965.855 535.100 ;
        RECT 4.000 531.740 965.855 533.940 ;
        RECT 4.300 530.580 965.855 531.740 ;
        RECT 4.000 528.380 965.855 530.580 ;
        RECT 4.300 527.220 965.855 528.380 ;
        RECT 4.000 525.020 965.855 527.220 ;
        RECT 4.300 523.860 965.855 525.020 ;
        RECT 4.000 521.660 965.855 523.860 ;
        RECT 4.300 520.500 965.855 521.660 ;
        RECT 4.000 518.300 965.855 520.500 ;
        RECT 4.300 517.140 965.855 518.300 ;
        RECT 4.000 514.940 965.855 517.140 ;
        RECT 4.300 513.780 965.855 514.940 ;
        RECT 4.000 511.580 965.855 513.780 ;
        RECT 4.300 510.420 965.855 511.580 ;
        RECT 4.000 508.220 965.855 510.420 ;
        RECT 4.300 507.060 965.855 508.220 ;
        RECT 4.000 504.860 965.855 507.060 ;
        RECT 4.300 503.700 965.855 504.860 ;
        RECT 4.000 501.500 965.855 503.700 ;
        RECT 4.300 500.340 965.855 501.500 ;
        RECT 4.000 498.140 965.855 500.340 ;
        RECT 4.300 496.980 965.855 498.140 ;
        RECT 4.000 494.780 965.855 496.980 ;
        RECT 4.300 493.620 965.855 494.780 ;
        RECT 4.000 491.420 965.855 493.620 ;
        RECT 4.300 490.260 965.855 491.420 ;
        RECT 4.000 488.060 965.855 490.260 ;
        RECT 4.300 486.900 965.855 488.060 ;
        RECT 4.000 484.700 965.855 486.900 ;
        RECT 4.300 483.540 965.855 484.700 ;
        RECT 4.000 481.340 965.855 483.540 ;
        RECT 4.300 480.180 965.855 481.340 ;
        RECT 4.000 54.620 965.855 480.180 ;
        RECT 4.300 53.460 965.855 54.620 ;
        RECT 4.000 47.900 965.855 53.460 ;
        RECT 4.300 46.740 965.855 47.900 ;
        RECT 4.000 44.540 965.855 46.740 ;
        RECT 4.300 43.380 965.855 44.540 ;
        RECT 4.000 34.460 965.855 43.380 ;
        RECT 4.300 33.300 965.855 34.460 ;
        RECT 4.000 31.100 965.855 33.300 ;
        RECT 4.300 29.940 965.855 31.100 ;
        RECT 4.000 27.740 965.855 29.940 ;
        RECT 4.300 26.580 965.855 27.740 ;
        RECT 4.000 24.380 965.855 26.580 ;
        RECT 4.300 23.220 965.855 24.380 ;
        RECT 4.000 21.020 965.855 23.220 ;
        RECT 4.300 19.860 965.855 21.020 ;
        RECT 4.000 15.540 965.855 19.860 ;
      LAYER Metal4 ;
        RECT 48.300 41.530 98.740 931.190 ;
        RECT 100.940 41.530 175.540 931.190 ;
        RECT 177.740 41.530 252.340 931.190 ;
        RECT 254.540 41.530 329.140 931.190 ;
        RECT 331.340 41.530 405.940 931.190 ;
        RECT 408.140 41.530 482.740 931.190 ;
        RECT 484.940 41.530 559.540 931.190 ;
        RECT 561.740 41.530 636.340 931.190 ;
        RECT 638.540 41.530 713.140 931.190 ;
        RECT 715.340 41.530 789.940 931.190 ;
        RECT 792.140 41.530 866.740 931.190 ;
        RECT 868.940 41.530 927.220 931.190 ;
  END
END top_ew_algofoogle
END LIBRARY

