magic
tech gf180mcuD
magscale 1 10
timestamp 1702221777
<< metal1 >>
rect 15138 57038 15150 57090
rect 15202 57087 15214 57090
rect 16034 57087 16046 57090
rect 15202 57041 16046 57087
rect 15202 57038 15214 57041
rect 16034 57038 16046 57041
rect 16098 57038 16110 57090
rect 44370 57038 44382 57090
rect 44434 57087 44446 57090
rect 44930 57087 44942 57090
rect 44434 57041 44942 57087
rect 44434 57038 44446 57041
rect 44930 57038 44942 57041
rect 44994 57038 45006 57090
rect 12562 56590 12574 56642
rect 12626 56639 12638 56642
rect 13122 56639 13134 56642
rect 12626 56593 13134 56639
rect 12626 56590 12638 56593
rect 13122 56590 13134 56593
rect 13186 56590 13198 56642
rect 18498 56590 18510 56642
rect 18562 56639 18574 56642
rect 18946 56639 18958 56642
rect 18562 56593 18958 56639
rect 18562 56590 18574 56593
rect 18946 56590 18958 56593
rect 19010 56590 19022 56642
rect 22082 56590 22094 56642
rect 22146 56639 22158 56642
rect 22866 56639 22878 56642
rect 22146 56593 22878 56639
rect 22146 56590 22158 56593
rect 22866 56590 22878 56593
rect 22930 56590 22942 56642
rect 23650 56590 23662 56642
rect 23714 56639 23726 56642
rect 24210 56639 24222 56642
rect 23714 56593 24222 56639
rect 23714 56590 23726 56593
rect 24210 56590 24222 56593
rect 24274 56590 24286 56642
rect 27346 56590 27358 56642
rect 27410 56639 27422 56642
rect 28354 56639 28366 56642
rect 27410 56593 28366 56639
rect 27410 56590 27422 56593
rect 28354 56590 28366 56593
rect 28418 56590 28430 56642
rect 29474 56590 29486 56642
rect 29538 56639 29550 56642
rect 30034 56639 30046 56642
rect 29538 56593 30046 56639
rect 29538 56590 29550 56593
rect 30034 56590 30046 56593
rect 30098 56590 30110 56642
rect 39218 56590 39230 56642
rect 39282 56639 39294 56642
rect 39890 56639 39902 56642
rect 39282 56593 39902 56639
rect 39282 56590 39294 56593
rect 39890 56590 39902 56593
rect 39954 56590 39966 56642
rect 54226 56590 54238 56642
rect 54290 56639 54302 56642
rect 55010 56639 55022 56642
rect 54290 56593 55022 56639
rect 54290 56590 54302 56593
rect 55010 56590 55022 56593
rect 55074 56590 55086 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 4622 56306 4674 56318
rect 4622 56242 4674 56254
rect 4958 56306 5010 56318
rect 4958 56242 5010 56254
rect 6974 56306 7026 56318
rect 6974 56242 7026 56254
rect 8206 56306 8258 56318
rect 8206 56242 8258 56254
rect 9662 56306 9714 56318
rect 9662 56242 9714 56254
rect 11006 56306 11058 56318
rect 11006 56242 11058 56254
rect 12350 56306 12402 56318
rect 12350 56242 12402 56254
rect 13694 56306 13746 56318
rect 13694 56242 13746 56254
rect 14702 56306 14754 56318
rect 14702 56242 14754 56254
rect 15150 56306 15202 56318
rect 15150 56242 15202 56254
rect 15598 56306 15650 56318
rect 15598 56242 15650 56254
rect 15934 56306 15986 56318
rect 15934 56242 15986 56254
rect 18286 56306 18338 56318
rect 18286 56242 18338 56254
rect 24670 56306 24722 56318
rect 24670 56242 24722 56254
rect 27022 56306 27074 56318
rect 27022 56242 27074 56254
rect 28366 56306 28418 56318
rect 28366 56242 28418 56254
rect 28926 56306 28978 56318
rect 28926 56242 28978 56254
rect 29486 56306 29538 56318
rect 29486 56242 29538 56254
rect 31502 56306 31554 56318
rect 31502 56242 31554 56254
rect 35310 56306 35362 56318
rect 35310 56242 35362 56254
rect 39118 56306 39170 56318
rect 39118 56242 39170 56254
rect 43598 56306 43650 56318
rect 43598 56242 43650 56254
rect 44942 56306 44994 56318
rect 44942 56242 44994 56254
rect 45950 56306 46002 56318
rect 45950 56242 46002 56254
rect 47406 56306 47458 56318
rect 47406 56242 47458 56254
rect 48638 56306 48690 56318
rect 48638 56242 48690 56254
rect 49982 56306 50034 56318
rect 49982 56242 50034 56254
rect 51326 56306 51378 56318
rect 51326 56242 51378 56254
rect 52670 56306 52722 56318
rect 52670 56242 52722 56254
rect 54014 56306 54066 56318
rect 54014 56242 54066 56254
rect 55470 56306 55522 56318
rect 55470 56242 55522 56254
rect 5518 56194 5570 56206
rect 5518 56130 5570 56142
rect 5854 56194 5906 56206
rect 17278 56194 17330 56206
rect 16258 56142 16270 56194
rect 16322 56142 16334 56194
rect 5854 56130 5906 56142
rect 17278 56130 17330 56142
rect 17614 56194 17666 56206
rect 17614 56130 17666 56142
rect 18622 56194 18674 56206
rect 18622 56130 18674 56142
rect 18958 56194 19010 56206
rect 18958 56130 19010 56142
rect 19854 56194 19906 56206
rect 22082 56142 22094 56194
rect 22146 56142 22158 56194
rect 23650 56142 23662 56194
rect 23714 56142 23726 56194
rect 19854 56130 19906 56142
rect 27806 56082 27858 56094
rect 20066 56030 20078 56082
rect 20130 56030 20142 56082
rect 21186 56030 21198 56082
rect 21250 56030 21262 56082
rect 22754 56030 22766 56082
rect 22818 56030 22830 56082
rect 26114 56030 26126 56082
rect 26178 56030 26190 56082
rect 27806 56018 27858 56030
rect 30270 56082 30322 56094
rect 30270 56018 30322 56030
rect 32174 56082 32226 56094
rect 32174 56018 32226 56030
rect 33742 56082 33794 56094
rect 33742 56018 33794 56030
rect 35982 56082 36034 56094
rect 35982 56018 36034 56030
rect 37550 56082 37602 56094
rect 37550 56018 37602 56030
rect 39790 56082 39842 56094
rect 39790 56018 39842 56030
rect 42590 56082 42642 56094
rect 42590 56018 42642 56030
rect 6190 55970 6242 55982
rect 6190 55906 6242 55918
rect 7422 55970 7474 55982
rect 7422 55906 7474 55918
rect 8654 55970 8706 55982
rect 8654 55906 8706 55918
rect 10110 55970 10162 55982
rect 10110 55906 10162 55918
rect 11454 55970 11506 55982
rect 11454 55906 11506 55918
rect 13134 55970 13186 55982
rect 13134 55906 13186 55918
rect 14142 55970 14194 55982
rect 14142 55906 14194 55918
rect 19406 55970 19458 55982
rect 19406 55906 19458 55918
rect 20750 55970 20802 55982
rect 29934 55970 29986 55982
rect 42926 55970 42978 55982
rect 25554 55918 25566 55970
rect 25618 55918 25630 55970
rect 30706 55918 30718 55970
rect 30770 55918 30782 55970
rect 32610 55918 32622 55970
rect 32674 55918 32686 55970
rect 34178 55918 34190 55970
rect 34242 55918 34254 55970
rect 36418 55918 36430 55970
rect 36482 55918 36494 55970
rect 37986 55918 37998 55970
rect 38050 55918 38062 55970
rect 40450 55918 40462 55970
rect 40514 55918 40526 55970
rect 42018 55918 42030 55970
rect 42082 55918 42094 55970
rect 20750 55906 20802 55918
rect 29934 55906 29986 55918
rect 42926 55906 42978 55918
rect 44046 55970 44098 55982
rect 44046 55906 44098 55918
rect 44494 55970 44546 55982
rect 44494 55906 44546 55918
rect 46398 55970 46450 55982
rect 46398 55906 46450 55918
rect 47854 55970 47906 55982
rect 47854 55906 47906 55918
rect 49086 55970 49138 55982
rect 49086 55906 49138 55918
rect 50430 55970 50482 55982
rect 50430 55906 50482 55918
rect 51774 55970 51826 55982
rect 51774 55906 51826 55918
rect 53118 55970 53170 55982
rect 53118 55906 53170 55918
rect 55022 55970 55074 55982
rect 55022 55906 55074 55918
rect 55918 55970 55970 55982
rect 55918 55906 55970 55918
rect 45390 55858 45442 55870
rect 45390 55794 45442 55806
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 15486 55522 15538 55534
rect 15486 55458 15538 55470
rect 16158 55522 16210 55534
rect 16158 55458 16210 55470
rect 19182 55522 19234 55534
rect 19182 55458 19234 55470
rect 14814 55410 14866 55422
rect 4610 55358 4622 55410
rect 4674 55358 4686 55410
rect 5842 55358 5854 55410
rect 5906 55358 5918 55410
rect 14814 55346 14866 55358
rect 18510 55410 18562 55422
rect 18510 55346 18562 55358
rect 20078 55410 20130 55422
rect 22418 55358 22430 55410
rect 22482 55358 22494 55410
rect 28578 55358 28590 55410
rect 28642 55358 28654 55410
rect 32050 55358 32062 55410
rect 32114 55358 32126 55410
rect 35298 55358 35310 55410
rect 35362 55358 35374 55410
rect 37426 55358 37438 55410
rect 37490 55358 37502 55410
rect 39666 55358 39678 55410
rect 39730 55358 39742 55410
rect 20078 55346 20130 55358
rect 15262 55298 15314 55310
rect 1810 55246 1822 55298
rect 1874 55246 1886 55298
rect 8754 55246 8766 55298
rect 8818 55246 8830 55298
rect 15262 55234 15314 55246
rect 16494 55298 16546 55310
rect 16494 55234 16546 55246
rect 17166 55298 17218 55310
rect 17166 55234 17218 55246
rect 17390 55298 17442 55310
rect 17390 55234 17442 55246
rect 17838 55298 17890 55310
rect 25218 55246 25230 55298
rect 25282 55246 25294 55298
rect 25778 55246 25790 55298
rect 25842 55246 25854 55298
rect 29138 55246 29150 55298
rect 29202 55246 29214 55298
rect 32498 55246 32510 55298
rect 32562 55246 32574 55298
rect 38098 55246 38110 55298
rect 38162 55246 38174 55298
rect 39106 55246 39118 55298
rect 39170 55246 39182 55298
rect 42578 55246 42590 55298
rect 42642 55246 42654 55298
rect 17838 55234 17890 55246
rect 16606 55186 16658 55198
rect 2482 55134 2494 55186
rect 2546 55134 2558 55186
rect 7970 55134 7982 55186
rect 8034 55134 8046 55186
rect 16606 55122 16658 55134
rect 16830 55186 16882 55198
rect 16830 55122 16882 55134
rect 17950 55186 18002 55198
rect 17950 55122 18002 55134
rect 18286 55186 18338 55198
rect 18286 55122 18338 55134
rect 20414 55186 20466 55198
rect 20414 55122 20466 55134
rect 21646 55186 21698 55198
rect 21646 55122 21698 55134
rect 22094 55186 22146 55198
rect 35982 55186 36034 55198
rect 24546 55134 24558 55186
rect 24610 55134 24622 55186
rect 26450 55134 26462 55186
rect 26514 55134 26526 55186
rect 29922 55134 29934 55186
rect 29986 55134 29998 55186
rect 33170 55134 33182 55186
rect 33234 55134 33246 55186
rect 22094 55122 22146 55134
rect 35982 55122 36034 55134
rect 36318 55186 36370 55198
rect 36318 55122 36370 55134
rect 38558 55186 38610 55198
rect 42926 55186 42978 55198
rect 41794 55134 41806 55186
rect 41858 55134 41870 55186
rect 38558 55122 38610 55134
rect 42926 55122 42978 55134
rect 43038 55186 43090 55198
rect 43038 55122 43090 55134
rect 43374 55186 43426 55198
rect 43374 55122 43426 55134
rect 5070 55074 5122 55086
rect 5070 55010 5122 55022
rect 9214 55074 9266 55086
rect 9214 55010 9266 55022
rect 17054 55074 17106 55086
rect 35646 55074 35698 55086
rect 18834 55022 18846 55074
rect 18898 55022 18910 55074
rect 17054 55010 17106 55022
rect 35646 55010 35698 55022
rect 39342 55074 39394 55086
rect 39342 55010 39394 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 2494 54738 2546 54750
rect 19182 54738 19234 54750
rect 16818 54686 16830 54738
rect 16882 54686 16894 54738
rect 2494 54674 2546 54686
rect 19182 54674 19234 54686
rect 19294 54738 19346 54750
rect 19294 54674 19346 54686
rect 20190 54738 20242 54750
rect 20190 54674 20242 54686
rect 26238 54738 26290 54750
rect 26238 54674 26290 54686
rect 29262 54738 29314 54750
rect 29262 54674 29314 54686
rect 30046 54738 30098 54750
rect 30046 54674 30098 54686
rect 33070 54738 33122 54750
rect 33070 54674 33122 54686
rect 39678 54738 39730 54750
rect 39678 54674 39730 54686
rect 40238 54738 40290 54750
rect 40238 54674 40290 54686
rect 40910 54738 40962 54750
rect 40910 54674 40962 54686
rect 2382 54626 2434 54638
rect 2382 54562 2434 54574
rect 7534 54626 7586 54638
rect 7534 54562 7586 54574
rect 19742 54626 19794 54638
rect 19742 54562 19794 54574
rect 24446 54626 24498 54638
rect 35634 54574 35646 54626
rect 35698 54574 35710 54626
rect 24446 54562 24498 54574
rect 2606 54514 2658 54526
rect 2606 54450 2658 54462
rect 2942 54514 2994 54526
rect 4398 54514 4450 54526
rect 6974 54514 7026 54526
rect 3378 54462 3390 54514
rect 3442 54462 3454 54514
rect 6514 54462 6526 54514
rect 6578 54462 6590 54514
rect 2942 54450 2994 54462
rect 4398 54450 4450 54462
rect 6974 54450 7026 54462
rect 7310 54514 7362 54526
rect 7310 54450 7362 54462
rect 12126 54514 12178 54526
rect 16270 54514 16322 54526
rect 19070 54514 19122 54526
rect 24334 54514 24386 54526
rect 30382 54514 30434 54526
rect 12450 54462 12462 54514
rect 12514 54462 12526 54514
rect 17826 54462 17838 54514
rect 17890 54462 17902 54514
rect 18274 54462 18286 54514
rect 18338 54462 18350 54514
rect 18610 54462 18622 54514
rect 18674 54462 18686 54514
rect 19506 54462 19518 54514
rect 19570 54462 19582 54514
rect 23090 54462 23102 54514
rect 23154 54462 23166 54514
rect 23874 54462 23886 54514
rect 23938 54462 23950 54514
rect 28578 54462 28590 54514
rect 28642 54462 28654 54514
rect 12126 54450 12178 54462
rect 16270 54450 16322 54462
rect 19070 54450 19122 54462
rect 24334 54450 24386 54462
rect 30382 54450 30434 54462
rect 34526 54514 34578 54526
rect 39230 54514 39282 54526
rect 34850 54462 34862 54514
rect 34914 54462 34926 54514
rect 45490 54462 45502 54514
rect 45554 54462 45566 54514
rect 34526 54450 34578 54462
rect 39230 54450 39282 54462
rect 4958 54402 5010 54414
rect 15374 54402 15426 54414
rect 25342 54402 25394 54414
rect 3266 54350 3278 54402
rect 3330 54350 3342 54402
rect 6738 54350 6750 54402
rect 6802 54350 6814 54402
rect 7634 54350 7646 54402
rect 7698 54350 7710 54402
rect 13234 54350 13246 54402
rect 13298 54350 13310 54402
rect 20962 54350 20974 54402
rect 21026 54350 21038 54402
rect 4958 54338 5010 54350
rect 15374 54338 15426 54350
rect 25342 54338 25394 54350
rect 25790 54402 25842 54414
rect 25790 54338 25842 54350
rect 29710 54402 29762 54414
rect 29710 54338 29762 54350
rect 32062 54402 32114 54414
rect 32062 54338 32114 54350
rect 32510 54402 32562 54414
rect 37762 54350 37774 54402
rect 37826 54350 37838 54402
rect 42690 54350 42702 54402
rect 42754 54350 42766 54402
rect 44818 54350 44830 54402
rect 44882 54350 44894 54402
rect 32510 54338 32562 54350
rect 16494 54290 16546 54302
rect 16494 54226 16546 54238
rect 24222 54290 24274 54302
rect 24222 54226 24274 54238
rect 39118 54290 39170 54302
rect 39118 54226 39170 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 13470 53954 13522 53966
rect 13470 53890 13522 53902
rect 17166 53954 17218 53966
rect 17166 53890 17218 53902
rect 24558 53954 24610 53966
rect 24558 53890 24610 53902
rect 9550 53842 9602 53854
rect 13582 53842 13634 53854
rect 23774 53842 23826 53854
rect 34190 53842 34242 53854
rect 38558 53842 38610 53854
rect 4610 53790 4622 53842
rect 4674 53790 4686 53842
rect 12786 53790 12798 53842
rect 12850 53790 12862 53842
rect 17378 53790 17390 53842
rect 17442 53790 17454 53842
rect 20738 53790 20750 53842
rect 20802 53790 20814 53842
rect 33730 53790 33742 53842
rect 33794 53790 33806 53842
rect 35186 53790 35198 53842
rect 35250 53790 35262 53842
rect 9550 53778 9602 53790
rect 13582 53778 13634 53790
rect 23774 53778 23826 53790
rect 34190 53778 34242 53790
rect 38558 53778 38610 53790
rect 39566 53842 39618 53854
rect 45938 53790 45950 53842
rect 46002 53790 46014 53842
rect 51538 53790 51550 53842
rect 51602 53790 51614 53842
rect 39566 53778 39618 53790
rect 22206 53730 22258 53742
rect 38670 53730 38722 53742
rect 39118 53730 39170 53742
rect 1810 53678 1822 53730
rect 1874 53678 1886 53730
rect 9986 53678 9998 53730
rect 10050 53678 10062 53730
rect 10658 53678 10670 53730
rect 10722 53678 10734 53730
rect 17490 53678 17502 53730
rect 17554 53678 17566 53730
rect 17826 53678 17838 53730
rect 17890 53678 17902 53730
rect 22866 53678 22878 53730
rect 22930 53678 22942 53730
rect 24546 53678 24558 53730
rect 24610 53678 24622 53730
rect 30930 53678 30942 53730
rect 30994 53678 31006 53730
rect 38770 53678 38782 53730
rect 38834 53678 38846 53730
rect 22206 53666 22258 53678
rect 38670 53666 38722 53678
rect 39118 53666 39170 53678
rect 42254 53730 42306 53742
rect 42254 53666 42306 53678
rect 42814 53730 42866 53742
rect 48738 53678 48750 53730
rect 48802 53678 48814 53730
rect 42814 53666 42866 53678
rect 23326 53618 23378 53630
rect 2482 53566 2494 53618
rect 2546 53566 2558 53618
rect 18610 53566 18622 53618
rect 18674 53566 18686 53618
rect 23326 53554 23378 53566
rect 23550 53618 23602 53630
rect 23550 53554 23602 53566
rect 23886 53618 23938 53630
rect 23886 53554 23938 53566
rect 24222 53618 24274 53630
rect 35534 53618 35586 53630
rect 31602 53566 31614 53618
rect 31666 53566 31678 53618
rect 24222 53554 24274 53566
rect 35534 53554 35586 53566
rect 35870 53618 35922 53630
rect 35870 53554 35922 53566
rect 35982 53618 36034 53630
rect 35982 53554 36034 53566
rect 37774 53618 37826 53630
rect 37774 53554 37826 53566
rect 39454 53618 39506 53630
rect 39454 53554 39506 53566
rect 39678 53618 39730 53630
rect 39678 53554 39730 53566
rect 39790 53618 39842 53630
rect 43374 53618 43426 53630
rect 39890 53566 39902 53618
rect 39954 53566 39966 53618
rect 39790 53554 39842 53566
rect 43374 53554 43426 53566
rect 43710 53618 43762 53630
rect 43710 53554 43762 53566
rect 46286 53618 46338 53630
rect 49410 53566 49422 53618
rect 49474 53566 49486 53618
rect 46286 53554 46338 53566
rect 5070 53506 5122 53518
rect 5070 53442 5122 53454
rect 13694 53506 13746 53518
rect 13694 53442 13746 53454
rect 16830 53506 16882 53518
rect 16830 53442 16882 53454
rect 25006 53506 25058 53518
rect 25006 53442 25058 53454
rect 35310 53506 35362 53518
rect 35310 53442 35362 53454
rect 36206 53506 36258 53518
rect 36206 53442 36258 53454
rect 37886 53506 37938 53518
rect 37886 53442 37938 53454
rect 38110 53506 38162 53518
rect 38110 53442 38162 53454
rect 38446 53506 38498 53518
rect 38446 53442 38498 53454
rect 46062 53506 46114 53518
rect 46062 53442 46114 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 2718 53170 2770 53182
rect 2718 53106 2770 53118
rect 3502 53170 3554 53182
rect 3502 53106 3554 53118
rect 18846 53170 18898 53182
rect 18846 53106 18898 53118
rect 19406 53170 19458 53182
rect 19406 53106 19458 53118
rect 23886 53170 23938 53182
rect 23886 53106 23938 53118
rect 24670 53170 24722 53182
rect 24670 53106 24722 53118
rect 30830 53170 30882 53182
rect 30830 53106 30882 53118
rect 31950 53170 32002 53182
rect 31950 53106 32002 53118
rect 33966 53170 34018 53182
rect 33966 53106 34018 53118
rect 34078 53170 34130 53182
rect 34078 53106 34130 53118
rect 34302 53170 34354 53182
rect 34302 53106 34354 53118
rect 34750 53170 34802 53182
rect 34750 53106 34802 53118
rect 36878 53170 36930 53182
rect 36878 53106 36930 53118
rect 39454 53170 39506 53182
rect 39454 53106 39506 53118
rect 41022 53170 41074 53182
rect 41022 53106 41074 53118
rect 42142 53170 42194 53182
rect 42142 53106 42194 53118
rect 42590 53170 42642 53182
rect 42590 53106 42642 53118
rect 49086 53170 49138 53182
rect 49086 53106 49138 53118
rect 4398 53058 4450 53070
rect 4398 52994 4450 53006
rect 8094 53058 8146 53070
rect 8094 52994 8146 53006
rect 12910 53058 12962 53070
rect 12910 52994 12962 53006
rect 18174 53058 18226 53070
rect 18174 52994 18226 53006
rect 25454 53058 25506 53070
rect 25454 52994 25506 53006
rect 26014 53058 26066 53070
rect 40238 53058 40290 53070
rect 28242 53006 28254 53058
rect 28306 53006 28318 53058
rect 38882 53006 38894 53058
rect 38946 53006 38958 53058
rect 26014 52994 26066 53006
rect 40238 52994 40290 53006
rect 41806 53058 41858 53070
rect 41806 52994 41858 53006
rect 43038 53058 43090 53070
rect 45714 53006 45726 53058
rect 45778 53006 45790 53058
rect 43038 52994 43090 53006
rect 3278 52946 3330 52958
rect 2930 52894 2942 52946
rect 2994 52894 3006 52946
rect 3278 52882 3330 52894
rect 3614 52946 3666 52958
rect 3614 52882 3666 52894
rect 3838 52946 3890 52958
rect 3838 52882 3890 52894
rect 4286 52946 4338 52958
rect 4286 52882 4338 52894
rect 4510 52946 4562 52958
rect 4510 52882 4562 52894
rect 11454 52946 11506 52958
rect 13470 52946 13522 52958
rect 12450 52894 12462 52946
rect 12514 52894 12526 52946
rect 11454 52882 11506 52894
rect 13470 52882 13522 52894
rect 13806 52946 13858 52958
rect 13806 52882 13858 52894
rect 14030 52946 14082 52958
rect 14030 52882 14082 52894
rect 18510 52946 18562 52958
rect 18510 52882 18562 52894
rect 19182 52946 19234 52958
rect 19182 52882 19234 52894
rect 19854 52946 19906 52958
rect 23774 52946 23826 52958
rect 20066 52894 20078 52946
rect 20130 52894 20142 52946
rect 23538 52894 23550 52946
rect 23602 52894 23614 52946
rect 19854 52882 19906 52894
rect 23774 52882 23826 52894
rect 23998 52946 24050 52958
rect 32286 52946 32338 52958
rect 35198 52946 35250 52958
rect 24210 52894 24222 52946
rect 24274 52894 24286 52946
rect 27570 52894 27582 52946
rect 27634 52894 27646 52946
rect 34514 52894 34526 52946
rect 34578 52894 34590 52946
rect 23998 52882 24050 52894
rect 32286 52882 32338 52894
rect 35198 52882 35250 52894
rect 35646 52946 35698 52958
rect 35646 52882 35698 52894
rect 36206 52946 36258 52958
rect 36206 52882 36258 52894
rect 37214 52946 37266 52958
rect 37214 52882 37266 52894
rect 38110 52946 38162 52958
rect 38110 52882 38162 52894
rect 38670 52946 38722 52958
rect 41134 52946 41186 52958
rect 38994 52894 39006 52946
rect 39058 52894 39070 52946
rect 38670 52882 38722 52894
rect 41134 52882 41186 52894
rect 42478 52946 42530 52958
rect 43934 52946 43986 52958
rect 43474 52894 43486 52946
rect 43538 52894 43550 52946
rect 45042 52894 45054 52946
rect 45106 52894 45118 52946
rect 48850 52894 48862 52946
rect 48914 52894 48926 52946
rect 49970 52894 49982 52946
rect 50034 52894 50046 52946
rect 42478 52882 42530 52894
rect 43934 52882 43986 52894
rect 10334 52834 10386 52846
rect 13582 52834 13634 52846
rect 10882 52782 10894 52834
rect 10946 52782 10958 52834
rect 12002 52782 12014 52834
rect 12066 52782 12078 52834
rect 10334 52770 10386 52782
rect 13582 52770 13634 52782
rect 16606 52834 16658 52846
rect 16606 52770 16658 52782
rect 17726 52834 17778 52846
rect 17726 52770 17778 52782
rect 18734 52834 18786 52846
rect 18734 52770 18786 52782
rect 19294 52834 19346 52846
rect 35982 52834 36034 52846
rect 20850 52782 20862 52834
rect 20914 52782 20926 52834
rect 22978 52782 22990 52834
rect 23042 52782 23054 52834
rect 30370 52782 30382 52834
rect 30434 52782 30446 52834
rect 19294 52770 19346 52782
rect 35982 52770 36034 52782
rect 38446 52834 38498 52846
rect 38446 52770 38498 52782
rect 39678 52834 39730 52846
rect 49198 52834 49250 52846
rect 47842 52782 47854 52834
rect 47906 52782 47918 52834
rect 39678 52770 39730 52782
rect 49198 52770 49250 52782
rect 49534 52834 49586 52846
rect 49858 52782 49870 52834
rect 49922 52782 49934 52834
rect 49534 52770 49586 52782
rect 2606 52722 2658 52734
rect 10558 52722 10610 52734
rect 4946 52670 4958 52722
rect 5010 52670 5022 52722
rect 2606 52658 2658 52670
rect 10558 52658 10610 52670
rect 11566 52722 11618 52734
rect 11566 52658 11618 52670
rect 16494 52722 16546 52734
rect 16494 52658 16546 52670
rect 17950 52722 18002 52734
rect 17950 52658 18002 52670
rect 25230 52722 25282 52734
rect 25230 52658 25282 52670
rect 25566 52722 25618 52734
rect 25566 52658 25618 52670
rect 35422 52722 35474 52734
rect 35422 52658 35474 52670
rect 36430 52722 36482 52734
rect 36430 52658 36482 52670
rect 37662 52722 37714 52734
rect 37662 52658 37714 52670
rect 37886 52722 37938 52734
rect 37886 52658 37938 52670
rect 40014 52722 40066 52734
rect 40014 52658 40066 52670
rect 41022 52722 41074 52734
rect 41022 52658 41074 52670
rect 42590 52722 42642 52734
rect 42590 52658 42642 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 4398 52386 4450 52398
rect 4398 52322 4450 52334
rect 20638 52386 20690 52398
rect 20638 52322 20690 52334
rect 37998 52386 38050 52398
rect 37998 52322 38050 52334
rect 39342 52386 39394 52398
rect 39342 52322 39394 52334
rect 40798 52386 40850 52398
rect 40798 52322 40850 52334
rect 41246 52386 41298 52398
rect 41246 52322 41298 52334
rect 49870 52386 49922 52398
rect 50530 52334 50542 52386
rect 50594 52334 50606 52386
rect 49870 52322 49922 52334
rect 7982 52274 8034 52286
rect 20190 52274 20242 52286
rect 33742 52274 33794 52286
rect 11330 52222 11342 52274
rect 11394 52222 11406 52274
rect 18274 52222 18286 52274
rect 18338 52222 18350 52274
rect 24546 52222 24558 52274
rect 24610 52222 24622 52274
rect 24994 52222 25006 52274
rect 25058 52222 25070 52274
rect 27122 52222 27134 52274
rect 27186 52222 27198 52274
rect 33282 52222 33294 52274
rect 33346 52222 33358 52274
rect 7982 52210 8034 52222
rect 20190 52210 20242 52222
rect 33742 52210 33794 52222
rect 36094 52274 36146 52286
rect 41806 52274 41858 52286
rect 38434 52222 38446 52274
rect 38498 52222 38510 52274
rect 36094 52210 36146 52222
rect 41806 52210 41858 52222
rect 46174 52274 46226 52286
rect 46174 52210 46226 52222
rect 49422 52274 49474 52286
rect 49422 52210 49474 52222
rect 4622 52162 4674 52174
rect 4162 52110 4174 52162
rect 4226 52110 4238 52162
rect 4622 52098 4674 52110
rect 6302 52162 6354 52174
rect 6302 52098 6354 52110
rect 6414 52162 6466 52174
rect 6862 52162 6914 52174
rect 6626 52110 6638 52162
rect 6690 52110 6702 52162
rect 6414 52098 6466 52110
rect 6862 52098 6914 52110
rect 7198 52162 7250 52174
rect 12574 52162 12626 52174
rect 12910 52162 12962 52174
rect 8530 52110 8542 52162
rect 8594 52110 8606 52162
rect 12786 52110 12798 52162
rect 12850 52110 12862 52162
rect 7198 52098 7250 52110
rect 12574 52098 12626 52110
rect 12910 52098 12962 52110
rect 13694 52162 13746 52174
rect 13694 52098 13746 52110
rect 13806 52162 13858 52174
rect 13806 52098 13858 52110
rect 13918 52162 13970 52174
rect 18734 52162 18786 52174
rect 14802 52110 14814 52162
rect 14866 52110 14878 52162
rect 15474 52110 15486 52162
rect 15538 52110 15550 52162
rect 13918 52098 13970 52110
rect 18734 52098 18786 52110
rect 19182 52162 19234 52174
rect 19182 52098 19234 52110
rect 19742 52162 19794 52174
rect 19742 52098 19794 52110
rect 20750 52162 20802 52174
rect 20750 52098 20802 52110
rect 23102 52162 23154 52174
rect 24446 52162 24498 52174
rect 39454 52162 39506 52174
rect 23538 52110 23550 52162
rect 23602 52110 23614 52162
rect 27906 52110 27918 52162
rect 27970 52110 27982 52162
rect 30482 52110 30494 52162
rect 30546 52110 30558 52162
rect 31154 52110 31166 52162
rect 31218 52110 31230 52162
rect 23102 52098 23154 52110
rect 24446 52098 24498 52110
rect 39454 52098 39506 52110
rect 40126 52162 40178 52174
rect 40126 52098 40178 52110
rect 40910 52162 40962 52174
rect 42030 52162 42082 52174
rect 41234 52110 41246 52162
rect 41298 52110 41310 52162
rect 40910 52098 40962 52110
rect 42030 52098 42082 52110
rect 47406 52162 47458 52174
rect 47406 52098 47458 52110
rect 47854 52162 47906 52174
rect 50766 52162 50818 52174
rect 50530 52110 50542 52162
rect 50594 52110 50606 52162
rect 51874 52110 51886 52162
rect 51938 52110 51950 52162
rect 47854 52098 47906 52110
rect 50766 52098 50818 52110
rect 7534 52050 7586 52062
rect 20638 52050 20690 52062
rect 9202 51998 9214 52050
rect 9266 51998 9278 52050
rect 16146 51998 16158 52050
rect 16210 51998 16222 52050
rect 7534 51986 7586 51998
rect 20638 51986 20690 51998
rect 23998 52050 24050 52062
rect 23998 51986 24050 51998
rect 35758 52050 35810 52062
rect 35758 51986 35810 51998
rect 36206 52050 36258 52062
rect 36206 51986 36258 51998
rect 38110 52050 38162 52062
rect 38110 51986 38162 51998
rect 38558 52050 38610 52062
rect 41582 52050 41634 52062
rect 49758 52050 49810 52062
rect 38770 51998 38782 52050
rect 38834 51998 38846 52050
rect 39778 51998 39790 52050
rect 39842 51998 39854 52050
rect 42130 51998 42142 52050
rect 42194 51998 42206 52050
rect 42690 51998 42702 52050
rect 42754 51998 42766 52050
rect 38558 51986 38610 51998
rect 41582 51986 41634 51998
rect 49758 51986 49810 51998
rect 51102 52050 51154 52062
rect 51102 51986 51154 51998
rect 51438 52050 51490 52062
rect 51438 51986 51490 51998
rect 4286 51938 4338 51950
rect 7086 51938 7138 51950
rect 24222 51938 24274 51950
rect 5842 51886 5854 51938
rect 5906 51886 5918 51938
rect 14354 51886 14366 51938
rect 14418 51886 14430 51938
rect 15026 51886 15038 51938
rect 15090 51886 15102 51938
rect 4286 51874 4338 51886
rect 7086 51874 7138 51886
rect 24222 51874 24274 51886
rect 24558 51938 24610 51950
rect 24558 51874 24610 51886
rect 28366 51938 28418 51950
rect 28366 51874 28418 51886
rect 35982 51938 36034 51950
rect 35982 51874 36034 51886
rect 37998 51938 38050 51950
rect 37998 51874 38050 51886
rect 39006 51938 39058 51950
rect 39006 51874 39058 51886
rect 40798 51938 40850 51950
rect 40798 51874 40850 51886
rect 46734 51938 46786 51950
rect 47742 51938 47794 51950
rect 47058 51886 47070 51938
rect 47122 51886 47134 51938
rect 46734 51874 46786 51886
rect 47742 51874 47794 51886
rect 49310 51938 49362 51950
rect 49310 51874 49362 51886
rect 49870 51938 49922 51950
rect 49870 51874 49922 51886
rect 50990 51938 51042 51950
rect 50990 51874 51042 51886
rect 51326 51938 51378 51950
rect 51326 51874 51378 51886
rect 51662 51938 51714 51950
rect 51662 51874 51714 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 16270 51602 16322 51614
rect 16270 51538 16322 51550
rect 22206 51602 22258 51614
rect 22206 51538 22258 51550
rect 22318 51602 22370 51614
rect 22318 51538 22370 51550
rect 23662 51602 23714 51614
rect 23662 51538 23714 51550
rect 31838 51602 31890 51614
rect 31838 51538 31890 51550
rect 33854 51602 33906 51614
rect 33854 51538 33906 51550
rect 34862 51602 34914 51614
rect 34862 51538 34914 51550
rect 35198 51602 35250 51614
rect 35198 51538 35250 51550
rect 35982 51602 36034 51614
rect 35982 51538 36034 51550
rect 38558 51602 38610 51614
rect 38558 51538 38610 51550
rect 49086 51602 49138 51614
rect 49086 51538 49138 51550
rect 7198 51490 7250 51502
rect 4610 51438 4622 51490
rect 4674 51438 4686 51490
rect 7198 51426 7250 51438
rect 11678 51490 11730 51502
rect 11678 51426 11730 51438
rect 12798 51490 12850 51502
rect 12798 51426 12850 51438
rect 13134 51490 13186 51502
rect 13134 51426 13186 51438
rect 13470 51490 13522 51502
rect 13470 51426 13522 51438
rect 15374 51490 15426 51502
rect 15374 51426 15426 51438
rect 15822 51490 15874 51502
rect 15822 51426 15874 51438
rect 17390 51490 17442 51502
rect 17390 51426 17442 51438
rect 18286 51490 18338 51502
rect 18286 51426 18338 51438
rect 19070 51490 19122 51502
rect 34190 51490 34242 51502
rect 23090 51438 23102 51490
rect 23154 51438 23166 51490
rect 19070 51426 19122 51438
rect 34190 51426 34242 51438
rect 35422 51490 35474 51502
rect 35422 51426 35474 51438
rect 37214 51490 37266 51502
rect 37214 51426 37266 51438
rect 38446 51490 38498 51502
rect 38446 51426 38498 51438
rect 38670 51490 38722 51502
rect 40014 51490 40066 51502
rect 38670 51426 38722 51438
rect 38782 51434 38834 51446
rect 6190 51378 6242 51390
rect 10558 51378 10610 51390
rect 6738 51326 6750 51378
rect 6802 51326 6814 51378
rect 6190 51314 6242 51326
rect 10558 51314 10610 51326
rect 11006 51378 11058 51390
rect 12126 51378 12178 51390
rect 11330 51326 11342 51378
rect 11394 51326 11406 51378
rect 11006 51314 11058 51326
rect 12126 51314 12178 51326
rect 13806 51378 13858 51390
rect 14478 51378 14530 51390
rect 14018 51326 14030 51378
rect 14082 51326 14094 51378
rect 13806 51314 13858 51326
rect 14478 51314 14530 51326
rect 15262 51378 15314 51390
rect 15262 51314 15314 51326
rect 15598 51378 15650 51390
rect 15598 51314 15650 51326
rect 16382 51378 16434 51390
rect 16382 51314 16434 51326
rect 16830 51378 16882 51390
rect 19854 51378 19906 51390
rect 18498 51326 18510 51378
rect 18562 51326 18574 51378
rect 16830 51314 16882 51326
rect 19854 51314 19906 51326
rect 20190 51378 20242 51390
rect 20190 51314 20242 51326
rect 20526 51378 20578 51390
rect 33966 51378 34018 51390
rect 22866 51326 22878 51378
rect 22930 51326 22942 51378
rect 28130 51326 28142 51378
rect 28194 51326 28206 51378
rect 28578 51326 28590 51378
rect 28642 51326 28654 51378
rect 20526 51314 20578 51326
rect 33966 51314 34018 51326
rect 34414 51378 34466 51390
rect 34414 51314 34466 51326
rect 34638 51378 34690 51390
rect 34638 51314 34690 51326
rect 34974 51378 35026 51390
rect 34974 51314 35026 51326
rect 35646 51378 35698 51390
rect 36654 51378 36706 51390
rect 40014 51426 40066 51438
rect 42030 51490 42082 51502
rect 43710 51490 43762 51502
rect 42690 51438 42702 51490
rect 42754 51438 42766 51490
rect 42914 51438 42926 51490
rect 42978 51438 42990 51490
rect 42030 51426 42082 51438
rect 43710 51426 43762 51438
rect 47630 51490 47682 51502
rect 47630 51426 47682 51438
rect 49422 51490 49474 51502
rect 52434 51438 52446 51490
rect 52498 51438 52510 51490
rect 49422 51426 49474 51438
rect 36194 51326 36206 51378
rect 36258 51326 36270 51378
rect 36418 51326 36430 51378
rect 36482 51326 36494 51378
rect 36978 51326 36990 51378
rect 37042 51326 37054 51378
rect 38782 51370 38834 51382
rect 39454 51378 39506 51390
rect 41470 51378 41522 51390
rect 39218 51326 39230 51378
rect 39282 51326 39294 51378
rect 39778 51326 39790 51378
rect 39842 51326 39854 51378
rect 35646 51314 35698 51326
rect 36654 51314 36706 51326
rect 39454 51314 39506 51326
rect 41470 51314 41522 51326
rect 42254 51378 42306 51390
rect 42254 51314 42306 51326
rect 43598 51378 43650 51390
rect 43598 51314 43650 51326
rect 46398 51378 46450 51390
rect 46398 51314 46450 51326
rect 46846 51378 46898 51390
rect 46846 51314 46898 51326
rect 47070 51378 47122 51390
rect 47070 51314 47122 51326
rect 47518 51378 47570 51390
rect 49758 51378 49810 51390
rect 48850 51326 48862 51378
rect 48914 51326 48926 51378
rect 47518 51314 47570 51326
rect 49758 51314 49810 51326
rect 49982 51378 50034 51390
rect 50754 51326 50766 51378
rect 50818 51326 50830 51378
rect 51650 51326 51662 51378
rect 51714 51326 51726 51378
rect 49982 51314 50034 51326
rect 16046 51266 16098 51278
rect 6066 51214 6078 51266
rect 6130 51214 6142 51266
rect 16046 51202 16098 51214
rect 17614 51266 17666 51278
rect 17614 51202 17666 51214
rect 20078 51266 20130 51278
rect 20078 51202 20130 51214
rect 22094 51266 22146 51278
rect 36878 51266 36930 51278
rect 23762 51214 23774 51266
rect 23826 51214 23838 51266
rect 25218 51214 25230 51266
rect 25282 51214 25294 51266
rect 27346 51214 27358 51266
rect 27410 51214 27422 51266
rect 29250 51214 29262 51266
rect 29314 51214 29326 51266
rect 31378 51214 31390 51266
rect 31442 51214 31454 51266
rect 22094 51202 22146 51214
rect 36878 51202 36930 51214
rect 39678 51266 39730 51278
rect 39678 51202 39730 51214
rect 41246 51266 41298 51278
rect 41246 51202 41298 51214
rect 45614 51266 45666 51278
rect 45614 51202 45666 51214
rect 46622 51266 46674 51278
rect 46622 51202 46674 51214
rect 49870 51266 49922 51278
rect 51326 51266 51378 51278
rect 50978 51214 50990 51266
rect 51042 51214 51054 51266
rect 54562 51214 54574 51266
rect 54626 51214 54638 51266
rect 49870 51202 49922 51214
rect 51326 51202 51378 51214
rect 10110 51154 10162 51166
rect 10110 51090 10162 51102
rect 10222 51154 10274 51166
rect 10222 51090 10274 51102
rect 10446 51154 10498 51166
rect 10446 51090 10498 51102
rect 11342 51154 11394 51166
rect 11342 51090 11394 51102
rect 11790 51154 11842 51166
rect 11790 51090 11842 51102
rect 12014 51154 12066 51166
rect 12014 51090 12066 51102
rect 13582 51154 13634 51166
rect 13582 51090 13634 51102
rect 14366 51154 14418 51166
rect 14366 51090 14418 51102
rect 16270 51154 16322 51166
rect 16270 51090 16322 51102
rect 17950 51154 18002 51166
rect 17950 51090 18002 51102
rect 18958 51154 19010 51166
rect 18958 51090 19010 51102
rect 23438 51154 23490 51166
rect 23438 51090 23490 51102
rect 35870 51154 35922 51166
rect 43710 51154 43762 51166
rect 41794 51102 41806 51154
rect 41858 51102 41870 51154
rect 35870 51090 35922 51102
rect 43710 51090 43762 51102
rect 45838 51154 45890 51166
rect 47630 51154 47682 51166
rect 46162 51102 46174 51154
rect 46226 51102 46238 51154
rect 45838 51090 45890 51102
rect 47630 51090 47682 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 34638 50818 34690 50830
rect 34638 50754 34690 50766
rect 34974 50818 35026 50830
rect 34974 50754 35026 50766
rect 36206 50818 36258 50830
rect 36206 50754 36258 50766
rect 42702 50818 42754 50830
rect 42702 50754 42754 50766
rect 43038 50818 43090 50830
rect 43038 50754 43090 50766
rect 45054 50818 45106 50830
rect 45054 50754 45106 50766
rect 45390 50818 45442 50830
rect 45390 50754 45442 50766
rect 49870 50818 49922 50830
rect 51090 50766 51102 50818
rect 51154 50766 51166 50818
rect 49870 50754 49922 50766
rect 6638 50706 6690 50718
rect 24334 50706 24386 50718
rect 2482 50654 2494 50706
rect 2546 50654 2558 50706
rect 4610 50654 4622 50706
rect 4674 50654 4686 50706
rect 8754 50654 8766 50706
rect 8818 50654 8830 50706
rect 10882 50654 10894 50706
rect 10946 50654 10958 50706
rect 14690 50654 14702 50706
rect 14754 50654 14766 50706
rect 6638 50642 6690 50654
rect 24334 50642 24386 50654
rect 25006 50706 25058 50718
rect 25006 50642 25058 50654
rect 28366 50706 28418 50718
rect 48190 50706 48242 50718
rect 39218 50654 39230 50706
rect 39282 50654 39294 50706
rect 42242 50654 42254 50706
rect 42306 50654 42318 50706
rect 47058 50654 47070 50706
rect 47122 50654 47134 50706
rect 50194 50654 50206 50706
rect 50258 50654 50270 50706
rect 55570 50654 55582 50706
rect 55634 50654 55646 50706
rect 28366 50642 28418 50654
rect 48190 50642 48242 50654
rect 5966 50594 6018 50606
rect 1810 50542 1822 50594
rect 1874 50542 1886 50594
rect 5966 50530 6018 50542
rect 6190 50594 6242 50606
rect 6190 50530 6242 50542
rect 6862 50594 6914 50606
rect 11230 50594 11282 50606
rect 7074 50542 7086 50594
rect 7138 50542 7150 50594
rect 8082 50542 8094 50594
rect 8146 50542 8158 50594
rect 6862 50530 6914 50542
rect 11230 50530 11282 50542
rect 12574 50594 12626 50606
rect 19070 50594 19122 50606
rect 15026 50542 15038 50594
rect 15090 50542 15102 50594
rect 15362 50542 15374 50594
rect 15426 50542 15438 50594
rect 18386 50542 18398 50594
rect 18450 50542 18462 50594
rect 12574 50530 12626 50542
rect 19070 50530 19122 50542
rect 19406 50594 19458 50606
rect 19406 50530 19458 50542
rect 19742 50594 19794 50606
rect 19742 50530 19794 50542
rect 20190 50594 20242 50606
rect 20190 50530 20242 50542
rect 20414 50594 20466 50606
rect 20414 50530 20466 50542
rect 23550 50594 23602 50606
rect 23550 50530 23602 50542
rect 24110 50594 24162 50606
rect 24110 50530 24162 50542
rect 35422 50594 35474 50606
rect 35422 50530 35474 50542
rect 35646 50594 35698 50606
rect 35646 50530 35698 50542
rect 35982 50594 36034 50606
rect 35982 50530 36034 50542
rect 36990 50594 37042 50606
rect 39902 50594 39954 50606
rect 37650 50542 37662 50594
rect 37714 50542 37726 50594
rect 38210 50542 38222 50594
rect 38274 50542 38286 50594
rect 39106 50542 39118 50594
rect 39170 50542 39182 50594
rect 36990 50530 37042 50542
rect 39902 50530 39954 50542
rect 41694 50594 41746 50606
rect 48078 50594 48130 50606
rect 42354 50542 42366 50594
rect 42418 50542 42430 50594
rect 43586 50542 43598 50594
rect 43650 50542 43662 50594
rect 46050 50542 46062 50594
rect 46114 50542 46126 50594
rect 46610 50542 46622 50594
rect 46674 50542 46686 50594
rect 47506 50542 47518 50594
rect 47570 50542 47582 50594
rect 41694 50530 41746 50542
rect 48078 50530 48130 50542
rect 48302 50594 48354 50606
rect 48302 50530 48354 50542
rect 49310 50594 49362 50606
rect 49310 50530 49362 50542
rect 49646 50594 49698 50606
rect 49646 50530 49698 50542
rect 50542 50594 50594 50606
rect 50542 50530 50594 50542
rect 50878 50594 50930 50606
rect 51202 50542 51214 50594
rect 51266 50542 51278 50594
rect 52658 50542 52670 50594
rect 52722 50542 52734 50594
rect 50878 50530 50930 50542
rect 6526 50482 6578 50494
rect 6526 50418 6578 50430
rect 7534 50482 7586 50494
rect 7534 50418 7586 50430
rect 11790 50482 11842 50494
rect 11790 50418 11842 50430
rect 12350 50482 12402 50494
rect 19182 50482 19234 50494
rect 14914 50430 14926 50482
rect 14978 50430 14990 50482
rect 15810 50430 15822 50482
rect 15874 50430 15886 50482
rect 18498 50430 18510 50482
rect 18562 50430 18574 50482
rect 18722 50430 18734 50482
rect 18786 50430 18798 50482
rect 12350 50418 12402 50430
rect 19182 50418 19234 50430
rect 19966 50482 20018 50494
rect 19966 50418 20018 50430
rect 22542 50482 22594 50494
rect 22542 50418 22594 50430
rect 22878 50482 22930 50494
rect 24558 50482 24610 50494
rect 23874 50430 23886 50482
rect 23938 50430 23950 50482
rect 22878 50418 22930 50430
rect 24558 50418 24610 50430
rect 24894 50482 24946 50494
rect 24894 50418 24946 50430
rect 25454 50482 25506 50494
rect 25454 50418 25506 50430
rect 30718 50482 30770 50494
rect 30718 50418 30770 50430
rect 34750 50482 34802 50494
rect 34750 50418 34802 50430
rect 37102 50482 37154 50494
rect 39342 50482 39394 50494
rect 42030 50482 42082 50494
rect 38322 50430 38334 50482
rect 38386 50430 38398 50482
rect 38994 50430 39006 50482
rect 39058 50430 39070 50482
rect 40114 50430 40126 50482
rect 40178 50430 40190 50482
rect 40674 50430 40686 50482
rect 40738 50430 40750 50482
rect 37102 50418 37154 50430
rect 39342 50418 39394 50430
rect 42030 50418 42082 50430
rect 42926 50482 42978 50494
rect 48526 50482 48578 50494
rect 43362 50430 43374 50482
rect 43426 50430 43438 50482
rect 46162 50430 46174 50482
rect 46226 50430 46238 50482
rect 47282 50430 47294 50482
rect 47346 50430 47358 50482
rect 42926 50418 42978 50430
rect 48526 50418 48578 50430
rect 49422 50482 49474 50494
rect 49422 50418 49474 50430
rect 50094 50482 50146 50494
rect 53442 50430 53454 50482
rect 53506 50430 53518 50482
rect 50094 50418 50146 50430
rect 5070 50370 5122 50382
rect 7422 50370 7474 50382
rect 24446 50370 24498 50382
rect 5618 50318 5630 50370
rect 5682 50318 5694 50370
rect 12898 50318 12910 50370
rect 12962 50318 12974 50370
rect 5070 50306 5122 50318
rect 7422 50306 7474 50318
rect 24446 50306 24498 50318
rect 35310 50370 35362 50382
rect 35310 50306 35362 50318
rect 39566 50370 39618 50382
rect 51326 50370 51378 50382
rect 40002 50318 40014 50370
rect 40066 50318 40078 50370
rect 41346 50318 41358 50370
rect 41410 50318 41422 50370
rect 39566 50306 39618 50318
rect 51326 50306 51378 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 12350 50034 12402 50046
rect 10546 49982 10558 50034
rect 10610 49982 10622 50034
rect 12350 49970 12402 49982
rect 16158 50034 16210 50046
rect 16158 49970 16210 49982
rect 17838 50034 17890 50046
rect 21982 50034 22034 50046
rect 24222 50034 24274 50046
rect 18946 49982 18958 50034
rect 19010 49982 19022 50034
rect 22978 49982 22990 50034
rect 23042 49982 23054 50034
rect 17838 49970 17890 49982
rect 21982 49970 22034 49982
rect 24222 49970 24274 49982
rect 34302 50034 34354 50046
rect 34302 49970 34354 49982
rect 35086 50034 35138 50046
rect 39790 50034 39842 50046
rect 41918 50034 41970 50046
rect 37538 49982 37550 50034
rect 37602 49982 37614 50034
rect 40898 49982 40910 50034
rect 40962 49982 40974 50034
rect 43586 49982 43598 50034
rect 43650 49982 43662 50034
rect 35086 49970 35138 49982
rect 39790 49970 39842 49982
rect 41918 49970 41970 49982
rect 12238 49922 12290 49934
rect 6178 49870 6190 49922
rect 6242 49870 6254 49922
rect 12238 49858 12290 49870
rect 15934 49922 15986 49934
rect 15934 49858 15986 49870
rect 18398 49922 18450 49934
rect 18398 49858 18450 49870
rect 31502 49922 31554 49934
rect 31502 49858 31554 49870
rect 31838 49922 31890 49934
rect 31838 49858 31890 49870
rect 32174 49922 32226 49934
rect 43038 49922 43090 49934
rect 36642 49870 36654 49922
rect 36706 49870 36718 49922
rect 39106 49870 39118 49922
rect 39170 49870 39182 49922
rect 32174 49858 32226 49870
rect 43038 49858 43090 49870
rect 43262 49922 43314 49934
rect 43262 49858 43314 49870
rect 48750 49922 48802 49934
rect 48750 49858 48802 49870
rect 9998 49810 10050 49822
rect 1810 49758 1822 49810
rect 1874 49758 1886 49810
rect 5394 49758 5406 49810
rect 5458 49758 5470 49810
rect 9998 49746 10050 49758
rect 11006 49810 11058 49822
rect 12574 49810 12626 49822
rect 11218 49758 11230 49810
rect 11282 49758 11294 49810
rect 11006 49746 11058 49758
rect 12574 49746 12626 49758
rect 13246 49810 13298 49822
rect 14142 49810 14194 49822
rect 13458 49758 13470 49810
rect 13522 49758 13534 49810
rect 13246 49746 13298 49758
rect 14142 49746 14194 49758
rect 14366 49810 14418 49822
rect 14366 49746 14418 49758
rect 15038 49810 15090 49822
rect 17278 49810 17330 49822
rect 18622 49810 18674 49822
rect 16370 49758 16382 49810
rect 16434 49758 16446 49810
rect 17602 49758 17614 49810
rect 17666 49758 17678 49810
rect 15038 49746 15090 49758
rect 17278 49746 17330 49758
rect 18622 49746 18674 49758
rect 19518 49810 19570 49822
rect 19518 49746 19570 49758
rect 19742 49810 19794 49822
rect 19742 49746 19794 49758
rect 20078 49810 20130 49822
rect 20078 49746 20130 49758
rect 20526 49810 20578 49822
rect 20526 49746 20578 49758
rect 21086 49810 21138 49822
rect 22542 49810 22594 49822
rect 22194 49758 22206 49810
rect 22258 49758 22270 49810
rect 21086 49746 21138 49758
rect 22542 49746 22594 49758
rect 22878 49810 22930 49822
rect 23662 49810 23714 49822
rect 23090 49758 23102 49810
rect 23154 49758 23166 49810
rect 22878 49746 22930 49758
rect 23662 49746 23714 49758
rect 24110 49810 24162 49822
rect 24110 49746 24162 49758
rect 24334 49810 24386 49822
rect 34190 49810 34242 49822
rect 27682 49758 27694 49810
rect 27746 49758 27758 49810
rect 24334 49746 24386 49758
rect 34190 49746 34242 49758
rect 34526 49810 34578 49822
rect 36878 49810 36930 49822
rect 41246 49810 41298 49822
rect 43934 49810 43986 49822
rect 34850 49758 34862 49810
rect 34914 49758 34926 49810
rect 35522 49758 35534 49810
rect 35586 49758 35598 49810
rect 36194 49758 36206 49810
rect 36258 49758 36270 49810
rect 37314 49758 37326 49810
rect 37378 49758 37390 49810
rect 37874 49758 37886 49810
rect 37938 49758 37950 49810
rect 38658 49758 38670 49810
rect 38722 49758 38734 49810
rect 39218 49758 39230 49810
rect 39282 49758 39294 49810
rect 40002 49758 40014 49810
rect 40066 49758 40078 49810
rect 42130 49758 42142 49810
rect 42194 49758 42206 49810
rect 45378 49758 45390 49810
rect 45442 49758 45454 49810
rect 48962 49758 48974 49810
rect 49026 49758 49038 49810
rect 49858 49758 49870 49810
rect 49922 49758 49934 49810
rect 34526 49746 34578 49758
rect 36878 49746 36930 49758
rect 41246 49746 41298 49758
rect 43934 49746 43986 49758
rect 5070 49698 5122 49710
rect 8766 49698 8818 49710
rect 2482 49646 2494 49698
rect 2546 49646 2558 49698
rect 4610 49646 4622 49698
rect 4674 49646 4686 49698
rect 8306 49646 8318 49698
rect 8370 49646 8382 49698
rect 5070 49634 5122 49646
rect 8766 49634 8818 49646
rect 11678 49698 11730 49710
rect 19630 49698 19682 49710
rect 13794 49646 13806 49698
rect 13858 49646 13870 49698
rect 17714 49646 17726 49698
rect 17778 49646 17790 49698
rect 11678 49634 11730 49646
rect 19630 49634 19682 49646
rect 22990 49698 23042 49710
rect 31278 49698 31330 49710
rect 28354 49646 28366 49698
rect 28418 49646 28430 49698
rect 30482 49646 30494 49698
rect 30546 49646 30558 49698
rect 22990 49634 23042 49646
rect 31278 49634 31330 49646
rect 33966 49698 34018 49710
rect 33966 49634 34018 49646
rect 34750 49698 34802 49710
rect 44494 49698 44546 49710
rect 42914 49646 42926 49698
rect 42978 49646 42990 49698
rect 34750 49634 34802 49646
rect 44494 49634 44546 49646
rect 44942 49698 44994 49710
rect 50990 49698 51042 49710
rect 47618 49646 47630 49698
rect 47682 49646 47694 49698
rect 49074 49646 49086 49698
rect 49138 49646 49150 49698
rect 49970 49646 49982 49698
rect 50034 49646 50046 49698
rect 44942 49634 44994 49646
rect 50990 49634 51042 49646
rect 10222 49586 10274 49598
rect 10222 49522 10274 49534
rect 10894 49586 10946 49598
rect 10894 49522 10946 49534
rect 14590 49586 14642 49598
rect 14590 49522 14642 49534
rect 14814 49586 14866 49598
rect 14814 49522 14866 49534
rect 15486 49586 15538 49598
rect 15486 49522 15538 49534
rect 15822 49586 15874 49598
rect 15822 49522 15874 49534
rect 20750 49586 20802 49598
rect 20750 49522 20802 49534
rect 21198 49586 21250 49598
rect 21198 49522 21250 49534
rect 21310 49586 21362 49598
rect 21310 49522 21362 49534
rect 21870 49586 21922 49598
rect 21870 49522 21922 49534
rect 30942 49586 30994 49598
rect 38670 49586 38722 49598
rect 35746 49534 35758 49586
rect 35810 49534 35822 49586
rect 30942 49522 30994 49534
rect 38670 49522 38722 49534
rect 39678 49586 39730 49598
rect 39678 49522 39730 49534
rect 41806 49586 41858 49598
rect 41806 49522 41858 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 4174 49250 4226 49262
rect 4174 49186 4226 49198
rect 4958 49250 5010 49262
rect 4958 49186 5010 49198
rect 6862 49250 6914 49262
rect 6862 49186 6914 49198
rect 7086 49250 7138 49262
rect 22654 49250 22706 49262
rect 21858 49198 21870 49250
rect 21922 49198 21934 49250
rect 7086 49186 7138 49198
rect 22654 49186 22706 49198
rect 36094 49250 36146 49262
rect 36094 49186 36146 49198
rect 39006 49250 39058 49262
rect 39006 49186 39058 49198
rect 43038 49250 43090 49262
rect 43038 49186 43090 49198
rect 49086 49250 49138 49262
rect 49086 49186 49138 49198
rect 50542 49250 50594 49262
rect 50542 49186 50594 49198
rect 7758 49138 7810 49150
rect 23998 49138 24050 49150
rect 16706 49086 16718 49138
rect 16770 49086 16782 49138
rect 19954 49086 19966 49138
rect 20018 49086 20030 49138
rect 7758 49074 7810 49086
rect 23998 49074 24050 49086
rect 28142 49138 28194 49150
rect 28142 49074 28194 49086
rect 29598 49138 29650 49150
rect 34066 49086 34078 49138
rect 34130 49086 34142 49138
rect 37538 49086 37550 49138
rect 37602 49086 37614 49138
rect 40226 49086 40238 49138
rect 40290 49086 40302 49138
rect 44818 49086 44830 49138
rect 44882 49086 44894 49138
rect 29598 49074 29650 49086
rect 4062 49026 4114 49038
rect 4734 49026 4786 49038
rect 4498 48974 4510 49026
rect 4562 48974 4574 49026
rect 4062 48962 4114 48974
rect 4734 48962 4786 48974
rect 5854 49026 5906 49038
rect 5854 48962 5906 48974
rect 6078 49026 6130 49038
rect 6078 48962 6130 48974
rect 7198 49026 7250 49038
rect 7198 48962 7250 48974
rect 9774 49026 9826 49038
rect 9774 48962 9826 48974
rect 9998 49026 10050 49038
rect 16606 49026 16658 49038
rect 21310 49026 21362 49038
rect 10210 48974 10222 49026
rect 10274 48974 10286 49026
rect 13458 48974 13470 49026
rect 13522 48974 13534 49026
rect 17154 48974 17166 49026
rect 17218 48974 17230 49026
rect 9998 48962 10050 48974
rect 16606 48962 16658 48974
rect 21310 48962 21362 48974
rect 21534 49026 21586 49038
rect 24110 49026 24162 49038
rect 22978 48974 22990 49026
rect 23042 48974 23054 49026
rect 21534 48962 21586 48974
rect 24110 48962 24162 48974
rect 27806 49026 27858 49038
rect 29486 49026 29538 49038
rect 28578 48974 28590 49026
rect 28642 48974 28654 49026
rect 29138 48974 29150 49026
rect 29202 48974 29214 49026
rect 27806 48962 27858 48974
rect 29486 48962 29538 48974
rect 30718 49026 30770 49038
rect 34302 49026 34354 49038
rect 31266 48974 31278 49026
rect 31330 48974 31342 49026
rect 30718 48962 30770 48974
rect 34302 48962 34354 48974
rect 36206 49026 36258 49038
rect 36206 48962 36258 48974
rect 37102 49026 37154 49038
rect 38334 49026 38386 49038
rect 37426 48974 37438 49026
rect 37490 48974 37502 49026
rect 37102 48962 37154 48974
rect 38334 48962 38386 48974
rect 39118 49026 39170 49038
rect 39118 48962 39170 48974
rect 39790 49026 39842 49038
rect 39790 48962 39842 48974
rect 40686 49026 40738 49038
rect 40686 48962 40738 48974
rect 41358 49026 41410 49038
rect 41358 48962 41410 48974
rect 41694 49026 41746 49038
rect 41694 48962 41746 48974
rect 42030 49026 42082 49038
rect 42030 48962 42082 48974
rect 42366 49026 42418 49038
rect 42366 48962 42418 48974
rect 43374 49026 43426 49038
rect 50654 49026 50706 49038
rect 44034 48974 44046 49026
rect 44098 48974 44110 49026
rect 47618 48974 47630 49026
rect 47682 48974 47694 49026
rect 49970 48974 49982 49026
rect 50034 48974 50046 49026
rect 43374 48962 43426 48974
rect 50654 48962 50706 48974
rect 50878 49026 50930 49038
rect 50878 48962 50930 48974
rect 3950 48914 4002 48926
rect 3950 48850 4002 48862
rect 6750 48914 6802 48926
rect 6750 48850 6802 48862
rect 7646 48914 7698 48926
rect 7646 48850 7698 48862
rect 9662 48914 9714 48926
rect 20302 48914 20354 48926
rect 14130 48862 14142 48914
rect 14194 48862 14206 48914
rect 15138 48862 15150 48914
rect 15202 48862 15214 48914
rect 17826 48862 17838 48914
rect 17890 48862 17902 48914
rect 9662 48850 9714 48862
rect 20302 48850 20354 48862
rect 20638 48914 20690 48926
rect 20638 48850 20690 48862
rect 23214 48914 23266 48926
rect 23214 48850 23266 48862
rect 23662 48914 23714 48926
rect 23662 48850 23714 48862
rect 23886 48914 23938 48926
rect 23886 48850 23938 48862
rect 27470 48914 27522 48926
rect 27470 48850 27522 48862
rect 27582 48914 27634 48926
rect 34750 48914 34802 48926
rect 30370 48862 30382 48914
rect 30434 48862 30446 48914
rect 31938 48862 31950 48914
rect 32002 48862 32014 48914
rect 27582 48850 27634 48862
rect 34750 48850 34802 48862
rect 34974 48914 35026 48926
rect 34974 48850 35026 48862
rect 37662 48914 37714 48926
rect 41582 48914 41634 48926
rect 39442 48862 39454 48914
rect 39506 48862 39518 48914
rect 37662 48850 37714 48862
rect 41582 48850 41634 48862
rect 42142 48914 42194 48926
rect 49310 48914 49362 48926
rect 50990 48914 51042 48926
rect 44146 48862 44158 48914
rect 44210 48862 44222 48914
rect 46946 48862 46958 48914
rect 47010 48862 47022 48914
rect 49746 48862 49758 48914
rect 49810 48862 49822 48914
rect 42142 48850 42194 48862
rect 49310 48850 49362 48862
rect 50990 48850 51042 48862
rect 4622 48802 4674 48814
rect 7870 48802 7922 48814
rect 6402 48750 6414 48802
rect 6466 48750 6478 48802
rect 4622 48738 4674 48750
rect 7870 48738 7922 48750
rect 8430 48802 8482 48814
rect 11342 48802 11394 48814
rect 10994 48750 11006 48802
rect 11058 48750 11070 48802
rect 8430 48738 8482 48750
rect 11342 48738 11394 48750
rect 22766 48802 22818 48814
rect 22766 48738 22818 48750
rect 25342 48802 25394 48814
rect 26798 48802 26850 48814
rect 25666 48750 25678 48802
rect 25730 48750 25742 48802
rect 25342 48738 25394 48750
rect 26798 48738 26850 48750
rect 27246 48802 27298 48814
rect 27246 48738 27298 48750
rect 28030 48802 28082 48814
rect 28030 48738 28082 48750
rect 28254 48802 28306 48814
rect 28254 48738 28306 48750
rect 29710 48802 29762 48814
rect 29710 48738 29762 48750
rect 34638 48802 34690 48814
rect 34638 48738 34690 48750
rect 35422 48802 35474 48814
rect 35422 48738 35474 48750
rect 36094 48802 36146 48814
rect 51438 48802 51490 48814
rect 37986 48750 37998 48802
rect 38050 48750 38062 48802
rect 48738 48750 48750 48802
rect 48802 48750 48814 48802
rect 36094 48738 36146 48750
rect 51438 48738 51490 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 17502 48466 17554 48478
rect 4274 48414 4286 48466
rect 4338 48414 4350 48466
rect 10322 48414 10334 48466
rect 10386 48414 10398 48466
rect 17502 48402 17554 48414
rect 18398 48466 18450 48478
rect 19854 48466 19906 48478
rect 19394 48414 19406 48466
rect 19458 48414 19470 48466
rect 18398 48402 18450 48414
rect 19854 48402 19906 48414
rect 20078 48466 20130 48478
rect 20078 48402 20130 48414
rect 20526 48466 20578 48478
rect 20526 48402 20578 48414
rect 20974 48466 21026 48478
rect 23998 48466 24050 48478
rect 23314 48414 23326 48466
rect 23378 48414 23390 48466
rect 20974 48402 21026 48414
rect 23998 48402 24050 48414
rect 27582 48466 27634 48478
rect 27582 48402 27634 48414
rect 27694 48466 27746 48478
rect 27694 48402 27746 48414
rect 28814 48466 28866 48478
rect 28814 48402 28866 48414
rect 12126 48354 12178 48366
rect 6738 48302 6750 48354
rect 6802 48302 6814 48354
rect 7858 48302 7870 48354
rect 7922 48302 7934 48354
rect 12126 48290 12178 48302
rect 14142 48354 14194 48366
rect 14142 48290 14194 48302
rect 15598 48354 15650 48366
rect 15598 48290 15650 48302
rect 17726 48354 17778 48366
rect 17726 48290 17778 48302
rect 18622 48354 18674 48366
rect 18622 48290 18674 48302
rect 20414 48354 20466 48366
rect 20414 48290 20466 48302
rect 23774 48354 23826 48366
rect 23774 48290 23826 48302
rect 24670 48354 24722 48366
rect 43262 48354 43314 48366
rect 26674 48302 26686 48354
rect 26738 48302 26750 48354
rect 30706 48302 30718 48354
rect 30770 48302 30782 48354
rect 24670 48290 24722 48302
rect 43262 48290 43314 48302
rect 44046 48354 44098 48366
rect 44046 48290 44098 48302
rect 44494 48354 44546 48366
rect 46946 48302 46958 48354
rect 47010 48302 47022 48354
rect 50082 48302 50094 48354
rect 50146 48302 50158 48354
rect 51202 48302 51214 48354
rect 51266 48302 51278 48354
rect 44494 48290 44546 48302
rect 2830 48242 2882 48254
rect 9774 48242 9826 48254
rect 14702 48242 14754 48254
rect 17278 48242 17330 48254
rect 3042 48190 3054 48242
rect 3106 48190 3118 48242
rect 4050 48190 4062 48242
rect 4114 48190 4126 48242
rect 7522 48190 7534 48242
rect 7586 48190 7598 48242
rect 8082 48190 8094 48242
rect 8146 48190 8158 48242
rect 8642 48190 8654 48242
rect 8706 48190 8718 48242
rect 11330 48190 11342 48242
rect 11394 48190 11406 48242
rect 16818 48190 16830 48242
rect 16882 48190 16894 48242
rect 2830 48178 2882 48190
rect 9774 48178 9826 48190
rect 14702 48178 14754 48190
rect 17278 48178 17330 48190
rect 17950 48242 18002 48254
rect 19742 48242 19794 48254
rect 19170 48190 19182 48242
rect 19234 48190 19246 48242
rect 17950 48178 18002 48190
rect 19742 48178 19794 48190
rect 23662 48242 23714 48254
rect 25790 48242 25842 48254
rect 24322 48190 24334 48242
rect 24386 48190 24398 48242
rect 23662 48178 23714 48190
rect 25790 48178 25842 48190
rect 26014 48242 26066 48254
rect 27806 48242 27858 48254
rect 26450 48190 26462 48242
rect 26514 48190 26526 48242
rect 27346 48190 27358 48242
rect 27410 48190 27422 48242
rect 26014 48178 26066 48190
rect 27806 48178 27858 48190
rect 27918 48242 27970 48254
rect 27918 48178 27970 48190
rect 28702 48242 28754 48254
rect 28702 48178 28754 48190
rect 28926 48242 28978 48254
rect 28926 48178 28978 48190
rect 29374 48242 29426 48254
rect 36206 48242 36258 48254
rect 32498 48190 32510 48242
rect 32562 48190 32574 48242
rect 33282 48190 33294 48242
rect 33346 48190 33358 48242
rect 29374 48178 29426 48190
rect 36206 48178 36258 48190
rect 43374 48242 43426 48254
rect 44606 48242 44658 48254
rect 48638 48242 48690 48254
rect 43810 48190 43822 48242
rect 43874 48190 43886 48242
rect 45378 48190 45390 48242
rect 45442 48190 45454 48242
rect 43374 48178 43426 48190
rect 44606 48178 44658 48190
rect 48638 48178 48690 48190
rect 48974 48242 49026 48254
rect 48974 48178 49026 48190
rect 49198 48242 49250 48254
rect 49198 48178 49250 48190
rect 49758 48242 49810 48254
rect 50530 48190 50542 48242
rect 50594 48190 50606 48242
rect 49758 48178 49810 48190
rect 14814 48130 14866 48142
rect 21422 48130 21474 48142
rect 4610 48078 4622 48130
rect 4674 48078 4686 48130
rect 8754 48078 8766 48130
rect 8818 48078 8830 48130
rect 11666 48078 11678 48130
rect 11730 48078 11742 48130
rect 18386 48078 18398 48130
rect 18450 48078 18462 48130
rect 14814 48066 14866 48078
rect 21422 48066 21474 48078
rect 22766 48130 22818 48142
rect 22766 48066 22818 48078
rect 29150 48130 29202 48142
rect 48190 48130 48242 48142
rect 34290 48078 34302 48130
rect 34354 48078 34366 48130
rect 29150 48066 29202 48078
rect 48190 48066 48242 48078
rect 48862 48130 48914 48142
rect 53330 48078 53342 48130
rect 53394 48078 53406 48130
rect 48862 48066 48914 48078
rect 2718 48018 2770 48030
rect 2718 47954 2770 47966
rect 8990 48018 9042 48030
rect 8990 47954 9042 47966
rect 9998 48018 10050 48030
rect 9998 47954 10050 47966
rect 12350 48018 12402 48030
rect 12350 47954 12402 47966
rect 12686 48018 12738 48030
rect 12686 47954 12738 47966
rect 22990 48018 23042 48030
rect 22990 47954 23042 47966
rect 24334 48018 24386 48030
rect 24334 47954 24386 47966
rect 25454 48018 25506 48030
rect 25454 47954 25506 47966
rect 29598 48018 29650 48030
rect 29598 47954 29650 47966
rect 43262 48018 43314 48030
rect 43262 47954 43314 47966
rect 44718 48018 44770 48030
rect 44718 47954 44770 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 13582 47682 13634 47694
rect 13582 47618 13634 47630
rect 25678 47682 25730 47694
rect 25678 47618 25730 47630
rect 33070 47682 33122 47694
rect 33070 47618 33122 47630
rect 45166 47682 45218 47694
rect 46386 47630 46398 47682
rect 46450 47630 46462 47682
rect 50194 47630 50206 47682
rect 50258 47630 50270 47682
rect 45166 47618 45218 47630
rect 12910 47570 12962 47582
rect 25118 47570 25170 47582
rect 2482 47518 2494 47570
rect 2546 47518 2558 47570
rect 4610 47518 4622 47570
rect 4674 47518 4686 47570
rect 8866 47518 8878 47570
rect 8930 47518 8942 47570
rect 10994 47518 11006 47570
rect 11058 47518 11070 47570
rect 18946 47518 18958 47570
rect 19010 47518 19022 47570
rect 12910 47506 12962 47518
rect 25118 47506 25170 47518
rect 27246 47570 27298 47582
rect 31054 47570 31106 47582
rect 29362 47518 29374 47570
rect 29426 47518 29438 47570
rect 29698 47518 29710 47570
rect 29762 47518 29774 47570
rect 27246 47506 27298 47518
rect 31054 47506 31106 47518
rect 31838 47570 31890 47582
rect 49646 47570 49698 47582
rect 36418 47518 36430 47570
rect 36482 47518 36494 47570
rect 44258 47518 44270 47570
rect 44322 47518 44334 47570
rect 47954 47518 47966 47570
rect 48018 47518 48030 47570
rect 31838 47506 31890 47518
rect 49646 47506 49698 47518
rect 51326 47570 51378 47582
rect 51326 47506 51378 47518
rect 13470 47458 13522 47470
rect 18510 47458 18562 47470
rect 21310 47458 21362 47470
rect 1810 47406 1822 47458
rect 1874 47406 1886 47458
rect 5954 47406 5966 47458
rect 6018 47406 6030 47458
rect 7074 47406 7086 47458
rect 7138 47406 7150 47458
rect 8082 47406 8094 47458
rect 8146 47406 8158 47458
rect 14018 47406 14030 47458
rect 14082 47406 14094 47458
rect 17826 47406 17838 47458
rect 17890 47406 17902 47458
rect 19618 47406 19630 47458
rect 19682 47406 19694 47458
rect 20514 47406 20526 47458
rect 20578 47406 20590 47458
rect 13470 47394 13522 47406
rect 18510 47394 18562 47406
rect 21310 47394 21362 47406
rect 22766 47458 22818 47470
rect 22766 47394 22818 47406
rect 23102 47458 23154 47470
rect 27694 47458 27746 47470
rect 25666 47406 25678 47458
rect 25730 47406 25742 47458
rect 23102 47394 23154 47406
rect 27694 47394 27746 47406
rect 27918 47458 27970 47470
rect 27918 47394 27970 47406
rect 28478 47458 28530 47470
rect 30830 47458 30882 47470
rect 32174 47458 32226 47470
rect 29026 47406 29038 47458
rect 29090 47406 29102 47458
rect 29810 47406 29822 47458
rect 29874 47406 29886 47458
rect 31154 47406 31166 47458
rect 31218 47406 31230 47458
rect 28478 47394 28530 47406
rect 30830 47394 30882 47406
rect 32174 47394 32226 47406
rect 32734 47458 32786 47470
rect 32734 47394 32786 47406
rect 33182 47458 33234 47470
rect 44942 47458 44994 47470
rect 45838 47458 45890 47470
rect 48302 47458 48354 47470
rect 33506 47406 33518 47458
rect 33570 47406 33582 47458
rect 41458 47406 41470 47458
rect 41522 47406 41534 47458
rect 45378 47406 45390 47458
rect 45442 47406 45454 47458
rect 46050 47406 46062 47458
rect 46114 47406 46126 47458
rect 46498 47406 46510 47458
rect 46562 47406 46574 47458
rect 47282 47406 47294 47458
rect 47346 47406 47358 47458
rect 47618 47406 47630 47458
rect 47682 47406 47694 47458
rect 33182 47394 33234 47406
rect 44942 47394 44994 47406
rect 45838 47394 45890 47406
rect 48302 47394 48354 47406
rect 48526 47458 48578 47470
rect 48526 47394 48578 47406
rect 48750 47458 48802 47470
rect 48750 47394 48802 47406
rect 49870 47458 49922 47470
rect 51214 47458 51266 47470
rect 50642 47406 50654 47458
rect 50706 47406 50718 47458
rect 51538 47406 51550 47458
rect 51602 47406 51614 47458
rect 49870 47394 49922 47406
rect 51214 47394 51266 47406
rect 17166 47346 17218 47358
rect 6066 47294 6078 47346
rect 6130 47294 6142 47346
rect 7522 47294 7534 47346
rect 7586 47294 7598 47346
rect 14130 47294 14142 47346
rect 14194 47294 14206 47346
rect 17166 47282 17218 47294
rect 19406 47346 19458 47358
rect 19406 47282 19458 47294
rect 22542 47346 22594 47358
rect 22542 47282 22594 47294
rect 25342 47346 25394 47358
rect 25342 47282 25394 47294
rect 27582 47346 27634 47358
rect 27582 47282 27634 47294
rect 28366 47346 28418 47358
rect 28366 47282 28418 47294
rect 31390 47346 31442 47358
rect 44830 47346 44882 47358
rect 34290 47294 34302 47346
rect 34354 47294 34366 47346
rect 42130 47294 42142 47346
rect 42194 47294 42206 47346
rect 31390 47282 31442 47294
rect 44830 47282 44882 47294
rect 49086 47346 49138 47358
rect 49086 47282 49138 47294
rect 5070 47234 5122 47246
rect 12798 47234 12850 47246
rect 6962 47182 6974 47234
rect 7026 47182 7038 47234
rect 5070 47170 5122 47182
rect 12798 47170 12850 47182
rect 13582 47234 13634 47246
rect 21422 47234 21474 47246
rect 15586 47182 15598 47234
rect 15650 47182 15662 47234
rect 20738 47182 20750 47234
rect 20802 47182 20814 47234
rect 13582 47170 13634 47182
rect 21422 47170 21474 47182
rect 21646 47234 21698 47246
rect 21646 47170 21698 47182
rect 22766 47234 22818 47246
rect 22766 47170 22818 47182
rect 24110 47234 24162 47246
rect 24110 47170 24162 47182
rect 24558 47234 24610 47246
rect 24558 47170 24610 47182
rect 26238 47234 26290 47246
rect 28142 47234 28194 47246
rect 26562 47182 26574 47234
rect 26626 47182 26638 47234
rect 26238 47170 26290 47182
rect 28142 47170 28194 47182
rect 37102 47234 37154 47246
rect 37102 47170 37154 47182
rect 46622 47234 46674 47246
rect 46622 47170 46674 47182
rect 48638 47234 48690 47246
rect 50866 47182 50878 47234
rect 50930 47182 50942 47234
rect 48638 47170 48690 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 15710 46898 15762 46910
rect 15710 46834 15762 46846
rect 16382 46898 16434 46910
rect 16382 46834 16434 46846
rect 19294 46898 19346 46910
rect 19294 46834 19346 46846
rect 19742 46898 19794 46910
rect 24110 46898 24162 46910
rect 20738 46846 20750 46898
rect 20802 46846 20814 46898
rect 19742 46834 19794 46846
rect 24110 46834 24162 46846
rect 27358 46898 27410 46910
rect 27358 46834 27410 46846
rect 28814 46898 28866 46910
rect 28814 46834 28866 46846
rect 28926 46898 28978 46910
rect 28926 46834 28978 46846
rect 29710 46898 29762 46910
rect 29710 46834 29762 46846
rect 30158 46898 30210 46910
rect 35758 46898 35810 46910
rect 33058 46846 33070 46898
rect 33122 46846 33134 46898
rect 30158 46834 30210 46846
rect 35758 46834 35810 46846
rect 51102 46898 51154 46910
rect 51102 46834 51154 46846
rect 2494 46786 2546 46798
rect 2494 46722 2546 46734
rect 3950 46786 4002 46798
rect 3950 46722 4002 46734
rect 6414 46786 6466 46798
rect 6414 46722 6466 46734
rect 12126 46786 12178 46798
rect 15486 46786 15538 46798
rect 13346 46734 13358 46786
rect 13410 46734 13422 46786
rect 13906 46734 13918 46786
rect 13970 46734 13982 46786
rect 12126 46722 12178 46734
rect 15486 46722 15538 46734
rect 16270 46786 16322 46798
rect 23102 46786 23154 46798
rect 22866 46734 22878 46786
rect 22930 46734 22942 46786
rect 16270 46722 16322 46734
rect 23102 46722 23154 46734
rect 26686 46786 26738 46798
rect 26686 46722 26738 46734
rect 28142 46786 28194 46798
rect 28142 46722 28194 46734
rect 28478 46786 28530 46798
rect 28478 46722 28530 46734
rect 28590 46786 28642 46798
rect 28590 46722 28642 46734
rect 29150 46786 29202 46798
rect 29150 46722 29202 46734
rect 29262 46786 29314 46798
rect 29262 46722 29314 46734
rect 29822 46786 29874 46798
rect 30942 46786 30994 46798
rect 30482 46734 30494 46786
rect 30546 46734 30558 46786
rect 29822 46722 29874 46734
rect 30942 46722 30994 46734
rect 31166 46786 31218 46798
rect 32398 46786 32450 46798
rect 32050 46734 32062 46786
rect 32114 46734 32126 46786
rect 31166 46722 31218 46734
rect 32398 46722 32450 46734
rect 34414 46786 34466 46798
rect 34414 46722 34466 46734
rect 34638 46786 34690 46798
rect 34638 46722 34690 46734
rect 47182 46786 47234 46798
rect 47182 46722 47234 46734
rect 3390 46674 3442 46686
rect 3154 46622 3166 46674
rect 3218 46622 3230 46674
rect 3390 46610 3442 46622
rect 3726 46674 3778 46686
rect 3726 46610 3778 46622
rect 4062 46674 4114 46686
rect 11230 46674 11282 46686
rect 10994 46622 11006 46674
rect 11058 46622 11070 46674
rect 4062 46610 4114 46622
rect 11230 46610 11282 46622
rect 11566 46674 11618 46686
rect 13694 46674 13746 46686
rect 16046 46674 16098 46686
rect 12002 46622 12014 46674
rect 12066 46622 12078 46674
rect 12786 46622 12798 46674
rect 12850 46622 12862 46674
rect 13122 46622 13134 46674
rect 13186 46622 13198 46674
rect 14354 46622 14366 46674
rect 14418 46622 14430 46674
rect 15138 46622 15150 46674
rect 15202 46622 15214 46674
rect 11566 46610 11618 46622
rect 13694 46610 13746 46622
rect 16046 46610 16098 46622
rect 17726 46674 17778 46686
rect 17726 46610 17778 46622
rect 17950 46674 18002 46686
rect 19518 46674 19570 46686
rect 18610 46622 18622 46674
rect 18674 46622 18686 46674
rect 17950 46610 18002 46622
rect 19518 46610 19570 46622
rect 20414 46674 20466 46686
rect 21758 46674 21810 46686
rect 21298 46622 21310 46674
rect 21362 46622 21374 46674
rect 20414 46610 20466 46622
rect 21758 46610 21810 46622
rect 22094 46674 22146 46686
rect 25342 46674 25394 46686
rect 28030 46674 28082 46686
rect 22306 46622 22318 46674
rect 22370 46622 22382 46674
rect 23426 46622 23438 46674
rect 23490 46622 23502 46674
rect 25666 46622 25678 46674
rect 25730 46622 25742 46674
rect 27122 46622 27134 46674
rect 27186 46622 27198 46674
rect 22094 46610 22146 46622
rect 25342 46610 25394 46622
rect 28030 46610 28082 46622
rect 30830 46674 30882 46686
rect 30830 46610 30882 46622
rect 31278 46674 31330 46686
rect 31278 46610 31330 46622
rect 31726 46674 31778 46686
rect 33966 46674 34018 46686
rect 39678 46674 39730 46686
rect 44494 46674 44546 46686
rect 33282 46622 33294 46674
rect 33346 46622 33358 46674
rect 36306 46622 36318 46674
rect 36370 46622 36382 46674
rect 40002 46622 40014 46674
rect 40066 46622 40078 46674
rect 41010 46622 41022 46674
rect 41074 46622 41086 46674
rect 31726 46610 31778 46622
rect 33966 46610 34018 46622
rect 39678 46610 39730 46622
rect 44494 46610 44546 46622
rect 44718 46674 44770 46686
rect 44718 46610 44770 46622
rect 45838 46674 45890 46686
rect 45838 46610 45890 46622
rect 46062 46674 46114 46686
rect 46062 46610 46114 46622
rect 47070 46674 47122 46686
rect 49758 46674 49810 46686
rect 50318 46674 50370 46686
rect 47394 46622 47406 46674
rect 47458 46622 47470 46674
rect 49298 46622 49310 46674
rect 49362 46622 49374 46674
rect 50082 46622 50094 46674
rect 50146 46622 50158 46674
rect 47070 46610 47122 46622
rect 49758 46610 49810 46622
rect 50318 46610 50370 46622
rect 50542 46674 50594 46686
rect 50542 46610 50594 46622
rect 7758 46562 7810 46574
rect 7758 46498 7810 46510
rect 10558 46562 10610 46574
rect 19406 46562 19458 46574
rect 18722 46510 18734 46562
rect 18786 46510 18798 46562
rect 10558 46498 10610 46510
rect 19406 46498 19458 46510
rect 20190 46562 20242 46574
rect 20190 46498 20242 46510
rect 24670 46562 24722 46574
rect 24670 46498 24722 46510
rect 26238 46562 26290 46574
rect 35422 46562 35474 46574
rect 40238 46562 40290 46574
rect 46174 46562 46226 46574
rect 34290 46510 34302 46562
rect 34354 46510 34366 46562
rect 37090 46510 37102 46562
rect 37154 46510 37166 46562
rect 39218 46510 39230 46562
rect 39282 46510 39294 46562
rect 41682 46510 41694 46562
rect 41746 46510 41758 46562
rect 43810 46510 43822 46562
rect 43874 46510 43886 46562
rect 46610 46510 46622 46562
rect 46674 46510 46686 46562
rect 48850 46510 48862 46562
rect 48914 46510 48926 46562
rect 26238 46498 26290 46510
rect 35422 46498 35474 46510
rect 40238 46498 40290 46510
rect 46174 46498 46226 46510
rect 6302 46450 6354 46462
rect 6302 46386 6354 46398
rect 6638 46450 6690 46462
rect 6638 46386 6690 46398
rect 10670 46450 10722 46462
rect 10670 46386 10722 46398
rect 11454 46450 11506 46462
rect 15822 46450 15874 46462
rect 14018 46398 14030 46450
rect 14082 46398 14094 46450
rect 11454 46386 11506 46398
rect 15822 46386 15874 46398
rect 16382 46450 16434 46462
rect 16382 46386 16434 46398
rect 17390 46450 17442 46462
rect 17390 46386 17442 46398
rect 26798 46450 26850 46462
rect 26798 46386 26850 46398
rect 27470 46450 27522 46462
rect 27470 46386 27522 46398
rect 29710 46450 29762 46462
rect 29710 46386 29762 46398
rect 32510 46450 32562 46462
rect 40350 46450 40402 46462
rect 45726 46450 45778 46462
rect 35410 46398 35422 46450
rect 35474 46447 35486 46450
rect 35970 46447 35982 46450
rect 35474 46401 35982 46447
rect 35474 46398 35486 46401
rect 35970 46398 35982 46401
rect 36034 46398 36046 46450
rect 45042 46398 45054 46450
rect 45106 46398 45118 46450
rect 32510 46386 32562 46398
rect 40350 46386 40402 46398
rect 45726 46386 45778 46398
rect 50654 46450 50706 46462
rect 50654 46386 50706 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 14926 46114 14978 46126
rect 6402 46062 6414 46114
rect 6466 46062 6478 46114
rect 14926 46050 14978 46062
rect 17166 46114 17218 46126
rect 17166 46050 17218 46062
rect 23438 46114 23490 46126
rect 23438 46050 23490 46062
rect 23662 46114 23714 46126
rect 23662 46050 23714 46062
rect 31390 46114 31442 46126
rect 51550 46114 51602 46126
rect 43810 46062 43822 46114
rect 43874 46111 43886 46114
rect 44370 46111 44382 46114
rect 43874 46065 44382 46111
rect 43874 46062 43886 46065
rect 44370 46062 44382 46065
rect 44434 46062 44446 46114
rect 31390 46050 31442 46062
rect 51550 46050 51602 46062
rect 11790 46002 11842 46014
rect 4610 45950 4622 46002
rect 4674 45950 4686 46002
rect 10882 45950 10894 46002
rect 10946 45950 10958 46002
rect 11790 45938 11842 45950
rect 13694 46002 13746 46014
rect 13694 45938 13746 45950
rect 14590 46002 14642 46014
rect 14590 45938 14642 45950
rect 15038 46002 15090 46014
rect 21758 46002 21810 46014
rect 29486 46002 29538 46014
rect 19842 45950 19854 46002
rect 19906 45950 19918 46002
rect 24210 45950 24222 46002
rect 24274 45950 24286 46002
rect 15038 45938 15090 45950
rect 21758 45938 21810 45950
rect 29486 45938 29538 45950
rect 31838 46002 31890 46014
rect 40238 46002 40290 46014
rect 32946 45950 32958 46002
rect 33010 45950 33022 46002
rect 39554 45950 39566 46002
rect 39618 45950 39630 46002
rect 47282 45950 47294 46002
rect 47346 45950 47358 46002
rect 49410 45950 49422 46002
rect 49474 45950 49486 46002
rect 31838 45938 31890 45950
rect 40238 45938 40290 45950
rect 5630 45890 5682 45902
rect 12574 45890 12626 45902
rect 18846 45890 18898 45902
rect 1810 45838 1822 45890
rect 1874 45838 1886 45890
rect 6178 45838 6190 45890
rect 6242 45838 6254 45890
rect 7074 45838 7086 45890
rect 7138 45838 7150 45890
rect 7970 45838 7982 45890
rect 8034 45838 8046 45890
rect 14130 45838 14142 45890
rect 14194 45838 14206 45890
rect 17714 45838 17726 45890
rect 17778 45838 17790 45890
rect 5630 45826 5682 45838
rect 12574 45826 12626 45838
rect 18846 45826 18898 45838
rect 20638 45890 20690 45902
rect 20638 45826 20690 45838
rect 21310 45890 21362 45902
rect 21310 45826 21362 45838
rect 21534 45890 21586 45902
rect 21534 45826 21586 45838
rect 22542 45890 22594 45902
rect 23886 45890 23938 45902
rect 22978 45838 22990 45890
rect 23042 45838 23054 45890
rect 22542 45826 22594 45838
rect 23886 45826 23938 45838
rect 25006 45890 25058 45902
rect 26798 45890 26850 45902
rect 25330 45838 25342 45890
rect 25394 45838 25406 45890
rect 25006 45826 25058 45838
rect 26798 45826 26850 45838
rect 27582 45890 27634 45902
rect 27582 45826 27634 45838
rect 28030 45890 28082 45902
rect 32510 45890 32562 45902
rect 39902 45890 39954 45902
rect 44046 45890 44098 45902
rect 29362 45838 29374 45890
rect 29426 45838 29438 45890
rect 29586 45838 29598 45890
rect 29650 45838 29662 45890
rect 30034 45838 30046 45890
rect 30098 45838 30110 45890
rect 31042 45838 31054 45890
rect 31106 45838 31118 45890
rect 32050 45838 32062 45890
rect 32114 45838 32126 45890
rect 39218 45838 39230 45890
rect 39282 45838 39294 45890
rect 40450 45838 40462 45890
rect 40514 45838 40526 45890
rect 40898 45838 40910 45890
rect 40962 45838 40974 45890
rect 28030 45826 28082 45838
rect 32510 45826 32562 45838
rect 39902 45826 39954 45838
rect 44046 45826 44098 45838
rect 44942 45890 44994 45902
rect 45826 45838 45838 45890
rect 45890 45838 45902 45890
rect 46610 45838 46622 45890
rect 46674 45838 46686 45890
rect 44942 45826 44994 45838
rect 15710 45778 15762 45790
rect 2482 45726 2494 45778
rect 2546 45726 2558 45778
rect 5842 45726 5854 45778
rect 5906 45726 5918 45778
rect 8754 45726 8766 45778
rect 8818 45726 8830 45778
rect 12898 45726 12910 45778
rect 12962 45726 12974 45778
rect 15710 45714 15762 45726
rect 15822 45778 15874 45790
rect 15822 45714 15874 45726
rect 17054 45778 17106 45790
rect 17054 45714 17106 45726
rect 18286 45778 18338 45790
rect 25902 45778 25954 45790
rect 20290 45726 20302 45778
rect 20354 45726 20366 45778
rect 18286 45714 18338 45726
rect 25902 45714 25954 45726
rect 28254 45778 28306 45790
rect 28254 45714 28306 45726
rect 29150 45778 29202 45790
rect 31726 45778 31778 45790
rect 51662 45778 51714 45790
rect 30146 45726 30158 45778
rect 30210 45726 30222 45778
rect 30706 45726 30718 45778
rect 30770 45726 30782 45778
rect 45602 45726 45614 45778
rect 45666 45726 45678 45778
rect 29150 45714 29202 45726
rect 31726 45714 31778 45726
rect 51662 45714 51714 45726
rect 5070 45666 5122 45678
rect 5070 45602 5122 45614
rect 7646 45666 7698 45678
rect 7646 45602 7698 45614
rect 16046 45666 16098 45678
rect 16046 45602 16098 45614
rect 17166 45666 17218 45678
rect 19406 45666 19458 45678
rect 17938 45614 17950 45666
rect 18002 45614 18014 45666
rect 17166 45602 17218 45614
rect 19406 45602 19458 45614
rect 22206 45666 22258 45678
rect 22206 45602 22258 45614
rect 24110 45666 24162 45678
rect 24110 45602 24162 45614
rect 24334 45666 24386 45678
rect 24334 45602 24386 45614
rect 25566 45666 25618 45678
rect 25566 45602 25618 45614
rect 25678 45666 25730 45678
rect 25678 45602 25730 45614
rect 26014 45666 26066 45678
rect 26014 45602 26066 45614
rect 26238 45666 26290 45678
rect 26238 45602 26290 45614
rect 26910 45666 26962 45678
rect 26910 45602 26962 45614
rect 27022 45666 27074 45678
rect 27022 45602 27074 45614
rect 27246 45666 27298 45678
rect 27246 45602 27298 45614
rect 27806 45666 27858 45678
rect 27806 45602 27858 45614
rect 31278 45666 31330 45678
rect 31278 45602 31330 45614
rect 49870 45666 49922 45678
rect 49870 45602 49922 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 2606 45330 2658 45342
rect 2606 45266 2658 45278
rect 5630 45330 5682 45342
rect 5630 45266 5682 45278
rect 9998 45330 10050 45342
rect 14478 45330 14530 45342
rect 12338 45278 12350 45330
rect 12402 45278 12414 45330
rect 9998 45266 10050 45278
rect 14478 45266 14530 45278
rect 14702 45330 14754 45342
rect 14702 45266 14754 45278
rect 15150 45330 15202 45342
rect 15150 45266 15202 45278
rect 16830 45330 16882 45342
rect 16830 45266 16882 45278
rect 25678 45330 25730 45342
rect 25678 45266 25730 45278
rect 39678 45330 39730 45342
rect 39678 45266 39730 45278
rect 44494 45330 44546 45342
rect 44494 45266 44546 45278
rect 2494 45218 2546 45230
rect 2494 45154 2546 45166
rect 4510 45218 4562 45230
rect 4510 45154 4562 45166
rect 5966 45218 6018 45230
rect 5966 45154 6018 45166
rect 8654 45218 8706 45230
rect 8654 45154 8706 45166
rect 8990 45218 9042 45230
rect 8990 45154 9042 45166
rect 15374 45218 15426 45230
rect 18398 45218 18450 45230
rect 32286 45218 32338 45230
rect 17714 45166 17726 45218
rect 17778 45166 17790 45218
rect 25890 45166 25902 45218
rect 25954 45166 25966 45218
rect 27906 45166 27918 45218
rect 27970 45166 27982 45218
rect 31378 45166 31390 45218
rect 31442 45166 31454 45218
rect 15374 45154 15426 45166
rect 18398 45154 18450 45166
rect 32286 45154 32338 45166
rect 32510 45218 32562 45230
rect 39566 45218 39618 45230
rect 38546 45166 38558 45218
rect 38610 45166 38622 45218
rect 32510 45154 32562 45166
rect 39566 45154 39618 45166
rect 40238 45218 40290 45230
rect 40238 45154 40290 45166
rect 40350 45218 40402 45230
rect 40350 45154 40402 45166
rect 41470 45218 41522 45230
rect 41470 45154 41522 45166
rect 42366 45218 42418 45230
rect 50194 45166 50206 45218
rect 50258 45166 50270 45218
rect 42366 45154 42418 45166
rect 2718 45106 2770 45118
rect 2718 45042 2770 45054
rect 3166 45106 3218 45118
rect 12014 45106 12066 45118
rect 4946 45054 4958 45106
rect 5010 45054 5022 45106
rect 5394 45054 5406 45106
rect 5458 45054 5470 45106
rect 10658 45054 10670 45106
rect 10722 45054 10734 45106
rect 10994 45054 11006 45106
rect 11058 45054 11070 45106
rect 3166 45042 3218 45054
rect 12014 45042 12066 45054
rect 14366 45106 14418 45118
rect 14366 45042 14418 45054
rect 15486 45106 15538 45118
rect 18958 45106 19010 45118
rect 33742 45106 33794 45118
rect 18050 45054 18062 45106
rect 18114 45054 18126 45106
rect 18610 45054 18622 45106
rect 18674 45054 18686 45106
rect 20626 45054 20638 45106
rect 20690 45054 20702 45106
rect 21522 45054 21534 45106
rect 21586 45054 21598 45106
rect 23202 45054 23214 45106
rect 23266 45054 23278 45106
rect 23874 45054 23886 45106
rect 23938 45054 23950 45106
rect 26674 45054 26686 45106
rect 26738 45054 26750 45106
rect 27234 45054 27246 45106
rect 27298 45054 27310 45106
rect 27458 45054 27470 45106
rect 27522 45054 27534 45106
rect 28914 45054 28926 45106
rect 28978 45054 28990 45106
rect 30034 45054 30046 45106
rect 30098 45054 30110 45106
rect 30706 45054 30718 45106
rect 30770 45054 30782 45106
rect 31266 45054 31278 45106
rect 31330 45054 31342 45106
rect 15486 45042 15538 45054
rect 18958 45042 19010 45054
rect 33742 45042 33794 45054
rect 33966 45106 34018 45118
rect 33966 45042 34018 45054
rect 34414 45106 34466 45118
rect 41022 45106 41074 45118
rect 34738 45054 34750 45106
rect 34802 45054 34814 45106
rect 38322 45054 38334 45106
rect 38386 45054 38398 45106
rect 34414 45042 34466 45054
rect 41022 45042 41074 45054
rect 41582 45106 41634 45118
rect 41582 45042 41634 45054
rect 41694 45106 41746 45118
rect 41694 45042 41746 45054
rect 41918 45106 41970 45118
rect 41918 45042 41970 45054
rect 42478 45106 42530 45118
rect 49410 45054 49422 45106
rect 49474 45054 49486 45106
rect 42478 45042 42530 45054
rect 11790 44994 11842 45006
rect 10546 44942 10558 44994
rect 10610 44942 10622 44994
rect 11790 44930 11842 44942
rect 15934 44994 15986 45006
rect 15934 44930 15986 44942
rect 16718 44994 16770 45006
rect 28702 44994 28754 45006
rect 33406 44994 33458 45006
rect 20290 44942 20302 44994
rect 20354 44942 20366 44994
rect 23538 44942 23550 44994
rect 23602 44942 23614 44994
rect 26338 44942 26350 44994
rect 26402 44942 26414 44994
rect 29250 44942 29262 44994
rect 29314 44942 29326 44994
rect 29586 44942 29598 44994
rect 29650 44942 29662 44994
rect 31378 44942 31390 44994
rect 31442 44942 31454 44994
rect 16718 44930 16770 44942
rect 28702 44930 28754 44942
rect 33406 44930 33458 44942
rect 34190 44994 34242 45006
rect 42142 44994 42194 45006
rect 35410 44942 35422 44994
rect 35474 44942 35486 44994
rect 37538 44942 37550 44994
rect 37602 44942 37614 44994
rect 40786 44942 40798 44994
rect 40850 44991 40862 44994
rect 41010 44991 41022 44994
rect 40850 44945 41022 44991
rect 40850 44942 40862 44945
rect 41010 44942 41022 44945
rect 41074 44942 41086 44994
rect 34190 44930 34242 44942
rect 42142 44930 42194 44942
rect 49086 44994 49138 45006
rect 52322 44942 52334 44994
rect 52386 44942 52398 44994
rect 49086 44930 49138 44942
rect 17950 44882 18002 44894
rect 17950 44818 18002 44830
rect 18286 44882 18338 44894
rect 18286 44818 18338 44830
rect 32174 44882 32226 44894
rect 32174 44818 32226 44830
rect 39678 44882 39730 44894
rect 39678 44818 39730 44830
rect 40238 44882 40290 44894
rect 40238 44818 40290 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 3614 44546 3666 44558
rect 3614 44482 3666 44494
rect 4174 44546 4226 44558
rect 4174 44482 4226 44494
rect 10110 44546 10162 44558
rect 10110 44482 10162 44494
rect 10446 44546 10498 44558
rect 17502 44546 17554 44558
rect 15474 44494 15486 44546
rect 15538 44543 15550 44546
rect 16482 44543 16494 44546
rect 15538 44497 16494 44543
rect 15538 44494 15550 44497
rect 16482 44494 16494 44497
rect 16546 44494 16558 44546
rect 10446 44482 10498 44494
rect 17502 44482 17554 44494
rect 29150 44546 29202 44558
rect 29150 44482 29202 44494
rect 29374 44546 29426 44558
rect 29374 44482 29426 44494
rect 32510 44546 32562 44558
rect 32510 44482 32562 44494
rect 34638 44546 34690 44558
rect 34638 44482 34690 44494
rect 2494 44434 2546 44446
rect 10222 44434 10274 44446
rect 8530 44382 8542 44434
rect 8594 44382 8606 44434
rect 2494 44370 2546 44382
rect 10222 44370 10274 44382
rect 11790 44434 11842 44446
rect 11790 44370 11842 44382
rect 16606 44434 16658 44446
rect 16606 44370 16658 44382
rect 17054 44434 17106 44446
rect 30942 44434 30994 44446
rect 37774 44434 37826 44446
rect 24994 44382 25006 44434
rect 25058 44382 25070 44434
rect 25778 44382 25790 44434
rect 25842 44382 25854 44434
rect 32834 44382 32846 44434
rect 32898 44382 32910 44434
rect 34066 44382 34078 44434
rect 34130 44382 34142 44434
rect 17054 44370 17106 44382
rect 30942 44370 30994 44382
rect 37774 44370 37826 44382
rect 39342 44434 39394 44446
rect 40798 44434 40850 44446
rect 40114 44382 40126 44434
rect 40178 44382 40190 44434
rect 41906 44382 41918 44434
rect 41970 44382 41982 44434
rect 44818 44382 44830 44434
rect 44882 44382 44894 44434
rect 39342 44370 39394 44382
rect 40798 44370 40850 44382
rect 2270 44322 2322 44334
rect 2270 44258 2322 44270
rect 2718 44322 2770 44334
rect 2718 44258 2770 44270
rect 2830 44322 2882 44334
rect 2830 44258 2882 44270
rect 3390 44322 3442 44334
rect 3390 44258 3442 44270
rect 3726 44322 3778 44334
rect 3726 44258 3778 44270
rect 4510 44322 4562 44334
rect 4510 44258 4562 44270
rect 4958 44322 5010 44334
rect 11118 44322 11170 44334
rect 5618 44270 5630 44322
rect 5682 44270 5694 44322
rect 10658 44270 10670 44322
rect 10722 44270 10734 44322
rect 4958 44258 5010 44270
rect 11118 44258 11170 44270
rect 11454 44322 11506 44334
rect 13582 44322 13634 44334
rect 12562 44270 12574 44322
rect 12626 44270 12638 44322
rect 11454 44258 11506 44270
rect 13582 44258 13634 44270
rect 13694 44322 13746 44334
rect 13694 44258 13746 44270
rect 14030 44322 14082 44334
rect 14030 44258 14082 44270
rect 14254 44322 14306 44334
rect 14254 44258 14306 44270
rect 14478 44322 14530 44334
rect 14478 44258 14530 44270
rect 15038 44322 15090 44334
rect 15038 44258 15090 44270
rect 17278 44322 17330 44334
rect 17278 44258 17330 44270
rect 17950 44322 18002 44334
rect 19854 44322 19906 44334
rect 28254 44322 28306 44334
rect 18274 44270 18286 44322
rect 18338 44270 18350 44322
rect 18610 44270 18622 44322
rect 18674 44270 18686 44322
rect 19394 44270 19406 44322
rect 19458 44270 19470 44322
rect 22306 44270 22318 44322
rect 22370 44270 22382 44322
rect 23314 44270 23326 44322
rect 23378 44270 23390 44322
rect 25666 44270 25678 44322
rect 25730 44270 25742 44322
rect 26450 44270 26462 44322
rect 26514 44270 26526 44322
rect 27346 44270 27358 44322
rect 27410 44270 27422 44322
rect 17950 44258 18002 44270
rect 19854 44258 19906 44270
rect 28254 44258 28306 44270
rect 28590 44322 28642 44334
rect 28590 44258 28642 44270
rect 29598 44322 29650 44334
rect 29598 44258 29650 44270
rect 29822 44322 29874 44334
rect 29822 44258 29874 44270
rect 30046 44322 30098 44334
rect 30046 44258 30098 44270
rect 30382 44322 30434 44334
rect 30382 44258 30434 44270
rect 31278 44322 31330 44334
rect 31278 44258 31330 44270
rect 31614 44322 31666 44334
rect 31614 44258 31666 44270
rect 31950 44322 32002 44334
rect 33742 44322 33794 44334
rect 33506 44270 33518 44322
rect 33570 44270 33582 44322
rect 31950 44258 32002 44270
rect 33742 44258 33794 44270
rect 38782 44322 38834 44334
rect 39778 44270 39790 44322
rect 39842 44270 39854 44322
rect 41234 44270 41246 44322
rect 41298 44270 41310 44322
rect 47730 44270 47742 44322
rect 47794 44270 47806 44322
rect 38782 44258 38834 44270
rect 3278 44210 3330 44222
rect 11230 44210 11282 44222
rect 6402 44158 6414 44210
rect 6466 44158 6478 44210
rect 3278 44146 3330 44158
rect 11230 44146 11282 44158
rect 12238 44210 12290 44222
rect 12238 44146 12290 44158
rect 14926 44210 14978 44222
rect 14926 44146 14978 44158
rect 15486 44210 15538 44222
rect 15486 44146 15538 44158
rect 15934 44210 15986 44222
rect 15934 44146 15986 44158
rect 17726 44210 17778 44222
rect 17726 44146 17778 44158
rect 19294 44210 19346 44222
rect 28478 44210 28530 44222
rect 22194 44158 22206 44210
rect 22258 44158 22270 44210
rect 23202 44158 23214 44210
rect 23266 44158 23278 44210
rect 26002 44158 26014 44210
rect 26066 44158 26078 44210
rect 26674 44158 26686 44210
rect 26738 44158 26750 44210
rect 19294 44146 19346 44158
rect 28478 44146 28530 44158
rect 33966 44210 34018 44222
rect 33966 44146 34018 44158
rect 34526 44210 34578 44222
rect 38434 44158 38446 44210
rect 38498 44158 38510 44210
rect 46946 44158 46958 44210
rect 47010 44158 47022 44210
rect 34526 44146 34578 44158
rect 4286 44098 4338 44110
rect 4286 44034 4338 44046
rect 5070 44098 5122 44110
rect 5070 44034 5122 44046
rect 9102 44098 9154 44110
rect 9102 44034 9154 44046
rect 9550 44098 9602 44110
rect 9550 44034 9602 44046
rect 12350 44098 12402 44110
rect 12350 44034 12402 44046
rect 13806 44098 13858 44110
rect 13806 44034 13858 44046
rect 14702 44098 14754 44110
rect 14702 44034 14754 44046
rect 16494 44098 16546 44110
rect 16494 44034 16546 44046
rect 20190 44098 20242 44110
rect 20190 44034 20242 44046
rect 29934 44098 29986 44110
rect 29934 44034 29986 44046
rect 30830 44098 30882 44110
rect 30830 44034 30882 44046
rect 31054 44098 31106 44110
rect 31054 44034 31106 44046
rect 31614 44098 31666 44110
rect 31614 44034 31666 44046
rect 32734 44098 32786 44110
rect 32734 44034 32786 44046
rect 34078 44098 34130 44110
rect 34078 44034 34130 44046
rect 34638 44098 34690 44110
rect 48190 44098 48242 44110
rect 44146 44046 44158 44098
rect 44210 44046 44222 44098
rect 34638 44034 34690 44046
rect 48190 44034 48242 44046
rect 50878 44098 50930 44110
rect 50878 44034 50930 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 5070 43762 5122 43774
rect 5070 43698 5122 43710
rect 5854 43762 5906 43774
rect 5854 43698 5906 43710
rect 12910 43762 12962 43774
rect 12910 43698 12962 43710
rect 19294 43762 19346 43774
rect 19294 43698 19346 43710
rect 22430 43762 22482 43774
rect 22430 43698 22482 43710
rect 23662 43762 23714 43774
rect 23662 43698 23714 43710
rect 26798 43762 26850 43774
rect 26798 43698 26850 43710
rect 39790 43762 39842 43774
rect 39790 43698 39842 43710
rect 41358 43762 41410 43774
rect 41358 43698 41410 43710
rect 46174 43762 46226 43774
rect 46174 43698 46226 43710
rect 4958 43650 5010 43662
rect 2482 43598 2494 43650
rect 2546 43598 2558 43650
rect 4958 43586 5010 43598
rect 10222 43650 10274 43662
rect 10222 43586 10274 43598
rect 10334 43650 10386 43662
rect 10334 43586 10386 43598
rect 10894 43650 10946 43662
rect 10894 43586 10946 43598
rect 11118 43650 11170 43662
rect 11118 43586 11170 43598
rect 11230 43650 11282 43662
rect 11230 43586 11282 43598
rect 12798 43650 12850 43662
rect 12798 43586 12850 43598
rect 13806 43650 13858 43662
rect 16382 43650 16434 43662
rect 15362 43598 15374 43650
rect 15426 43598 15438 43650
rect 13806 43586 13858 43598
rect 16382 43586 16434 43598
rect 17726 43650 17778 43662
rect 17726 43586 17778 43598
rect 18846 43650 18898 43662
rect 18846 43586 18898 43598
rect 20638 43650 20690 43662
rect 20638 43586 20690 43598
rect 24222 43650 24274 43662
rect 24222 43586 24274 43598
rect 24670 43650 24722 43662
rect 24670 43586 24722 43598
rect 25342 43650 25394 43662
rect 25342 43586 25394 43598
rect 27022 43650 27074 43662
rect 34414 43650 34466 43662
rect 29586 43598 29598 43650
rect 29650 43598 29662 43650
rect 33394 43598 33406 43650
rect 33458 43598 33470 43650
rect 27022 43586 27074 43598
rect 34414 43586 34466 43598
rect 34638 43650 34690 43662
rect 34638 43586 34690 43598
rect 38558 43650 38610 43662
rect 38558 43586 38610 43598
rect 39118 43650 39170 43662
rect 39118 43586 39170 43598
rect 39230 43650 39282 43662
rect 39230 43586 39282 43598
rect 39566 43650 39618 43662
rect 39566 43586 39618 43598
rect 40350 43650 40402 43662
rect 40350 43586 40402 43598
rect 41918 43650 41970 43662
rect 41918 43586 41970 43598
rect 42366 43650 42418 43662
rect 42366 43586 42418 43598
rect 46846 43650 46898 43662
rect 46846 43586 46898 43598
rect 50094 43650 50146 43662
rect 50418 43598 50430 43650
rect 50482 43598 50494 43650
rect 50094 43586 50146 43598
rect 5518 43538 5570 43550
rect 1810 43486 1822 43538
rect 1874 43486 1886 43538
rect 5518 43474 5570 43486
rect 5742 43538 5794 43550
rect 11454 43538 11506 43550
rect 6626 43486 6638 43538
rect 6690 43486 6702 43538
rect 5742 43474 5794 43486
rect 11454 43474 11506 43486
rect 11790 43538 11842 43550
rect 11790 43474 11842 43486
rect 12014 43538 12066 43550
rect 12686 43538 12738 43550
rect 12226 43486 12238 43538
rect 12290 43486 12302 43538
rect 12014 43474 12066 43486
rect 12686 43474 12738 43486
rect 13134 43538 13186 43550
rect 13134 43474 13186 43486
rect 13358 43538 13410 43550
rect 13358 43474 13410 43486
rect 13694 43538 13746 43550
rect 13694 43474 13746 43486
rect 13918 43538 13970 43550
rect 13918 43474 13970 43486
rect 14366 43538 14418 43550
rect 16270 43538 16322 43550
rect 16942 43538 16994 43550
rect 15138 43486 15150 43538
rect 15202 43486 15214 43538
rect 16594 43486 16606 43538
rect 16658 43486 16670 43538
rect 14366 43474 14418 43486
rect 16270 43474 16322 43486
rect 16942 43474 16994 43486
rect 18174 43538 18226 43550
rect 18174 43474 18226 43486
rect 18398 43538 18450 43550
rect 21534 43538 21586 43550
rect 19506 43486 19518 43538
rect 19570 43486 19582 43538
rect 18398 43474 18450 43486
rect 21534 43474 21586 43486
rect 21870 43538 21922 43550
rect 23550 43538 23602 43550
rect 23202 43486 23214 43538
rect 23266 43486 23278 43538
rect 21870 43474 21922 43486
rect 23550 43474 23602 43486
rect 23774 43538 23826 43550
rect 23774 43474 23826 43486
rect 24446 43538 24498 43550
rect 24446 43474 24498 43486
rect 25678 43538 25730 43550
rect 26462 43538 26514 43550
rect 26114 43486 26126 43538
rect 26178 43486 26190 43538
rect 25678 43474 25730 43486
rect 26462 43474 26514 43486
rect 27358 43538 27410 43550
rect 28254 43538 28306 43550
rect 27794 43486 27806 43538
rect 27858 43486 27870 43538
rect 27358 43474 27410 43486
rect 28254 43474 28306 43486
rect 28478 43538 28530 43550
rect 28478 43474 28530 43486
rect 28702 43538 28754 43550
rect 28702 43474 28754 43486
rect 28926 43538 28978 43550
rect 31054 43538 31106 43550
rect 33070 43538 33122 43550
rect 38446 43538 38498 43550
rect 29698 43486 29710 43538
rect 29762 43486 29774 43538
rect 30370 43486 30382 43538
rect 30434 43486 30446 43538
rect 31154 43486 31166 43538
rect 31218 43486 31230 43538
rect 35074 43486 35086 43538
rect 35138 43486 35150 43538
rect 28926 43474 28978 43486
rect 31054 43474 31106 43486
rect 33070 43474 33122 43486
rect 38446 43474 38498 43486
rect 38782 43538 38834 43550
rect 38782 43474 38834 43486
rect 38894 43538 38946 43550
rect 38894 43474 38946 43486
rect 40798 43538 40850 43550
rect 40798 43474 40850 43486
rect 41246 43538 41298 43550
rect 41246 43474 41298 43486
rect 41470 43538 41522 43550
rect 41470 43474 41522 43486
rect 42142 43538 42194 43550
rect 45278 43538 45330 43550
rect 49646 43538 49698 43550
rect 44818 43486 44830 43538
rect 44882 43486 44894 43538
rect 49074 43486 49086 43538
rect 49138 43486 49150 43538
rect 42142 43474 42194 43486
rect 45278 43474 45330 43486
rect 49646 43474 49698 43486
rect 9886 43426 9938 43438
rect 4610 43374 4622 43426
rect 4674 43374 4686 43426
rect 7410 43374 7422 43426
rect 7474 43374 7486 43426
rect 9886 43362 9938 43374
rect 14814 43426 14866 43438
rect 14814 43362 14866 43374
rect 16158 43426 16210 43438
rect 16158 43362 16210 43374
rect 17502 43426 17554 43438
rect 17502 43362 17554 43374
rect 24558 43426 24610 43438
rect 24558 43362 24610 43374
rect 27134 43426 27186 43438
rect 42254 43426 42306 43438
rect 30482 43374 30494 43426
rect 30546 43374 30558 43426
rect 34738 43374 34750 43426
rect 34802 43374 34814 43426
rect 35858 43374 35870 43426
rect 35922 43374 35934 43426
rect 37986 43374 37998 43426
rect 38050 43374 38062 43426
rect 39890 43374 39902 43426
rect 39954 43374 39966 43426
rect 27134 43362 27186 43374
rect 42254 43362 42306 43374
rect 45390 43426 45442 43438
rect 45390 43362 45442 43374
rect 46174 43426 46226 43438
rect 46174 43362 46226 43374
rect 47294 43426 47346 43438
rect 47294 43362 47346 43374
rect 49758 43426 49810 43438
rect 49758 43362 49810 43374
rect 51102 43426 51154 43438
rect 51102 43362 51154 43374
rect 5854 43314 5906 43326
rect 5854 43250 5906 43262
rect 10222 43314 10274 43326
rect 10222 43250 10274 43262
rect 11678 43314 11730 43326
rect 11678 43250 11730 43262
rect 18622 43314 18674 43326
rect 18622 43250 18674 43262
rect 19182 43314 19234 43326
rect 19182 43250 19234 43262
rect 28814 43314 28866 43326
rect 28814 43250 28866 43262
rect 45838 43314 45890 43326
rect 45838 43250 45890 43262
rect 46062 43314 46114 43326
rect 46062 43250 46114 43262
rect 51326 43314 51378 43326
rect 51326 43250 51378 43262
rect 51662 43314 51714 43326
rect 51662 43250 51714 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 3726 42978 3778 42990
rect 3378 42926 3390 42978
rect 3442 42926 3454 42978
rect 3726 42914 3778 42926
rect 7198 42978 7250 42990
rect 11678 42978 11730 42990
rect 7522 42926 7534 42978
rect 7586 42926 7598 42978
rect 7198 42914 7250 42926
rect 11678 42914 11730 42926
rect 12910 42978 12962 42990
rect 12910 42914 12962 42926
rect 16046 42978 16098 42990
rect 16046 42914 16098 42926
rect 18846 42978 18898 42990
rect 18846 42914 18898 42926
rect 22654 42978 22706 42990
rect 22654 42914 22706 42926
rect 30046 42978 30098 42990
rect 30046 42914 30098 42926
rect 34526 42978 34578 42990
rect 45266 42926 45278 42978
rect 45330 42975 45342 42978
rect 45826 42975 45838 42978
rect 45330 42929 45838 42975
rect 45330 42926 45342 42929
rect 45826 42926 45838 42929
rect 45890 42926 45902 42978
rect 34526 42914 34578 42926
rect 3950 42866 4002 42878
rect 3950 42802 4002 42814
rect 4734 42866 4786 42878
rect 11454 42866 11506 42878
rect 6514 42814 6526 42866
rect 6578 42814 6590 42866
rect 8642 42814 8654 42866
rect 8706 42814 8718 42866
rect 10770 42814 10782 42866
rect 10834 42814 10846 42866
rect 4734 42802 4786 42814
rect 11454 42802 11506 42814
rect 14702 42866 14754 42878
rect 17054 42866 17106 42878
rect 15810 42814 15822 42866
rect 15874 42814 15886 42866
rect 14702 42802 14754 42814
rect 17054 42802 17106 42814
rect 20526 42866 20578 42878
rect 25566 42866 25618 42878
rect 23538 42814 23550 42866
rect 23602 42814 23614 42866
rect 20526 42802 20578 42814
rect 25566 42802 25618 42814
rect 26350 42866 26402 42878
rect 26350 42802 26402 42814
rect 27582 42866 27634 42878
rect 27582 42802 27634 42814
rect 29150 42866 29202 42878
rect 42142 42866 42194 42878
rect 29474 42814 29486 42866
rect 29538 42814 29550 42866
rect 30930 42814 30942 42866
rect 30994 42814 31006 42866
rect 36082 42814 36094 42866
rect 36146 42814 36158 42866
rect 39890 42814 39902 42866
rect 39954 42814 39966 42866
rect 29150 42802 29202 42814
rect 42142 42802 42194 42814
rect 45838 42866 45890 42878
rect 50194 42814 50206 42866
rect 50258 42814 50270 42866
rect 45838 42802 45890 42814
rect 6974 42754 7026 42766
rect 12798 42754 12850 42766
rect 5842 42702 5854 42754
rect 5906 42702 5918 42754
rect 6626 42702 6638 42754
rect 6690 42702 6702 42754
rect 7858 42702 7870 42754
rect 7922 42702 7934 42754
rect 6974 42690 7026 42702
rect 12798 42690 12850 42702
rect 13358 42754 13410 42766
rect 13918 42754 13970 42766
rect 13682 42702 13694 42754
rect 13746 42702 13758 42754
rect 13358 42690 13410 42702
rect 13918 42690 13970 42702
rect 14142 42754 14194 42766
rect 14142 42690 14194 42702
rect 15598 42754 15650 42766
rect 15598 42690 15650 42702
rect 16270 42754 16322 42766
rect 16270 42690 16322 42702
rect 16942 42754 16994 42766
rect 16942 42690 16994 42702
rect 17726 42754 17778 42766
rect 22318 42754 22370 42766
rect 25454 42754 25506 42766
rect 19394 42702 19406 42754
rect 19458 42702 19470 42754
rect 19842 42702 19854 42754
rect 19906 42702 19918 42754
rect 22978 42702 22990 42754
rect 23042 42702 23054 42754
rect 24882 42702 24894 42754
rect 24946 42702 24958 42754
rect 17726 42690 17778 42702
rect 22318 42690 22370 42702
rect 25454 42690 25506 42702
rect 26462 42754 26514 42766
rect 26462 42690 26514 42702
rect 26798 42754 26850 42766
rect 26798 42690 26850 42702
rect 28254 42754 28306 42766
rect 28254 42690 28306 42702
rect 28590 42754 28642 42766
rect 28590 42690 28642 42702
rect 29934 42754 29986 42766
rect 30830 42754 30882 42766
rect 30594 42702 30606 42754
rect 30658 42702 30670 42754
rect 29934 42690 29986 42702
rect 30830 42690 30882 42702
rect 34750 42754 34802 42766
rect 42366 42754 42418 42766
rect 36978 42702 36990 42754
rect 37042 42702 37054 42754
rect 40338 42702 40350 42754
rect 40402 42702 40414 42754
rect 41122 42702 41134 42754
rect 41186 42702 41198 42754
rect 41682 42702 41694 42754
rect 41746 42702 41758 42754
rect 34750 42690 34802 42702
rect 42366 42690 42418 42702
rect 46286 42754 46338 42766
rect 50542 42754 50594 42766
rect 46834 42702 46846 42754
rect 46898 42702 46910 42754
rect 47394 42702 47406 42754
rect 47458 42702 47470 42754
rect 46286 42690 46338 42702
rect 50542 42690 50594 42702
rect 50766 42754 50818 42766
rect 50766 42690 50818 42702
rect 6302 42642 6354 42654
rect 5618 42590 5630 42642
rect 5682 42590 5694 42642
rect 6302 42578 6354 42590
rect 14366 42642 14418 42654
rect 14366 42578 14418 42590
rect 14814 42642 14866 42654
rect 14814 42578 14866 42590
rect 15486 42642 15538 42654
rect 15486 42578 15538 42590
rect 17166 42642 17218 42654
rect 17166 42578 17218 42590
rect 17950 42642 18002 42654
rect 17950 42578 18002 42590
rect 18062 42642 18114 42654
rect 18062 42578 18114 42590
rect 18510 42642 18562 42654
rect 18510 42578 18562 42590
rect 18734 42642 18786 42654
rect 18734 42578 18786 42590
rect 22094 42642 22146 42654
rect 26238 42642 26290 42654
rect 28478 42642 28530 42654
rect 51438 42642 51490 42654
rect 23202 42590 23214 42642
rect 23266 42590 23278 42642
rect 27122 42590 27134 42642
rect 27186 42590 27198 42642
rect 37762 42590 37774 42642
rect 37826 42590 37838 42642
rect 41794 42590 41806 42642
rect 41858 42590 41870 42642
rect 46610 42590 46622 42642
rect 46674 42590 46686 42642
rect 48066 42590 48078 42642
rect 48130 42590 48142 42642
rect 51090 42590 51102 42642
rect 51154 42590 51166 42642
rect 22094 42578 22146 42590
rect 26238 42578 26290 42590
rect 28478 42578 28530 42590
rect 51438 42578 51490 42590
rect 51662 42642 51714 42654
rect 51662 42578 51714 42590
rect 51998 42642 52050 42654
rect 51998 42578 52050 42590
rect 5070 42530 5122 42542
rect 12686 42530 12738 42542
rect 17390 42530 17442 42542
rect 12002 42478 12014 42530
rect 12066 42478 12078 42530
rect 13794 42478 13806 42530
rect 13858 42478 13870 42530
rect 5070 42466 5122 42478
rect 12686 42466 12738 42478
rect 17390 42466 17442 42478
rect 19966 42530 20018 42542
rect 19966 42466 20018 42478
rect 26014 42530 26066 42542
rect 26014 42466 26066 42478
rect 28030 42530 28082 42542
rect 28030 42466 28082 42478
rect 29374 42530 29426 42542
rect 29374 42466 29426 42478
rect 30382 42530 30434 42542
rect 30382 42466 30434 42478
rect 31390 42530 31442 42542
rect 31390 42466 31442 42478
rect 32622 42530 32674 42542
rect 32622 42466 32674 42478
rect 34190 42530 34242 42542
rect 34190 42466 34242 42478
rect 34974 42530 35026 42542
rect 34974 42466 35026 42478
rect 35086 42530 35138 42542
rect 35086 42466 35138 42478
rect 35198 42530 35250 42542
rect 35198 42466 35250 42478
rect 35646 42530 35698 42542
rect 45390 42530 45442 42542
rect 42690 42478 42702 42530
rect 42754 42478 42766 42530
rect 35646 42466 35698 42478
rect 45390 42466 45442 42478
rect 51774 42530 51826 42542
rect 51774 42466 51826 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 14366 42194 14418 42206
rect 4386 42142 4398 42194
rect 4450 42142 4462 42194
rect 11106 42142 11118 42194
rect 11170 42142 11182 42194
rect 27470 42194 27522 42206
rect 14366 42130 14418 42142
rect 18622 42138 18674 42150
rect 14478 42082 14530 42094
rect 14478 42018 14530 42030
rect 14926 42082 14978 42094
rect 14926 42018 14978 42030
rect 17838 42082 17890 42094
rect 17838 42018 17890 42030
rect 18510 42082 18562 42094
rect 27470 42130 27522 42142
rect 28366 42194 28418 42206
rect 28366 42130 28418 42142
rect 28590 42194 28642 42206
rect 28590 42130 28642 42142
rect 29710 42194 29762 42206
rect 32286 42194 32338 42206
rect 31266 42142 31278 42194
rect 31330 42142 31342 42194
rect 29710 42130 29762 42142
rect 32286 42130 32338 42142
rect 36654 42194 36706 42206
rect 36654 42130 36706 42142
rect 37102 42194 37154 42206
rect 37102 42130 37154 42142
rect 18622 42074 18674 42086
rect 19294 42082 19346 42094
rect 18510 42018 18562 42030
rect 19294 42018 19346 42030
rect 19742 42082 19794 42094
rect 19742 42018 19794 42030
rect 19966 42082 20018 42094
rect 19966 42018 20018 42030
rect 22878 42082 22930 42094
rect 22878 42018 22930 42030
rect 27134 42082 27186 42094
rect 27134 42018 27186 42030
rect 27246 42082 27298 42094
rect 32062 42082 32114 42094
rect 30370 42030 30382 42082
rect 30434 42030 30446 42082
rect 27246 42018 27298 42030
rect 32062 42018 32114 42030
rect 33294 42082 33346 42094
rect 33294 42018 33346 42030
rect 35534 42082 35586 42094
rect 35534 42018 35586 42030
rect 36094 42082 36146 42094
rect 36094 42018 36146 42030
rect 53006 42082 53058 42094
rect 53778 42030 53790 42082
rect 53842 42030 53854 42082
rect 53006 42018 53058 42030
rect 3390 41970 3442 41982
rect 2818 41918 2830 41970
rect 2882 41918 2894 41970
rect 3390 41906 3442 41918
rect 3838 41970 3890 41982
rect 3838 41906 3890 41918
rect 4062 41970 4114 41982
rect 4062 41906 4114 41918
rect 4734 41970 4786 41982
rect 4734 41906 4786 41918
rect 4958 41970 5010 41982
rect 12238 41970 12290 41982
rect 5282 41918 5294 41970
rect 5346 41918 5358 41970
rect 8754 41918 8766 41970
rect 8818 41918 8830 41970
rect 11330 41918 11342 41970
rect 11394 41918 11406 41970
rect 4958 41906 5010 41918
rect 12238 41906 12290 41918
rect 15486 41970 15538 41982
rect 15486 41906 15538 41918
rect 16046 41970 16098 41982
rect 16046 41906 16098 41918
rect 16270 41970 16322 41982
rect 16270 41906 16322 41918
rect 16494 41970 16546 41982
rect 16494 41906 16546 41918
rect 16942 41970 16994 41982
rect 17950 41970 18002 41982
rect 20302 41970 20354 41982
rect 21982 41970 22034 41982
rect 17378 41918 17390 41970
rect 17442 41918 17454 41970
rect 18162 41918 18174 41970
rect 18226 41918 18238 41970
rect 20738 41918 20750 41970
rect 20802 41918 20814 41970
rect 21522 41918 21534 41970
rect 21586 41918 21598 41970
rect 16942 41906 16994 41918
rect 17950 41906 18002 41918
rect 20302 41906 20354 41918
rect 21982 41906 22034 41918
rect 22990 41970 23042 41982
rect 22990 41906 23042 41918
rect 23102 41970 23154 41982
rect 27806 41970 27858 41982
rect 25330 41918 25342 41970
rect 25394 41918 25406 41970
rect 26002 41918 26014 41970
rect 26066 41918 26078 41970
rect 26450 41918 26462 41970
rect 26514 41918 26526 41970
rect 23102 41906 23154 41918
rect 27806 41906 27858 41918
rect 28142 41970 28194 41982
rect 28142 41906 28194 41918
rect 28814 41970 28866 41982
rect 28814 41906 28866 41918
rect 29038 41970 29090 41982
rect 29038 41906 29090 41918
rect 29486 41970 29538 41982
rect 29486 41906 29538 41918
rect 30046 41970 30098 41982
rect 30046 41906 30098 41918
rect 30942 41970 30994 41982
rect 30942 41906 30994 41918
rect 31614 41970 31666 41982
rect 35310 41970 35362 41982
rect 34962 41918 34974 41970
rect 35026 41918 35038 41970
rect 31614 41906 31666 41918
rect 35310 41906 35362 41918
rect 35870 41970 35922 41982
rect 38894 41970 38946 41982
rect 40126 41970 40178 41982
rect 38658 41918 38670 41970
rect 38722 41918 38734 41970
rect 39778 41918 39790 41970
rect 39842 41918 39854 41970
rect 42242 41918 42254 41970
rect 42306 41918 42318 41970
rect 43250 41918 43262 41970
rect 43314 41918 43326 41970
rect 44034 41918 44046 41970
rect 44098 41918 44110 41970
rect 45378 41918 45390 41970
rect 45442 41918 45454 41970
rect 49410 41918 49422 41970
rect 49474 41918 49486 41970
rect 49746 41918 49758 41970
rect 49810 41918 49822 41970
rect 51762 41918 51774 41970
rect 51826 41918 51838 41970
rect 52770 41918 52782 41970
rect 52834 41918 52846 41970
rect 53666 41918 53678 41970
rect 53730 41918 53742 41970
rect 35870 41906 35922 41918
rect 38894 41906 38946 41918
rect 40126 41906 40178 41918
rect 3166 41858 3218 41870
rect 3166 41794 3218 41806
rect 3950 41858 4002 41870
rect 3950 41794 4002 41806
rect 5854 41858 5906 41870
rect 9662 41858 9714 41870
rect 7634 41806 7646 41858
rect 7698 41806 7710 41858
rect 5854 41794 5906 41806
rect 9662 41794 9714 41806
rect 13918 41858 13970 41870
rect 13918 41794 13970 41806
rect 16382 41858 16434 41870
rect 27694 41858 27746 41870
rect 19394 41806 19406 41858
rect 19458 41806 19470 41858
rect 19954 41806 19966 41858
rect 20018 41806 20030 41858
rect 16382 41794 16434 41806
rect 27694 41794 27746 41806
rect 29598 41858 29650 41870
rect 29598 41794 29650 41806
rect 31838 41858 31890 41870
rect 31838 41794 31890 41806
rect 32174 41858 32226 41870
rect 32174 41794 32226 41806
rect 33182 41858 33234 41870
rect 33182 41794 33234 41806
rect 35422 41858 35474 41870
rect 38334 41858 38386 41870
rect 36194 41806 36206 41858
rect 36258 41806 36270 41858
rect 45602 41806 45614 41858
rect 45666 41806 45678 41858
rect 48850 41806 48862 41858
rect 48914 41806 48926 41858
rect 50754 41806 50766 41858
rect 50818 41806 50830 41858
rect 51650 41806 51662 41858
rect 51714 41806 51726 41858
rect 53554 41806 53566 41858
rect 53618 41806 53630 41858
rect 35422 41794 35474 41806
rect 38334 41794 38386 41806
rect 2830 41746 2882 41758
rect 2830 41682 2882 41694
rect 5630 41746 5682 41758
rect 5630 41682 5682 41694
rect 14366 41746 14418 41758
rect 14366 41682 14418 41694
rect 14814 41746 14866 41758
rect 14814 41682 14866 41694
rect 18622 41746 18674 41758
rect 18622 41682 18674 41694
rect 19070 41746 19122 41758
rect 19070 41682 19122 41694
rect 20750 41746 20802 41758
rect 20750 41682 20802 41694
rect 21086 41746 21138 41758
rect 28702 41746 28754 41758
rect 23538 41694 23550 41746
rect 23602 41694 23614 41746
rect 26226 41694 26238 41746
rect 26290 41694 26302 41746
rect 21086 41682 21138 41694
rect 28702 41682 28754 41694
rect 33070 41746 33122 41758
rect 33070 41682 33122 41694
rect 39118 41746 39170 41758
rect 39118 41682 39170 41694
rect 39342 41746 39394 41758
rect 39342 41682 39394 41694
rect 39454 41746 39506 41758
rect 39454 41682 39506 41694
rect 39790 41746 39842 41758
rect 46050 41694 46062 41746
rect 46114 41694 46126 41746
rect 39790 41682 39842 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 6414 41410 6466 41422
rect 6414 41346 6466 41358
rect 6862 41410 6914 41422
rect 6862 41346 6914 41358
rect 13470 41410 13522 41422
rect 13470 41346 13522 41358
rect 13582 41410 13634 41422
rect 13582 41346 13634 41358
rect 15262 41410 15314 41422
rect 15262 41346 15314 41358
rect 18286 41410 18338 41422
rect 18286 41346 18338 41358
rect 18622 41410 18674 41422
rect 18622 41346 18674 41358
rect 19966 41410 20018 41422
rect 19966 41346 20018 41358
rect 20302 41410 20354 41422
rect 20302 41346 20354 41358
rect 22542 41410 22594 41422
rect 22542 41346 22594 41358
rect 25342 41410 25394 41422
rect 49982 41410 50034 41422
rect 27570 41358 27582 41410
rect 27634 41358 27646 41410
rect 51762 41358 51774 41410
rect 51826 41358 51838 41410
rect 25342 41346 25394 41358
rect 49982 41346 50034 41358
rect 5070 41298 5122 41310
rect 2482 41246 2494 41298
rect 2546 41246 2558 41298
rect 4610 41246 4622 41298
rect 4674 41246 4686 41298
rect 5070 41234 5122 41246
rect 7758 41298 7810 41310
rect 11902 41298 11954 41310
rect 8866 41246 8878 41298
rect 8930 41246 8942 41298
rect 10994 41246 11006 41298
rect 11058 41246 11070 41298
rect 7758 41234 7810 41246
rect 11902 41234 11954 41246
rect 14254 41298 14306 41310
rect 16158 41298 16210 41310
rect 14466 41246 14478 41298
rect 14530 41295 14542 41298
rect 14802 41295 14814 41298
rect 14530 41249 14814 41295
rect 14530 41246 14542 41249
rect 14802 41246 14814 41249
rect 14866 41246 14878 41298
rect 14254 41234 14306 41246
rect 16158 41234 16210 41246
rect 16606 41298 16658 41310
rect 16606 41234 16658 41246
rect 19630 41298 19682 41310
rect 19630 41234 19682 41246
rect 23326 41298 23378 41310
rect 36206 41298 36258 41310
rect 48862 41298 48914 41310
rect 32722 41246 32734 41298
rect 32786 41246 32798 41298
rect 34850 41246 34862 41298
rect 34914 41246 34926 41298
rect 43026 41246 43038 41298
rect 43090 41246 43102 41298
rect 44818 41246 44830 41298
rect 44882 41246 44894 41298
rect 23326 41234 23378 41246
rect 36206 41234 36258 41246
rect 48862 41234 48914 41246
rect 6190 41186 6242 41198
rect 1810 41134 1822 41186
rect 1874 41134 1886 41186
rect 5954 41134 5966 41186
rect 6018 41134 6030 41186
rect 6190 41122 6242 41134
rect 6974 41186 7026 41198
rect 12238 41186 12290 41198
rect 8082 41134 8094 41186
rect 8146 41134 8158 41186
rect 6974 41122 7026 41134
rect 12238 41122 12290 41134
rect 13694 41186 13746 41198
rect 13694 41122 13746 41134
rect 14030 41186 14082 41198
rect 14030 41122 14082 41134
rect 15038 41186 15090 41198
rect 15038 41122 15090 41134
rect 17390 41186 17442 41198
rect 17390 41122 17442 41134
rect 17726 41186 17778 41198
rect 17726 41122 17778 41134
rect 17950 41186 18002 41198
rect 19742 41186 19794 41198
rect 18274 41134 18286 41186
rect 18338 41134 18350 41186
rect 17950 41122 18002 41134
rect 19742 41122 19794 41134
rect 20190 41186 20242 41198
rect 22654 41186 22706 41198
rect 21410 41134 21422 41186
rect 21474 41134 21486 41186
rect 21970 41134 21982 41186
rect 22034 41134 22046 41186
rect 22194 41134 22206 41186
rect 22258 41134 22270 41186
rect 20190 41122 20242 41134
rect 22654 41122 22706 41134
rect 25454 41186 25506 41198
rect 25454 41122 25506 41134
rect 25790 41186 25842 41198
rect 27134 41186 27186 41198
rect 35310 41186 35362 41198
rect 26226 41134 26238 41186
rect 26290 41134 26302 41186
rect 26786 41134 26798 41186
rect 26850 41134 26862 41186
rect 27682 41134 27694 41186
rect 27746 41134 27758 41186
rect 29922 41134 29934 41186
rect 29986 41134 29998 41186
rect 32050 41134 32062 41186
rect 32114 41134 32126 41186
rect 25790 41122 25842 41134
rect 27134 41122 27186 41134
rect 35310 41122 35362 41134
rect 35758 41186 35810 41198
rect 35758 41122 35810 41134
rect 36990 41186 37042 41198
rect 39566 41186 39618 41198
rect 51214 41186 51266 41198
rect 37538 41134 37550 41186
rect 37602 41134 37614 41186
rect 42018 41134 42030 41186
rect 42082 41134 42094 41186
rect 42802 41134 42814 41186
rect 42866 41134 42878 41186
rect 43810 41134 43822 41186
rect 43874 41134 43886 41186
rect 47730 41134 47742 41186
rect 47794 41134 47806 41186
rect 50978 41134 50990 41186
rect 51042 41134 51054 41186
rect 36990 41122 37042 41134
rect 39566 41122 39618 41134
rect 51214 41122 51266 41134
rect 51326 41186 51378 41198
rect 51326 41122 51378 41134
rect 6526 41074 6578 41086
rect 6526 41010 6578 41022
rect 7086 41074 7138 41086
rect 7086 41010 7138 41022
rect 19182 41074 19234 41086
rect 19182 41010 19234 41022
rect 19294 41074 19346 41086
rect 19294 41010 19346 41022
rect 22430 41074 22482 41086
rect 22430 41010 22482 41022
rect 22990 41074 23042 41086
rect 22990 41010 23042 41022
rect 23438 41074 23490 41086
rect 23438 41010 23490 41022
rect 29486 41074 29538 41086
rect 35422 41074 35474 41086
rect 30594 41022 30606 41074
rect 30658 41022 30670 41074
rect 29486 41010 29538 41022
rect 35422 41010 35474 41022
rect 37214 41074 37266 41086
rect 37214 41010 37266 41022
rect 39678 41074 39730 41086
rect 39678 41010 39730 41022
rect 41582 41074 41634 41086
rect 44270 41074 44322 41086
rect 49982 41074 50034 41086
rect 42466 41022 42478 41074
rect 42530 41022 42542 41074
rect 46946 41022 46958 41074
rect 47010 41022 47022 41074
rect 41582 41010 41634 41022
rect 44270 41010 44322 41022
rect 49982 41010 50034 41022
rect 50094 41074 50146 41086
rect 50094 41010 50146 41022
rect 50430 41074 50482 41086
rect 50430 41010 50482 41022
rect 50542 41074 50594 41086
rect 50542 41010 50594 41022
rect 16046 40962 16098 40974
rect 12562 40910 12574 40962
rect 12626 40910 12638 40962
rect 15586 40910 15598 40962
rect 15650 40910 15662 40962
rect 16046 40898 16098 40910
rect 17054 40962 17106 40974
rect 17054 40898 17106 40910
rect 17614 40962 17666 40974
rect 17614 40898 17666 40910
rect 19070 40962 19122 40974
rect 22878 40962 22930 40974
rect 21634 40910 21646 40962
rect 21698 40910 21710 40962
rect 19070 40898 19122 40910
rect 22878 40898 22930 40910
rect 25342 40962 25394 40974
rect 25342 40898 25394 40910
rect 29150 40962 29202 40974
rect 29150 40898 29202 40910
rect 29262 40962 29314 40974
rect 29262 40898 29314 40910
rect 29374 40962 29426 40974
rect 29374 40898 29426 40910
rect 30270 40962 30322 40974
rect 30270 40898 30322 40910
rect 35646 40962 35698 40974
rect 35646 40898 35698 40910
rect 37102 40962 37154 40974
rect 37102 40898 37154 40910
rect 38110 40962 38162 40974
rect 39230 40962 39282 40974
rect 38882 40910 38894 40962
rect 38946 40910 38958 40962
rect 38110 40898 38162 40910
rect 39230 40898 39282 40910
rect 39902 40962 39954 40974
rect 39902 40898 39954 40910
rect 41470 40962 41522 40974
rect 41470 40898 41522 40910
rect 41694 40962 41746 40974
rect 44158 40962 44210 40974
rect 43698 40910 43710 40962
rect 43762 40910 43774 40962
rect 41694 40898 41746 40910
rect 44158 40898 44210 40910
rect 48190 40962 48242 40974
rect 48190 40898 48242 40910
rect 49422 40962 49474 40974
rect 49422 40898 49474 40910
rect 50766 40962 50818 40974
rect 50766 40898 50818 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 4510 40626 4562 40638
rect 4510 40562 4562 40574
rect 8990 40626 9042 40638
rect 8990 40562 9042 40574
rect 13918 40626 13970 40638
rect 13918 40562 13970 40574
rect 14478 40626 14530 40638
rect 14478 40562 14530 40574
rect 14590 40626 14642 40638
rect 16382 40626 16434 40638
rect 15698 40574 15710 40626
rect 15762 40574 15774 40626
rect 14590 40562 14642 40574
rect 16382 40562 16434 40574
rect 22094 40626 22146 40638
rect 22094 40562 22146 40574
rect 24670 40626 24722 40638
rect 24670 40562 24722 40574
rect 28702 40626 28754 40638
rect 28702 40562 28754 40574
rect 29710 40626 29762 40638
rect 38446 40626 38498 40638
rect 32274 40574 32286 40626
rect 32338 40574 32350 40626
rect 29710 40562 29762 40574
rect 38446 40562 38498 40574
rect 44382 40626 44434 40638
rect 44382 40562 44434 40574
rect 45278 40626 45330 40638
rect 45278 40562 45330 40574
rect 45950 40626 46002 40638
rect 45950 40562 46002 40574
rect 46846 40626 46898 40638
rect 46846 40562 46898 40574
rect 47182 40626 47234 40638
rect 47182 40562 47234 40574
rect 48974 40626 49026 40638
rect 48974 40562 49026 40574
rect 49198 40626 49250 40638
rect 49198 40562 49250 40574
rect 51438 40626 51490 40638
rect 51438 40562 51490 40574
rect 51662 40626 51714 40638
rect 51662 40562 51714 40574
rect 51998 40626 52050 40638
rect 51998 40562 52050 40574
rect 52222 40626 52274 40638
rect 52222 40562 52274 40574
rect 52558 40626 52610 40638
rect 52558 40562 52610 40574
rect 16046 40514 16098 40526
rect 7746 40462 7758 40514
rect 7810 40462 7822 40514
rect 10322 40462 10334 40514
rect 10386 40462 10398 40514
rect 13122 40462 13134 40514
rect 13186 40462 13198 40514
rect 16046 40450 16098 40462
rect 16158 40514 16210 40526
rect 16158 40450 16210 40462
rect 16718 40514 16770 40526
rect 16718 40450 16770 40462
rect 16830 40514 16882 40526
rect 16830 40450 16882 40462
rect 22318 40514 22370 40526
rect 22318 40450 22370 40462
rect 22430 40514 22482 40526
rect 22430 40450 22482 40462
rect 24558 40514 24610 40526
rect 26798 40514 26850 40526
rect 26226 40462 26238 40514
rect 26290 40462 26302 40514
rect 24558 40450 24610 40462
rect 26798 40450 26850 40462
rect 26910 40514 26962 40526
rect 26910 40450 26962 40462
rect 27358 40514 27410 40526
rect 27358 40450 27410 40462
rect 27470 40514 27522 40526
rect 38222 40514 38274 40526
rect 50990 40514 51042 40526
rect 28354 40462 28366 40514
rect 28418 40462 28430 40514
rect 29026 40462 29038 40514
rect 29090 40462 29102 40514
rect 30930 40462 30942 40514
rect 30994 40462 31006 40514
rect 32498 40462 32510 40514
rect 32562 40462 32574 40514
rect 35746 40462 35758 40514
rect 35810 40462 35822 40514
rect 39778 40462 39790 40514
rect 39842 40462 39854 40514
rect 45602 40462 45614 40514
rect 45666 40462 45678 40514
rect 46274 40462 46286 40514
rect 46338 40462 46350 40514
rect 27470 40450 27522 40462
rect 38222 40450 38274 40462
rect 50990 40450 51042 40462
rect 51326 40514 51378 40526
rect 51326 40450 51378 40462
rect 51886 40514 51938 40526
rect 51886 40450 51938 40462
rect 12798 40402 12850 40414
rect 14702 40402 14754 40414
rect 16494 40402 16546 40414
rect 8418 40350 8430 40402
rect 8482 40350 8494 40402
rect 9538 40350 9550 40402
rect 9602 40350 9614 40402
rect 13906 40350 13918 40402
rect 13970 40350 13982 40402
rect 15026 40350 15038 40402
rect 15090 40350 15102 40402
rect 15474 40350 15486 40402
rect 15538 40350 15550 40402
rect 12798 40338 12850 40350
rect 14702 40338 14754 40350
rect 16494 40338 16546 40350
rect 17502 40402 17554 40414
rect 17502 40338 17554 40350
rect 18734 40402 18786 40414
rect 18734 40338 18786 40350
rect 19630 40402 19682 40414
rect 19630 40338 19682 40350
rect 19966 40402 20018 40414
rect 19966 40338 20018 40350
rect 20414 40402 20466 40414
rect 20414 40338 20466 40350
rect 21198 40402 21250 40414
rect 21198 40338 21250 40350
rect 21646 40402 21698 40414
rect 21646 40338 21698 40350
rect 21870 40402 21922 40414
rect 29934 40402 29986 40414
rect 31950 40402 32002 40414
rect 39006 40402 39058 40414
rect 41918 40402 41970 40414
rect 25218 40350 25230 40402
rect 25282 40350 25294 40402
rect 26002 40350 26014 40402
rect 26066 40350 26078 40402
rect 28130 40350 28142 40402
rect 28194 40350 28206 40402
rect 29362 40350 29374 40402
rect 29426 40350 29438 40402
rect 30818 40350 30830 40402
rect 30882 40350 30894 40402
rect 35074 40350 35086 40402
rect 35138 40350 35150 40402
rect 40002 40350 40014 40402
rect 40066 40350 40078 40402
rect 41346 40350 41358 40402
rect 41410 40350 41422 40402
rect 21870 40338 21922 40350
rect 29934 40338 29986 40350
rect 31950 40338 32002 40350
rect 39006 40338 39058 40350
rect 41918 40338 41970 40350
rect 42254 40402 42306 40414
rect 42254 40338 42306 40350
rect 42590 40402 42642 40414
rect 42590 40338 42642 40350
rect 42926 40402 42978 40414
rect 43598 40402 43650 40414
rect 43250 40350 43262 40402
rect 43314 40350 43326 40402
rect 42926 40338 42978 40350
rect 43598 40338 43650 40350
rect 43822 40402 43874 40414
rect 43822 40338 43874 40350
rect 44942 40402 44994 40414
rect 44942 40338 44994 40350
rect 48190 40402 48242 40414
rect 49534 40402 49586 40414
rect 48738 40350 48750 40402
rect 48802 40350 48814 40402
rect 48190 40338 48242 40350
rect 49534 40338 49586 40350
rect 49758 40402 49810 40414
rect 49758 40338 49810 40350
rect 50094 40402 50146 40414
rect 50094 40338 50146 40350
rect 50318 40402 50370 40414
rect 50318 40338 50370 40350
rect 50766 40402 50818 40414
rect 50766 40338 50818 40350
rect 4622 40290 4674 40302
rect 4622 40226 4674 40238
rect 4846 40290 4898 40302
rect 18062 40290 18114 40302
rect 5618 40238 5630 40290
rect 5682 40238 5694 40290
rect 12450 40238 12462 40290
rect 12514 40238 12526 40290
rect 4846 40226 4898 40238
rect 18062 40226 18114 40238
rect 18510 40290 18562 40302
rect 18510 40226 18562 40238
rect 21758 40290 21810 40302
rect 29822 40290 29874 40302
rect 38334 40290 38386 40302
rect 25666 40238 25678 40290
rect 25730 40238 25742 40290
rect 37874 40238 37886 40290
rect 37938 40238 37950 40290
rect 21758 40226 21810 40238
rect 29822 40226 29874 40238
rect 38334 40226 38386 40238
rect 42030 40290 42082 40302
rect 42030 40226 42082 40238
rect 42478 40290 42530 40302
rect 42478 40226 42530 40238
rect 47742 40290 47794 40302
rect 49646 40290 49698 40302
rect 49186 40238 49198 40290
rect 49250 40238 49262 40290
rect 47742 40226 47794 40238
rect 49646 40226 49698 40238
rect 50878 40290 50930 40302
rect 50878 40226 50930 40238
rect 4510 40178 4562 40190
rect 4510 40114 4562 40126
rect 18286 40178 18338 40190
rect 18286 40114 18338 40126
rect 19182 40178 19234 40190
rect 19182 40114 19234 40126
rect 26910 40178 26962 40190
rect 26910 40114 26962 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 6190 39842 6242 39854
rect 6190 39778 6242 39790
rect 15374 39842 15426 39854
rect 15374 39778 15426 39790
rect 15822 39842 15874 39854
rect 15822 39778 15874 39790
rect 26686 39842 26738 39854
rect 28590 39842 28642 39854
rect 27234 39790 27246 39842
rect 27298 39790 27310 39842
rect 26686 39778 26738 39790
rect 28590 39778 28642 39790
rect 29934 39842 29986 39854
rect 29934 39778 29986 39790
rect 5070 39730 5122 39742
rect 5070 39666 5122 39678
rect 8766 39730 8818 39742
rect 8766 39666 8818 39678
rect 11454 39730 11506 39742
rect 20750 39730 20802 39742
rect 30046 39730 30098 39742
rect 12674 39678 12686 39730
rect 12738 39678 12750 39730
rect 16146 39678 16158 39730
rect 16210 39678 16222 39730
rect 18050 39678 18062 39730
rect 18114 39678 18126 39730
rect 23538 39678 23550 39730
rect 23602 39678 23614 39730
rect 25106 39678 25118 39730
rect 25170 39678 25182 39730
rect 11454 39666 11506 39678
rect 20750 39666 20802 39678
rect 30046 39666 30098 39678
rect 36430 39730 36482 39742
rect 41918 39730 41970 39742
rect 48862 39730 48914 39742
rect 37762 39678 37774 39730
rect 37826 39678 37838 39730
rect 39890 39678 39902 39730
rect 39954 39678 39966 39730
rect 42466 39678 42478 39730
rect 42530 39678 42542 39730
rect 36430 39666 36482 39678
rect 41918 39666 41970 39678
rect 48862 39666 48914 39678
rect 4734 39618 4786 39630
rect 4734 39554 4786 39566
rect 5518 39618 5570 39630
rect 15486 39618 15538 39630
rect 19630 39618 19682 39630
rect 12226 39566 12238 39618
rect 12290 39566 12302 39618
rect 12562 39566 12574 39618
rect 12626 39566 12638 39618
rect 17826 39566 17838 39618
rect 17890 39566 17902 39618
rect 5518 39554 5570 39566
rect 15486 39554 15538 39566
rect 19630 39554 19682 39566
rect 21310 39618 21362 39630
rect 21310 39554 21362 39566
rect 21870 39618 21922 39630
rect 21870 39554 21922 39566
rect 22430 39618 22482 39630
rect 25342 39618 25394 39630
rect 24994 39566 25006 39618
rect 25058 39566 25070 39618
rect 22430 39554 22482 39566
rect 25342 39554 25394 39566
rect 25678 39618 25730 39630
rect 25678 39554 25730 39566
rect 26574 39618 26626 39630
rect 27918 39618 27970 39630
rect 29038 39618 29090 39630
rect 27682 39566 27694 39618
rect 27746 39566 27758 39618
rect 28578 39566 28590 39618
rect 28642 39566 28654 39618
rect 26574 39554 26626 39566
rect 27918 39554 27970 39566
rect 29038 39554 29090 39566
rect 32510 39618 32562 39630
rect 32510 39554 32562 39566
rect 33406 39618 33458 39630
rect 44830 39618 44882 39630
rect 37090 39566 37102 39618
rect 37154 39566 37166 39618
rect 41234 39566 41246 39618
rect 41298 39566 41310 39618
rect 41682 39566 41694 39618
rect 41746 39566 41758 39618
rect 42690 39566 42702 39618
rect 42754 39566 42766 39618
rect 33406 39554 33458 39566
rect 44830 39554 44882 39566
rect 45390 39618 45442 39630
rect 45390 39554 45442 39566
rect 46286 39618 46338 39630
rect 46286 39554 46338 39566
rect 47182 39618 47234 39630
rect 47182 39554 47234 39566
rect 47518 39618 47570 39630
rect 48414 39618 48466 39630
rect 47954 39566 47966 39618
rect 48018 39566 48030 39618
rect 47518 39554 47570 39566
rect 48414 39554 48466 39566
rect 48638 39618 48690 39630
rect 48638 39554 48690 39566
rect 49310 39618 49362 39630
rect 49310 39554 49362 39566
rect 49758 39618 49810 39630
rect 49758 39554 49810 39566
rect 49870 39618 49922 39630
rect 49870 39554 49922 39566
rect 50318 39618 50370 39630
rect 50318 39554 50370 39566
rect 50654 39618 50706 39630
rect 50654 39554 50706 39566
rect 13022 39506 13074 39518
rect 13022 39442 13074 39454
rect 14590 39506 14642 39518
rect 14590 39442 14642 39454
rect 14926 39506 14978 39518
rect 28254 39506 28306 39518
rect 17042 39454 17054 39506
rect 17106 39454 17118 39506
rect 18274 39454 18286 39506
rect 18338 39454 18350 39506
rect 26002 39454 26014 39506
rect 26066 39454 26078 39506
rect 14926 39442 14978 39454
rect 28254 39442 28306 39454
rect 29598 39506 29650 39518
rect 29598 39442 29650 39454
rect 32286 39506 32338 39518
rect 32286 39442 32338 39454
rect 32846 39506 32898 39518
rect 32846 39442 32898 39454
rect 33070 39506 33122 39518
rect 33070 39442 33122 39454
rect 44270 39506 44322 39518
rect 44270 39442 44322 39454
rect 45838 39506 45890 39518
rect 45838 39442 45890 39454
rect 46174 39506 46226 39518
rect 46174 39442 46226 39454
rect 46846 39506 46898 39518
rect 46846 39442 46898 39454
rect 46958 39506 47010 39518
rect 46958 39442 47010 39454
rect 49086 39506 49138 39518
rect 49086 39442 49138 39454
rect 49646 39506 49698 39518
rect 51202 39454 51214 39506
rect 51266 39454 51278 39506
rect 51650 39454 51662 39506
rect 51714 39454 51726 39506
rect 49646 39442 49698 39454
rect 4062 39394 4114 39406
rect 4062 39330 4114 39342
rect 4174 39394 4226 39406
rect 4174 39330 4226 39342
rect 4286 39394 4338 39406
rect 4286 39330 4338 39342
rect 5854 39394 5906 39406
rect 5854 39330 5906 39342
rect 6078 39394 6130 39406
rect 6078 39330 6130 39342
rect 6414 39394 6466 39406
rect 15374 39394 15426 39406
rect 6738 39342 6750 39394
rect 6802 39342 6814 39394
rect 6414 39330 6466 39342
rect 15374 39330 15426 39342
rect 16046 39394 16098 39406
rect 16046 39330 16098 39342
rect 20190 39394 20242 39406
rect 20190 39330 20242 39342
rect 22542 39394 22594 39406
rect 22542 39330 22594 39342
rect 22766 39394 22818 39406
rect 22766 39330 22818 39342
rect 23102 39394 23154 39406
rect 23102 39330 23154 39342
rect 23998 39394 24050 39406
rect 23998 39330 24050 39342
rect 26686 39394 26738 39406
rect 26686 39330 26738 39342
rect 29374 39394 29426 39406
rect 29374 39330 29426 39342
rect 29710 39394 29762 39406
rect 29710 39330 29762 39342
rect 30158 39394 30210 39406
rect 30158 39330 30210 39342
rect 31950 39394 32002 39406
rect 31950 39330 32002 39342
rect 32622 39394 32674 39406
rect 32622 39330 32674 39342
rect 33294 39394 33346 39406
rect 33294 39330 33346 39342
rect 43710 39394 43762 39406
rect 43710 39330 43762 39342
rect 45278 39394 45330 39406
rect 45278 39330 45330 39342
rect 45502 39394 45554 39406
rect 45502 39330 45554 39342
rect 46062 39394 46114 39406
rect 50978 39342 50990 39394
rect 51042 39342 51054 39394
rect 46062 39330 46114 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 7646 39058 7698 39070
rect 6178 39006 6190 39058
rect 6242 39006 6254 39058
rect 7646 38994 7698 39006
rect 15150 39058 15202 39070
rect 15150 38994 15202 39006
rect 16270 39058 16322 39070
rect 16270 38994 16322 39006
rect 18846 39058 18898 39070
rect 29038 39058 29090 39070
rect 25218 39006 25230 39058
rect 25282 39006 25294 39058
rect 18846 38994 18898 39006
rect 29038 38994 29090 39006
rect 29262 39058 29314 39070
rect 29262 38994 29314 39006
rect 33742 39058 33794 39070
rect 33742 38994 33794 39006
rect 34190 39058 34242 39070
rect 34190 38994 34242 39006
rect 37662 39058 37714 39070
rect 41570 39006 41582 39058
rect 41634 39006 41646 39058
rect 46946 39006 46958 39058
rect 47010 39006 47022 39058
rect 37662 38994 37714 39006
rect 5182 38946 5234 38958
rect 2482 38894 2494 38946
rect 2546 38894 2558 38946
rect 5182 38882 5234 38894
rect 5294 38946 5346 38958
rect 13806 38946 13858 38958
rect 5842 38894 5854 38946
rect 5906 38894 5918 38946
rect 5294 38882 5346 38894
rect 13806 38882 13858 38894
rect 14478 38946 14530 38958
rect 14478 38882 14530 38894
rect 15374 38946 15426 38958
rect 15374 38882 15426 38894
rect 16158 38946 16210 38958
rect 16158 38882 16210 38894
rect 18398 38946 18450 38958
rect 18398 38882 18450 38894
rect 19742 38946 19794 38958
rect 28926 38946 28978 38958
rect 22530 38894 22542 38946
rect 22594 38894 22606 38946
rect 19742 38882 19794 38894
rect 28926 38882 28978 38894
rect 37438 38946 37490 38958
rect 37438 38882 37490 38894
rect 37998 38946 38050 38958
rect 37998 38882 38050 38894
rect 38558 38946 38610 38958
rect 45502 38946 45554 38958
rect 41906 38894 41918 38946
rect 41970 38894 41982 38946
rect 38558 38882 38610 38894
rect 45502 38882 45554 38894
rect 45950 38946 46002 38958
rect 45950 38882 46002 38894
rect 47742 38946 47794 38958
rect 47742 38882 47794 38894
rect 47854 38946 47906 38958
rect 47854 38882 47906 38894
rect 47966 38946 48018 38958
rect 47966 38882 48018 38894
rect 49758 38946 49810 38958
rect 51202 38894 51214 38946
rect 51266 38894 51278 38946
rect 49758 38882 49810 38894
rect 5406 38834 5458 38846
rect 1810 38782 1822 38834
rect 1874 38782 1886 38834
rect 5406 38770 5458 38782
rect 6526 38834 6578 38846
rect 6526 38770 6578 38782
rect 6974 38834 7026 38846
rect 6974 38770 7026 38782
rect 7422 38834 7474 38846
rect 7422 38770 7474 38782
rect 14590 38834 14642 38846
rect 15262 38834 15314 38846
rect 17726 38834 17778 38846
rect 14914 38782 14926 38834
rect 14978 38782 14990 38834
rect 15586 38782 15598 38834
rect 15650 38782 15662 38834
rect 16482 38782 16494 38834
rect 16546 38782 16558 38834
rect 14590 38770 14642 38782
rect 15262 38770 15314 38782
rect 17726 38770 17778 38782
rect 17950 38834 18002 38846
rect 20526 38834 20578 38846
rect 33966 38834 34018 38846
rect 20290 38782 20302 38834
rect 20354 38782 20366 38834
rect 21746 38782 21758 38834
rect 21810 38782 21822 38834
rect 25442 38782 25454 38834
rect 25506 38782 25518 38834
rect 31266 38782 31278 38834
rect 31330 38782 31342 38834
rect 17950 38770 18002 38782
rect 20526 38770 20578 38782
rect 33966 38770 34018 38782
rect 37326 38834 37378 38846
rect 37326 38770 37378 38782
rect 37886 38834 37938 38846
rect 37886 38770 37938 38782
rect 38222 38834 38274 38846
rect 38222 38770 38274 38782
rect 38670 38834 38722 38846
rect 43374 38834 43426 38846
rect 44606 38834 44658 38846
rect 46622 38834 46674 38846
rect 49646 38834 49698 38846
rect 41570 38782 41582 38834
rect 41634 38782 41646 38834
rect 42578 38782 42590 38834
rect 42642 38782 42654 38834
rect 43922 38782 43934 38834
rect 43986 38782 43998 38834
rect 45042 38782 45054 38834
rect 45106 38782 45118 38834
rect 49186 38782 49198 38834
rect 49250 38782 49262 38834
rect 50418 38782 50430 38834
rect 50482 38782 50494 38834
rect 38670 38770 38722 38782
rect 43374 38770 43426 38782
rect 44606 38770 44658 38782
rect 46622 38770 46674 38782
rect 49646 38770 49698 38782
rect 6750 38722 6802 38734
rect 4610 38670 4622 38722
rect 4674 38670 4686 38722
rect 6750 38658 6802 38670
rect 7534 38722 7586 38734
rect 7534 38658 7586 38670
rect 12798 38722 12850 38734
rect 12798 38658 12850 38670
rect 14254 38722 14306 38734
rect 14254 38658 14306 38670
rect 18286 38722 18338 38734
rect 26014 38722 26066 38734
rect 24658 38670 24670 38722
rect 24722 38670 24734 38722
rect 18286 38658 18338 38670
rect 26014 38658 26066 38670
rect 26462 38722 26514 38734
rect 26462 38658 26514 38670
rect 27694 38722 27746 38734
rect 27694 38658 27746 38670
rect 30830 38722 30882 38734
rect 30830 38658 30882 38670
rect 34078 38722 34130 38734
rect 34078 38658 34130 38670
rect 39230 38722 39282 38734
rect 46398 38722 46450 38734
rect 42466 38670 42478 38722
rect 42530 38670 42542 38722
rect 44146 38670 44158 38722
rect 44210 38670 44222 38722
rect 53330 38670 53342 38722
rect 53394 38670 53406 38722
rect 39230 38658 39282 38670
rect 46398 38658 46450 38670
rect 38558 38610 38610 38622
rect 17378 38558 17390 38610
rect 17442 38558 17454 38610
rect 47282 38558 47294 38610
rect 47346 38558 47358 38610
rect 38558 38546 38610 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 27022 38274 27074 38286
rect 27022 38210 27074 38222
rect 45838 38274 45890 38286
rect 45838 38210 45890 38222
rect 19966 38162 20018 38174
rect 4610 38110 4622 38162
rect 4674 38110 4686 38162
rect 8754 38110 8766 38162
rect 8818 38110 8830 38162
rect 9650 38110 9662 38162
rect 9714 38110 9726 38162
rect 17602 38110 17614 38162
rect 17666 38110 17678 38162
rect 19966 38098 20018 38110
rect 21758 38162 21810 38174
rect 21758 38098 21810 38110
rect 22990 38162 23042 38174
rect 27918 38162 27970 38174
rect 27346 38110 27358 38162
rect 27410 38110 27422 38162
rect 32498 38110 32510 38162
rect 32562 38110 32574 38162
rect 34626 38110 34638 38162
rect 34690 38110 34702 38162
rect 55010 38110 55022 38162
rect 55074 38110 55086 38162
rect 22990 38098 23042 38110
rect 27918 38098 27970 38110
rect 14702 38050 14754 38062
rect 1810 37998 1822 38050
rect 1874 37998 1886 38050
rect 5954 37998 5966 38050
rect 6018 37998 6030 38050
rect 12562 37998 12574 38050
rect 12626 37998 12638 38050
rect 14702 37986 14754 37998
rect 15038 38050 15090 38062
rect 25230 38050 25282 38062
rect 15810 37998 15822 38050
rect 15874 37998 15886 38050
rect 18162 37998 18174 38050
rect 18226 37998 18238 38050
rect 24770 37998 24782 38050
rect 24834 37998 24846 38050
rect 15038 37986 15090 37998
rect 25230 37986 25282 37998
rect 28590 38050 28642 38062
rect 28590 37986 28642 37998
rect 29486 38050 29538 38062
rect 29486 37986 29538 37998
rect 30270 38050 30322 38062
rect 37214 38050 37266 38062
rect 31714 37998 31726 38050
rect 31778 37998 31790 38050
rect 30270 37986 30322 37998
rect 37214 37986 37266 37998
rect 37998 38050 38050 38062
rect 37998 37986 38050 37998
rect 38110 38050 38162 38062
rect 38110 37986 38162 37998
rect 38222 38050 38274 38062
rect 38222 37986 38274 37998
rect 38446 38050 38498 38062
rect 43710 38050 43762 38062
rect 39666 37998 39678 38050
rect 39730 37998 39742 38050
rect 38446 37986 38498 37998
rect 43710 37986 43762 37998
rect 44718 38050 44770 38062
rect 44718 37986 44770 37998
rect 45726 38050 45778 38062
rect 48974 38050 49026 38062
rect 51326 38050 51378 38062
rect 54574 38050 54626 38062
rect 47058 37998 47070 38050
rect 47122 37998 47134 38050
rect 48290 37998 48302 38050
rect 48354 37998 48366 38050
rect 49634 37998 49646 38050
rect 49698 37998 49710 38050
rect 51762 37998 51774 38050
rect 51826 37998 51838 38050
rect 52882 37998 52894 38050
rect 52946 37998 52958 38050
rect 45726 37986 45778 37998
rect 48974 37986 49026 37998
rect 51326 37986 51378 37998
rect 54574 37986 54626 37998
rect 14366 37938 14418 37950
rect 2482 37886 2494 37938
rect 2546 37886 2558 37938
rect 6626 37886 6638 37938
rect 6690 37886 6702 37938
rect 11778 37886 11790 37938
rect 11842 37886 11854 37938
rect 14366 37874 14418 37886
rect 14814 37938 14866 37950
rect 14814 37874 14866 37886
rect 18734 37938 18786 37950
rect 18734 37874 18786 37886
rect 21422 37938 21474 37950
rect 21422 37874 21474 37886
rect 23998 37938 24050 37950
rect 23998 37874 24050 37886
rect 24334 37938 24386 37950
rect 29822 37938 29874 37950
rect 26562 37886 26574 37938
rect 26626 37886 26638 37938
rect 24334 37874 24386 37886
rect 29822 37874 29874 37886
rect 30718 37938 30770 37950
rect 30718 37874 30770 37886
rect 31054 37938 31106 37950
rect 31054 37874 31106 37886
rect 37326 37938 37378 37950
rect 37326 37874 37378 37886
rect 38782 37938 38834 37950
rect 38782 37874 38834 37886
rect 39342 37938 39394 37950
rect 39342 37874 39394 37886
rect 42478 37938 42530 37950
rect 42478 37874 42530 37886
rect 42814 37938 42866 37950
rect 42814 37874 42866 37886
rect 44942 37938 44994 37950
rect 44942 37874 44994 37886
rect 45166 37938 45218 37950
rect 45166 37874 45218 37886
rect 45390 37938 45442 37950
rect 45390 37874 45442 37886
rect 45838 37938 45890 37950
rect 45838 37874 45890 37886
rect 46398 37938 46450 37950
rect 46398 37874 46450 37886
rect 48862 37938 48914 37950
rect 52770 37886 52782 37938
rect 52834 37886 52846 37938
rect 53330 37886 53342 37938
rect 53394 37886 53406 37938
rect 48862 37874 48914 37886
rect 5070 37826 5122 37838
rect 5070 37762 5122 37774
rect 9214 37826 9266 37838
rect 9214 37762 9266 37774
rect 13694 37826 13746 37838
rect 19630 37826 19682 37838
rect 14018 37774 14030 37826
rect 14082 37774 14094 37826
rect 13694 37762 13746 37774
rect 19630 37762 19682 37774
rect 21310 37826 21362 37838
rect 21310 37762 21362 37774
rect 21870 37826 21922 37838
rect 21870 37762 21922 37774
rect 22542 37826 22594 37838
rect 22542 37762 22594 37774
rect 26014 37826 26066 37838
rect 26014 37762 26066 37774
rect 26238 37826 26290 37838
rect 26238 37762 26290 37774
rect 27246 37826 27298 37838
rect 35086 37826 35138 37838
rect 28242 37774 28254 37826
rect 28306 37774 28318 37826
rect 27246 37762 27298 37774
rect 35086 37762 35138 37774
rect 36206 37826 36258 37838
rect 36206 37762 36258 37774
rect 37102 37826 37154 37838
rect 37102 37762 37154 37774
rect 37774 37826 37826 37838
rect 37774 37762 37826 37774
rect 38670 37826 38722 37838
rect 38670 37762 38722 37774
rect 39454 37826 39506 37838
rect 39454 37762 39506 37774
rect 43486 37826 43538 37838
rect 43486 37762 43538 37774
rect 43822 37826 43874 37838
rect 43822 37762 43874 37774
rect 44382 37826 44434 37838
rect 44382 37762 44434 37774
rect 51102 37826 51154 37838
rect 51102 37762 51154 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 3502 37490 3554 37502
rect 3502 37426 3554 37438
rect 4398 37490 4450 37502
rect 4398 37426 4450 37438
rect 5182 37490 5234 37502
rect 5182 37426 5234 37438
rect 6526 37490 6578 37502
rect 6526 37426 6578 37438
rect 6638 37490 6690 37502
rect 6638 37426 6690 37438
rect 14142 37490 14194 37502
rect 14142 37426 14194 37438
rect 17502 37490 17554 37502
rect 17502 37426 17554 37438
rect 18174 37490 18226 37502
rect 18174 37426 18226 37438
rect 22990 37490 23042 37502
rect 36430 37490 36482 37502
rect 31490 37438 31502 37490
rect 31554 37438 31566 37490
rect 22990 37426 23042 37438
rect 36430 37426 36482 37438
rect 40238 37490 40290 37502
rect 40238 37426 40290 37438
rect 50206 37490 50258 37502
rect 50206 37426 50258 37438
rect 50990 37490 51042 37502
rect 50990 37426 51042 37438
rect 3726 37378 3778 37390
rect 3726 37314 3778 37326
rect 3950 37378 4002 37390
rect 3950 37314 4002 37326
rect 4622 37378 4674 37390
rect 4622 37314 4674 37326
rect 4846 37378 4898 37390
rect 4846 37314 4898 37326
rect 5518 37378 5570 37390
rect 5518 37314 5570 37326
rect 6750 37378 6802 37390
rect 17390 37378 17442 37390
rect 24334 37378 24386 37390
rect 36206 37378 36258 37390
rect 11778 37326 11790 37378
rect 11842 37326 11854 37378
rect 15362 37326 15374 37378
rect 15426 37326 15438 37378
rect 16370 37326 16382 37378
rect 16434 37326 16446 37378
rect 17826 37326 17838 37378
rect 17890 37326 17902 37378
rect 20850 37326 20862 37378
rect 20914 37326 20926 37378
rect 22082 37326 22094 37378
rect 22146 37326 22158 37378
rect 27906 37326 27918 37378
rect 27970 37326 27982 37378
rect 6750 37314 6802 37326
rect 17390 37314 17442 37326
rect 24334 37314 24386 37326
rect 36206 37314 36258 37326
rect 37102 37378 37154 37390
rect 37102 37314 37154 37326
rect 37214 37378 37266 37390
rect 56142 37378 56194 37390
rect 37650 37326 37662 37378
rect 37714 37326 37726 37378
rect 37986 37326 37998 37378
rect 38050 37326 38062 37378
rect 44146 37326 44158 37378
rect 44210 37326 44222 37378
rect 45714 37326 45726 37378
rect 45778 37326 45790 37378
rect 37214 37314 37266 37326
rect 56142 37314 56194 37326
rect 3390 37266 3442 37278
rect 3390 37202 3442 37214
rect 4286 37266 4338 37278
rect 19630 37266 19682 37278
rect 11106 37214 11118 37266
rect 11170 37214 11182 37266
rect 14354 37214 14366 37266
rect 14418 37214 14430 37266
rect 15586 37214 15598 37266
rect 15650 37214 15662 37266
rect 16034 37214 16046 37266
rect 16098 37214 16110 37266
rect 18610 37214 18622 37266
rect 18674 37214 18686 37266
rect 19058 37214 19070 37266
rect 19122 37214 19134 37266
rect 4286 37202 4338 37214
rect 19630 37202 19682 37214
rect 20078 37266 20130 37278
rect 20078 37202 20130 37214
rect 20302 37266 20354 37278
rect 20302 37202 20354 37214
rect 21198 37266 21250 37278
rect 22430 37266 22482 37278
rect 21634 37214 21646 37266
rect 21698 37214 21710 37266
rect 21198 37202 21250 37214
rect 22430 37202 22482 37214
rect 23326 37266 23378 37278
rect 23326 37202 23378 37214
rect 23886 37266 23938 37278
rect 25230 37266 25282 37278
rect 30494 37266 30546 37278
rect 24658 37214 24670 37266
rect 24722 37214 24734 37266
rect 25890 37214 25902 37266
rect 25954 37214 25966 37266
rect 27234 37214 27246 37266
rect 27298 37214 27310 37266
rect 23886 37202 23938 37214
rect 25230 37202 25282 37214
rect 30494 37202 30546 37214
rect 31166 37266 31218 37278
rect 36542 37266 36594 37278
rect 32386 37214 32398 37266
rect 32450 37214 32462 37266
rect 33058 37214 33070 37266
rect 33122 37214 33134 37266
rect 31166 37202 31218 37214
rect 36542 37202 36594 37214
rect 36990 37266 37042 37278
rect 48750 37266 48802 37278
rect 38210 37214 38222 37266
rect 38274 37214 38286 37266
rect 39778 37214 39790 37266
rect 39842 37214 39854 37266
rect 43810 37214 43822 37266
rect 43874 37214 43886 37266
rect 44818 37214 44830 37266
rect 44882 37214 44894 37266
rect 45826 37214 45838 37266
rect 45890 37214 45902 37266
rect 36990 37202 37042 37214
rect 48750 37202 48802 37214
rect 48974 37266 49026 37278
rect 48974 37202 49026 37214
rect 49422 37266 49474 37278
rect 55022 37266 55074 37278
rect 54114 37214 54126 37266
rect 54178 37214 54190 37266
rect 49422 37202 49474 37214
rect 55022 37202 55074 37214
rect 19854 37154 19906 37166
rect 13906 37102 13918 37154
rect 13970 37102 13982 37154
rect 19854 37090 19906 37102
rect 24446 37154 24498 37166
rect 26686 37154 26738 37166
rect 30942 37154 30994 37166
rect 48190 37154 48242 37166
rect 26114 37102 26126 37154
rect 26178 37102 26190 37154
rect 30034 37102 30046 37154
rect 30098 37102 30110 37154
rect 32050 37102 32062 37154
rect 32114 37102 32126 37154
rect 33842 37102 33854 37154
rect 33906 37102 33918 37154
rect 35970 37102 35982 37154
rect 36034 37102 36046 37154
rect 40898 37102 40910 37154
rect 40962 37102 40974 37154
rect 43026 37102 43038 37154
rect 43090 37102 43102 37154
rect 45266 37102 45278 37154
rect 45330 37102 45342 37154
rect 24446 37090 24498 37102
rect 26686 37090 26738 37102
rect 30942 37090 30994 37102
rect 48190 37090 48242 37102
rect 49198 37154 49250 37166
rect 49198 37090 49250 37102
rect 50430 37154 50482 37166
rect 54574 37154 54626 37166
rect 51314 37102 51326 37154
rect 51378 37102 51390 37154
rect 53442 37102 53454 37154
rect 53506 37102 53518 37154
rect 50430 37090 50482 37102
rect 54574 37090 54626 37102
rect 56702 37154 56754 37166
rect 56702 37090 56754 37102
rect 57262 37154 57314 37166
rect 57262 37090 57314 37102
rect 54798 37042 54850 37054
rect 18610 36990 18622 37042
rect 18674 36990 18686 37042
rect 22642 36990 22654 37042
rect 22706 37039 22718 37042
rect 22978 37039 22990 37042
rect 22706 36993 22990 37039
rect 22706 36990 22718 36993
rect 22978 36990 22990 36993
rect 23042 36990 23054 37042
rect 54798 36978 54850 36990
rect 55470 37042 55522 37054
rect 55470 36978 55522 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 14590 36706 14642 36718
rect 33742 36706 33794 36718
rect 15586 36654 15598 36706
rect 15650 36654 15662 36706
rect 14590 36642 14642 36654
rect 33742 36642 33794 36654
rect 37214 36706 37266 36718
rect 37214 36642 37266 36654
rect 37550 36706 37602 36718
rect 37550 36642 37602 36654
rect 48862 36706 48914 36718
rect 48862 36642 48914 36654
rect 16158 36594 16210 36606
rect 28142 36594 28194 36606
rect 22082 36542 22094 36594
rect 22146 36542 22158 36594
rect 22530 36542 22542 36594
rect 22594 36542 22606 36594
rect 16158 36530 16210 36542
rect 28142 36530 28194 36542
rect 28590 36594 28642 36606
rect 28590 36530 28642 36542
rect 30046 36594 30098 36606
rect 30046 36530 30098 36542
rect 33854 36594 33906 36606
rect 39006 36594 39058 36606
rect 46846 36594 46898 36606
rect 38546 36542 38558 36594
rect 38610 36542 38622 36594
rect 40338 36542 40350 36594
rect 40402 36542 40414 36594
rect 42466 36542 42478 36594
rect 42530 36542 42542 36594
rect 33854 36530 33906 36542
rect 39006 36530 39058 36542
rect 46846 36530 46898 36542
rect 47630 36594 47682 36606
rect 47630 36530 47682 36542
rect 51662 36594 51714 36606
rect 51662 36530 51714 36542
rect 54686 36594 54738 36606
rect 55570 36542 55582 36594
rect 55634 36542 55646 36594
rect 54686 36530 54738 36542
rect 13694 36482 13746 36494
rect 13694 36418 13746 36430
rect 14030 36482 14082 36494
rect 14478 36482 14530 36494
rect 14242 36430 14254 36482
rect 14306 36430 14318 36482
rect 14030 36418 14082 36430
rect 14478 36418 14530 36430
rect 15262 36482 15314 36494
rect 15262 36418 15314 36430
rect 15934 36482 15986 36494
rect 15934 36418 15986 36430
rect 17278 36482 17330 36494
rect 17278 36418 17330 36430
rect 18958 36482 19010 36494
rect 18958 36418 19010 36430
rect 19406 36482 19458 36494
rect 19406 36418 19458 36430
rect 19742 36482 19794 36494
rect 19742 36418 19794 36430
rect 20078 36482 20130 36494
rect 20078 36418 20130 36430
rect 20526 36482 20578 36494
rect 23326 36482 23378 36494
rect 21970 36430 21982 36482
rect 22034 36430 22046 36482
rect 22418 36430 22430 36482
rect 22482 36430 22494 36482
rect 20526 36418 20578 36430
rect 23326 36418 23378 36430
rect 23998 36482 24050 36494
rect 23998 36418 24050 36430
rect 27358 36482 27410 36494
rect 27358 36418 27410 36430
rect 29486 36482 29538 36494
rect 29486 36418 29538 36430
rect 31166 36482 31218 36494
rect 31166 36418 31218 36430
rect 31502 36482 31554 36494
rect 36990 36482 37042 36494
rect 43934 36482 43986 36494
rect 45166 36482 45218 36494
rect 36082 36430 36094 36482
rect 36146 36430 36158 36482
rect 38322 36430 38334 36482
rect 38386 36430 38398 36482
rect 39554 36430 39566 36482
rect 39618 36430 39630 36482
rect 44818 36430 44830 36482
rect 44882 36430 44894 36482
rect 31502 36418 31554 36430
rect 36990 36418 37042 36430
rect 43934 36418 43986 36430
rect 45166 36418 45218 36430
rect 45278 36482 45330 36494
rect 45278 36418 45330 36430
rect 45502 36482 45554 36494
rect 45502 36418 45554 36430
rect 45726 36482 45778 36494
rect 45726 36418 45778 36430
rect 46062 36482 46114 36494
rect 46062 36418 46114 36430
rect 47742 36482 47794 36494
rect 47742 36418 47794 36430
rect 48190 36482 48242 36494
rect 56030 36482 56082 36494
rect 49858 36430 49870 36482
rect 49922 36430 49934 36482
rect 50194 36430 50206 36482
rect 50258 36430 50270 36482
rect 52658 36430 52670 36482
rect 52722 36430 52734 36482
rect 54114 36430 54126 36482
rect 54178 36430 54190 36482
rect 54786 36430 54798 36482
rect 54850 36430 54862 36482
rect 55458 36430 55470 36482
rect 55522 36430 55534 36482
rect 48190 36418 48242 36430
rect 56030 36418 56082 36430
rect 56366 36482 56418 36494
rect 56366 36418 56418 36430
rect 13806 36370 13858 36382
rect 13806 36306 13858 36318
rect 18062 36370 18114 36382
rect 18062 36306 18114 36318
rect 20750 36370 20802 36382
rect 33966 36370 34018 36382
rect 47518 36370 47570 36382
rect 56702 36370 56754 36382
rect 25218 36318 25230 36370
rect 25282 36318 25294 36370
rect 27682 36318 27694 36370
rect 27746 36318 27758 36370
rect 32498 36318 32510 36370
rect 32562 36318 32574 36370
rect 35858 36318 35870 36370
rect 35922 36318 35934 36370
rect 46386 36318 46398 36370
rect 46450 36318 46462 36370
rect 50866 36318 50878 36370
rect 50930 36318 50942 36370
rect 52882 36318 52894 36370
rect 52946 36318 52958 36370
rect 20750 36306 20802 36318
rect 33966 36306 34018 36318
rect 47518 36306 47570 36318
rect 56702 36306 56754 36318
rect 57038 36370 57090 36382
rect 57038 36306 57090 36318
rect 12910 36258 12962 36270
rect 19518 36258 19570 36270
rect 14914 36206 14926 36258
rect 14978 36206 14990 36258
rect 17154 36206 17166 36258
rect 17218 36206 17230 36258
rect 12910 36194 12962 36206
rect 19518 36194 19570 36206
rect 20302 36258 20354 36270
rect 20302 36194 20354 36206
rect 23102 36258 23154 36270
rect 23102 36194 23154 36206
rect 23774 36258 23826 36270
rect 23774 36194 23826 36206
rect 23886 36258 23938 36270
rect 24894 36258 24946 36270
rect 24546 36206 24558 36258
rect 24610 36206 24622 36258
rect 23886 36194 23938 36206
rect 24894 36194 24946 36206
rect 25566 36258 25618 36270
rect 25566 36194 25618 36206
rect 30830 36258 30882 36270
rect 30830 36194 30882 36206
rect 31838 36258 31890 36270
rect 31838 36194 31890 36206
rect 32174 36258 32226 36270
rect 32174 36194 32226 36206
rect 42926 36258 42978 36270
rect 42926 36194 42978 36206
rect 43598 36258 43650 36270
rect 48638 36258 48690 36270
rect 44258 36206 44270 36258
rect 44322 36206 44334 36258
rect 45154 36206 45166 36258
rect 45218 36206 45230 36258
rect 43598 36194 43650 36206
rect 48638 36194 48690 36206
rect 48750 36258 48802 36270
rect 48750 36194 48802 36206
rect 52110 36258 52162 36270
rect 56254 36258 56306 36270
rect 53106 36206 53118 36258
rect 53170 36206 53182 36258
rect 54002 36206 54014 36258
rect 54066 36206 54078 36258
rect 52110 36194 52162 36206
rect 56254 36194 56306 36206
rect 57150 36258 57202 36270
rect 57150 36194 57202 36206
rect 57262 36258 57314 36270
rect 57262 36194 57314 36206
rect 57822 36258 57874 36270
rect 57822 36194 57874 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 17390 35922 17442 35934
rect 14914 35870 14926 35922
rect 14978 35870 14990 35922
rect 17390 35858 17442 35870
rect 18398 35922 18450 35934
rect 18398 35858 18450 35870
rect 18622 35922 18674 35934
rect 18622 35858 18674 35870
rect 18958 35922 19010 35934
rect 25566 35922 25618 35934
rect 25218 35870 25230 35922
rect 25282 35870 25294 35922
rect 18958 35858 19010 35870
rect 25566 35858 25618 35870
rect 28030 35922 28082 35934
rect 28030 35858 28082 35870
rect 29262 35922 29314 35934
rect 29262 35858 29314 35870
rect 29374 35922 29426 35934
rect 29374 35858 29426 35870
rect 29710 35922 29762 35934
rect 29710 35858 29762 35870
rect 30270 35922 30322 35934
rect 30270 35858 30322 35870
rect 30718 35922 30770 35934
rect 30718 35858 30770 35870
rect 43486 35922 43538 35934
rect 43486 35858 43538 35870
rect 43822 35922 43874 35934
rect 43822 35858 43874 35870
rect 45502 35922 45554 35934
rect 45502 35858 45554 35870
rect 45950 35922 46002 35934
rect 45950 35858 46002 35870
rect 54574 35922 54626 35934
rect 54574 35858 54626 35870
rect 57934 35922 57986 35934
rect 57934 35858 57986 35870
rect 15822 35810 15874 35822
rect 15822 35746 15874 35758
rect 16830 35810 16882 35822
rect 16830 35746 16882 35758
rect 19070 35810 19122 35822
rect 30494 35810 30546 35822
rect 36654 35810 36706 35822
rect 21522 35758 21534 35810
rect 21586 35758 21598 35810
rect 28578 35758 28590 35810
rect 28642 35758 28654 35810
rect 33730 35758 33742 35810
rect 33794 35758 33806 35810
rect 19070 35746 19122 35758
rect 30494 35746 30546 35758
rect 36654 35746 36706 35758
rect 47070 35810 47122 35822
rect 47070 35746 47122 35758
rect 54462 35810 54514 35822
rect 54462 35746 54514 35758
rect 56030 35810 56082 35822
rect 56030 35746 56082 35758
rect 16046 35698 16098 35710
rect 12002 35646 12014 35698
rect 12066 35646 12078 35698
rect 16046 35634 16098 35646
rect 17726 35698 17778 35710
rect 17726 35634 17778 35646
rect 17950 35698 18002 35710
rect 26126 35698 26178 35710
rect 29486 35698 29538 35710
rect 22306 35646 22318 35698
rect 22370 35646 22382 35698
rect 23202 35646 23214 35698
rect 23266 35646 23278 35698
rect 23874 35646 23886 35698
rect 23938 35646 23950 35698
rect 28242 35646 28254 35698
rect 28306 35646 28318 35698
rect 28802 35646 28814 35698
rect 28866 35646 28878 35698
rect 17950 35634 18002 35646
rect 26126 35634 26178 35646
rect 29486 35634 29538 35646
rect 34078 35698 34130 35710
rect 37550 35698 37602 35710
rect 39118 35698 39170 35710
rect 37314 35646 37326 35698
rect 37378 35646 37390 35698
rect 38210 35646 38222 35698
rect 38274 35646 38286 35698
rect 34078 35634 34130 35646
rect 37550 35634 37602 35646
rect 39118 35634 39170 35646
rect 39454 35698 39506 35710
rect 40238 35698 40290 35710
rect 39778 35646 39790 35698
rect 39842 35646 39854 35698
rect 39454 35634 39506 35646
rect 40238 35634 40290 35646
rect 44718 35698 44770 35710
rect 44718 35634 44770 35646
rect 44942 35698 44994 35710
rect 45726 35698 45778 35710
rect 47966 35698 48018 35710
rect 54798 35698 54850 35710
rect 56590 35698 56642 35710
rect 45154 35646 45166 35698
rect 45218 35646 45230 35698
rect 47618 35646 47630 35698
rect 47682 35646 47694 35698
rect 48738 35646 48750 35698
rect 48802 35646 48814 35698
rect 49634 35646 49646 35698
rect 49698 35646 49710 35698
rect 50754 35646 50766 35698
rect 50818 35646 50830 35698
rect 51426 35646 51438 35698
rect 51490 35646 51502 35698
rect 52546 35646 52558 35698
rect 52610 35646 52622 35698
rect 55346 35646 55358 35698
rect 55410 35646 55422 35698
rect 44942 35634 44994 35646
rect 45726 35634 45778 35646
rect 47966 35634 48018 35646
rect 54798 35634 54850 35646
rect 56590 35634 56642 35646
rect 56926 35698 56978 35710
rect 57138 35646 57150 35698
rect 57202 35646 57214 35698
rect 56926 35634 56978 35646
rect 15598 35586 15650 35598
rect 12674 35534 12686 35586
rect 12738 35534 12750 35586
rect 15598 35522 15650 35534
rect 18510 35586 18562 35598
rect 27918 35586 27970 35598
rect 19394 35534 19406 35586
rect 19458 35534 19470 35586
rect 23426 35534 23438 35586
rect 23490 35534 23502 35586
rect 18510 35522 18562 35534
rect 27918 35522 27970 35534
rect 30382 35586 30434 35598
rect 44382 35586 44434 35598
rect 38322 35534 38334 35586
rect 38386 35534 38398 35586
rect 30382 35522 30434 35534
rect 44382 35522 44434 35534
rect 45614 35586 45666 35598
rect 45614 35522 45666 35534
rect 46622 35586 46674 35598
rect 56702 35586 56754 35598
rect 50418 35534 50430 35586
rect 50482 35534 50494 35586
rect 53330 35534 53342 35586
rect 53394 35534 53406 35586
rect 55122 35534 55134 35586
rect 55186 35534 55198 35586
rect 46622 35522 46674 35534
rect 56702 35522 56754 35534
rect 57822 35586 57874 35598
rect 57822 35522 57874 35534
rect 16382 35474 16434 35486
rect 16382 35410 16434 35422
rect 16718 35474 16770 35486
rect 39790 35474 39842 35486
rect 23314 35422 23326 35474
rect 23378 35422 23390 35474
rect 16718 35410 16770 35422
rect 39790 35410 39842 35422
rect 44606 35474 44658 35486
rect 44606 35410 44658 35422
rect 48750 35474 48802 35486
rect 48750 35410 48802 35422
rect 49086 35474 49138 35486
rect 57710 35474 57762 35486
rect 57138 35422 57150 35474
rect 57202 35422 57214 35474
rect 49086 35410 49138 35422
rect 57710 35410 57762 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 13806 35138 13858 35150
rect 13806 35074 13858 35086
rect 18958 35138 19010 35150
rect 18958 35074 19010 35086
rect 29486 35138 29538 35150
rect 29486 35074 29538 35086
rect 30606 35138 30658 35150
rect 30606 35074 30658 35086
rect 34638 35138 34690 35150
rect 34638 35074 34690 35086
rect 35086 35138 35138 35150
rect 35086 35074 35138 35086
rect 43822 35138 43874 35150
rect 43822 35074 43874 35086
rect 45278 35138 45330 35150
rect 51538 35086 51550 35138
rect 51602 35086 51614 35138
rect 52882 35086 52894 35138
rect 52946 35086 52958 35138
rect 57138 35086 57150 35138
rect 57202 35086 57214 35138
rect 45278 35074 45330 35086
rect 15038 35026 15090 35038
rect 18734 35026 18786 35038
rect 34414 35026 34466 35038
rect 13570 34974 13582 35026
rect 13634 34974 13646 35026
rect 18162 34974 18174 35026
rect 18226 34974 18238 35026
rect 20514 34974 20526 35026
rect 20578 34974 20590 35026
rect 22418 34974 22430 35026
rect 22482 34974 22494 35026
rect 23874 34974 23886 35026
rect 23938 34974 23950 35026
rect 26002 34974 26014 35026
rect 26066 34974 26078 35026
rect 15038 34962 15090 34974
rect 18734 34962 18786 34974
rect 34414 34962 34466 34974
rect 34862 35026 34914 35038
rect 47182 35026 47234 35038
rect 53342 35026 53394 35038
rect 38098 34974 38110 35026
rect 38162 34974 38174 35026
rect 40002 34974 40014 35026
rect 40066 34974 40078 35026
rect 42130 34974 42142 35026
rect 42194 34974 42206 35026
rect 51090 34974 51102 35026
rect 51154 34974 51166 35026
rect 54114 34974 54126 35026
rect 54178 34974 54190 35026
rect 34862 34962 34914 34974
rect 47182 34962 47234 34974
rect 53342 34962 53394 34974
rect 21310 34914 21362 34926
rect 15362 34862 15374 34914
rect 15426 34862 15438 34914
rect 19282 34862 19294 34914
rect 19346 34862 19358 34914
rect 19618 34862 19630 34914
rect 19682 34862 19694 34914
rect 20626 34862 20638 34914
rect 20690 34862 20702 34914
rect 21310 34850 21362 34862
rect 21422 34914 21474 34926
rect 26462 34914 26514 34926
rect 23202 34862 23214 34914
rect 23266 34862 23278 34914
rect 21422 34850 21474 34862
rect 26462 34850 26514 34862
rect 27022 34914 27074 34926
rect 33406 34914 33458 34926
rect 44718 34914 44770 34926
rect 29138 34862 29150 34914
rect 29202 34862 29214 34914
rect 30258 34862 30270 34914
rect 30322 34862 30334 34914
rect 39330 34862 39342 34914
rect 39394 34862 39406 34914
rect 44146 34862 44158 34914
rect 44210 34862 44222 34914
rect 27022 34850 27074 34862
rect 33406 34850 33458 34862
rect 44718 34850 44770 34862
rect 45166 34914 45218 34926
rect 45166 34850 45218 34862
rect 45502 34914 45554 34926
rect 45502 34850 45554 34862
rect 46286 34914 46338 34926
rect 46286 34850 46338 34862
rect 47070 34914 47122 34926
rect 47070 34850 47122 34862
rect 47294 34914 47346 34926
rect 48514 34862 48526 34914
rect 48578 34862 48590 34914
rect 49298 34862 49310 34914
rect 49362 34862 49374 34914
rect 49522 34862 49534 34914
rect 49586 34862 49598 34914
rect 50978 34862 50990 34914
rect 51042 34862 51054 34914
rect 52658 34862 52670 34914
rect 52722 34862 52734 34914
rect 56802 34862 56814 34914
rect 56866 34862 56878 34914
rect 57138 34862 57150 34914
rect 57202 34862 57214 34914
rect 47294 34850 47346 34862
rect 13582 34802 13634 34814
rect 21982 34802 22034 34814
rect 16034 34750 16046 34802
rect 16098 34750 16110 34802
rect 20738 34750 20750 34802
rect 20802 34750 20814 34802
rect 13582 34738 13634 34750
rect 21982 34738 22034 34750
rect 33182 34802 33234 34814
rect 45726 34802 45778 34814
rect 37874 34750 37886 34802
rect 37938 34750 37950 34802
rect 33182 34738 33234 34750
rect 45726 34738 45778 34750
rect 46398 34802 46450 34814
rect 53454 34802 53506 34814
rect 56590 34802 56642 34814
rect 53218 34750 53230 34802
rect 53282 34750 53294 34802
rect 54338 34750 54350 34802
rect 54402 34750 54414 34802
rect 56018 34750 56030 34802
rect 56082 34750 56094 34802
rect 46398 34738 46450 34750
rect 53454 34738 53506 34750
rect 56590 34738 56642 34750
rect 57822 34802 57874 34814
rect 57822 34738 57874 34750
rect 19070 34690 19122 34702
rect 19070 34626 19122 34638
rect 29374 34690 29426 34702
rect 29374 34626 29426 34638
rect 30494 34690 30546 34702
rect 30494 34626 30546 34638
rect 33854 34690 33906 34702
rect 33854 34626 33906 34638
rect 33966 34690 34018 34702
rect 33966 34626 34018 34638
rect 34078 34690 34130 34702
rect 34078 34626 34130 34638
rect 35534 34690 35586 34702
rect 35534 34626 35586 34638
rect 36318 34690 36370 34702
rect 36318 34626 36370 34638
rect 37102 34690 37154 34702
rect 37102 34626 37154 34638
rect 42590 34690 42642 34702
rect 42590 34626 42642 34638
rect 43486 34690 43538 34702
rect 43486 34626 43538 34638
rect 43934 34690 43986 34702
rect 46846 34690 46898 34702
rect 57710 34690 57762 34702
rect 45154 34638 45166 34690
rect 45218 34638 45230 34690
rect 55906 34638 55918 34690
rect 55970 34638 55982 34690
rect 57026 34638 57038 34690
rect 57090 34638 57102 34690
rect 43934 34626 43986 34638
rect 46846 34626 46898 34638
rect 57710 34626 57762 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 15598 34354 15650 34366
rect 15598 34290 15650 34302
rect 16382 34354 16434 34366
rect 16382 34290 16434 34302
rect 21870 34354 21922 34366
rect 21870 34290 21922 34302
rect 22766 34354 22818 34366
rect 22766 34290 22818 34302
rect 25454 34354 25506 34366
rect 25454 34290 25506 34302
rect 36430 34354 36482 34366
rect 36430 34290 36482 34302
rect 46398 34354 46450 34366
rect 46398 34290 46450 34302
rect 48974 34354 49026 34366
rect 48974 34290 49026 34302
rect 49982 34354 50034 34366
rect 49982 34290 50034 34302
rect 16606 34242 16658 34254
rect 16606 34178 16658 34190
rect 16830 34242 16882 34254
rect 16830 34178 16882 34190
rect 25902 34242 25954 34254
rect 36542 34242 36594 34254
rect 48190 34242 48242 34254
rect 27122 34190 27134 34242
rect 27186 34190 27198 34242
rect 30370 34190 30382 34242
rect 30434 34190 30446 34242
rect 41010 34190 41022 34242
rect 41074 34190 41086 34242
rect 42578 34190 42590 34242
rect 42642 34190 42654 34242
rect 43810 34190 43822 34242
rect 43874 34190 43886 34242
rect 25902 34178 25954 34190
rect 36542 34178 36594 34190
rect 48190 34178 48242 34190
rect 50206 34242 50258 34254
rect 50206 34178 50258 34190
rect 50654 34242 50706 34254
rect 50654 34178 50706 34190
rect 56030 34242 56082 34254
rect 56030 34178 56082 34190
rect 16270 34130 16322 34142
rect 20862 34130 20914 34142
rect 48750 34130 48802 34142
rect 56478 34130 56530 34142
rect 14466 34078 14478 34130
rect 14530 34078 14542 34130
rect 17938 34078 17950 34130
rect 18002 34078 18014 34130
rect 24658 34078 24670 34130
rect 24722 34078 24734 34130
rect 26450 34078 26462 34130
rect 26514 34078 26526 34130
rect 29586 34078 29598 34130
rect 29650 34078 29662 34130
rect 33170 34078 33182 34130
rect 33234 34078 33246 34130
rect 37090 34078 37102 34130
rect 37154 34078 37166 34130
rect 38770 34078 38782 34130
rect 38834 34078 38846 34130
rect 40898 34078 40910 34130
rect 40962 34078 40974 34130
rect 42018 34078 42030 34130
rect 42082 34078 42094 34130
rect 43138 34078 43150 34130
rect 43202 34078 43214 34130
rect 47618 34078 47630 34130
rect 47682 34078 47694 34130
rect 48066 34078 48078 34130
rect 48130 34078 48142 34130
rect 49186 34078 49198 34130
rect 49250 34078 49262 34130
rect 49410 34078 49422 34130
rect 49474 34078 49486 34130
rect 51762 34078 51774 34130
rect 51826 34078 51838 34130
rect 53106 34078 53118 34130
rect 53170 34078 53182 34130
rect 53554 34078 53566 34130
rect 53618 34078 53630 34130
rect 53890 34078 53902 34130
rect 53954 34078 53966 34130
rect 16270 34066 16322 34078
rect 20862 34066 20914 34078
rect 48750 34066 48802 34078
rect 56478 34066 56530 34078
rect 56814 34130 56866 34142
rect 57250 34078 57262 34130
rect 57314 34078 57326 34130
rect 56814 34066 56866 34078
rect 20302 34018 20354 34030
rect 19730 33966 19742 34018
rect 19794 33966 19806 34018
rect 20302 33954 20354 33966
rect 21310 34018 21362 34030
rect 21310 33954 21362 33966
rect 23214 34018 23266 34030
rect 23214 33954 23266 33966
rect 24446 34018 24498 34030
rect 55582 34018 55634 34030
rect 29250 33966 29262 34018
rect 29314 33966 29326 34018
rect 32498 33966 32510 34018
rect 32562 33966 32574 34018
rect 33842 33966 33854 34018
rect 33906 33966 33918 34018
rect 35970 33966 35982 34018
rect 36034 33966 36046 34018
rect 37202 33966 37214 34018
rect 37266 33966 37278 34018
rect 41682 33966 41694 34018
rect 41746 33966 41758 34018
rect 45938 33966 45950 34018
rect 46002 33966 46014 34018
rect 49074 33966 49086 34018
rect 49138 33966 49150 34018
rect 49858 33966 49870 34018
rect 49922 33966 49934 34018
rect 57362 33966 57374 34018
rect 57426 33966 57438 34018
rect 24446 33954 24498 33966
rect 55582 33954 55634 33966
rect 14478 33906 14530 33918
rect 14478 33842 14530 33854
rect 14814 33906 14866 33918
rect 14814 33842 14866 33854
rect 24334 33906 24386 33918
rect 24334 33842 24386 33854
rect 26014 33906 26066 33918
rect 26014 33842 26066 33854
rect 36430 33906 36482 33918
rect 38210 33854 38222 33906
rect 38274 33854 38286 33906
rect 51202 33854 51214 33906
rect 51266 33854 51278 33906
rect 36430 33842 36482 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 44046 33570 44098 33582
rect 44046 33506 44098 33518
rect 47182 33570 47234 33582
rect 47182 33506 47234 33518
rect 50094 33570 50146 33582
rect 50094 33506 50146 33518
rect 17278 33458 17330 33470
rect 14242 33406 14254 33458
rect 14306 33406 14318 33458
rect 16370 33406 16382 33458
rect 16434 33406 16446 33458
rect 17278 33394 17330 33406
rect 19406 33458 19458 33470
rect 29934 33458 29986 33470
rect 20066 33406 20078 33458
rect 20130 33406 20142 33458
rect 24434 33406 24446 33458
rect 24498 33406 24510 33458
rect 19406 33394 19458 33406
rect 29934 33394 29986 33406
rect 30382 33458 30434 33470
rect 30382 33394 30434 33406
rect 32734 33458 32786 33470
rect 42254 33458 42306 33470
rect 33506 33406 33518 33458
rect 33570 33406 33582 33458
rect 39890 33406 39902 33458
rect 39954 33406 39966 33458
rect 32734 33394 32786 33406
rect 42254 33394 42306 33406
rect 51214 33458 51266 33470
rect 57934 33458 57986 33470
rect 51650 33406 51662 33458
rect 51714 33406 51726 33458
rect 55794 33406 55806 33458
rect 55858 33406 55870 33458
rect 51214 33394 51266 33406
rect 57934 33394 57986 33406
rect 35758 33346 35810 33358
rect 13570 33294 13582 33346
rect 13634 33294 13646 33346
rect 18050 33294 18062 33346
rect 18114 33294 18126 33346
rect 18834 33294 18846 33346
rect 18898 33294 18910 33346
rect 22530 33294 22542 33346
rect 22594 33294 22606 33346
rect 23650 33294 23662 33346
rect 23714 33294 23726 33346
rect 29474 33294 29486 33346
rect 29538 33294 29550 33346
rect 35074 33294 35086 33346
rect 35138 33294 35150 33346
rect 35758 33282 35810 33294
rect 36318 33346 36370 33358
rect 43934 33346 43986 33358
rect 37090 33294 37102 33346
rect 37154 33294 37166 33346
rect 36318 33282 36370 33294
rect 43934 33282 43986 33294
rect 47070 33346 47122 33358
rect 47070 33282 47122 33294
rect 49982 33346 50034 33358
rect 49982 33282 50034 33294
rect 50878 33346 50930 33358
rect 51090 33294 51102 33346
rect 51154 33294 51166 33346
rect 53554 33294 53566 33346
rect 53618 33294 53630 33346
rect 54002 33294 54014 33346
rect 54066 33294 54078 33346
rect 55010 33294 55022 33346
rect 55074 33294 55086 33346
rect 50878 33282 50930 33294
rect 16830 33234 16882 33246
rect 22206 33234 22258 33246
rect 18722 33182 18734 33234
rect 18786 33182 18798 33234
rect 16830 33170 16882 33182
rect 22206 33170 22258 33182
rect 29150 33234 29202 33246
rect 29150 33170 29202 33182
rect 33070 33234 33122 33246
rect 36206 33234 36258 33246
rect 46510 33234 46562 33246
rect 34738 33182 34750 33234
rect 34802 33182 34814 33234
rect 35410 33182 35422 33234
rect 35474 33182 35486 33234
rect 37762 33182 37774 33234
rect 37826 33182 37838 33234
rect 33070 33170 33122 33182
rect 36206 33170 36258 33182
rect 46510 33170 46562 33182
rect 46734 33234 46786 33246
rect 46734 33170 46786 33182
rect 52110 33234 52162 33246
rect 52994 33182 53006 33234
rect 53058 33182 53070 33234
rect 54674 33182 54686 33234
rect 54738 33182 54750 33234
rect 52110 33170 52162 33182
rect 20526 33122 20578 33134
rect 17938 33070 17950 33122
rect 18002 33070 18014 33122
rect 20526 33058 20578 33070
rect 21422 33122 21474 33134
rect 21422 33058 21474 33070
rect 21870 33122 21922 33134
rect 21870 33058 21922 33070
rect 22318 33122 22370 33134
rect 22318 33058 22370 33070
rect 23326 33122 23378 33134
rect 29262 33122 29314 33134
rect 26674 33070 26686 33122
rect 26738 33070 26750 33122
rect 23326 33058 23378 33070
rect 29262 33058 29314 33070
rect 36430 33122 36482 33134
rect 36430 33058 36482 33070
rect 40350 33122 40402 33134
rect 40350 33058 40402 33070
rect 42814 33122 42866 33134
rect 42814 33058 42866 33070
rect 43262 33122 43314 33134
rect 43262 33058 43314 33070
rect 43822 33122 43874 33134
rect 43822 33058 43874 33070
rect 46622 33122 46674 33134
rect 46622 33058 46674 33070
rect 47182 33122 47234 33134
rect 54114 33070 54126 33122
rect 54178 33070 54190 33122
rect 47182 33058 47234 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 16382 32786 16434 32798
rect 16382 32722 16434 32734
rect 31950 32786 32002 32798
rect 31950 32722 32002 32734
rect 34078 32786 34130 32798
rect 34078 32722 34130 32734
rect 35646 32786 35698 32798
rect 35646 32722 35698 32734
rect 37326 32786 37378 32798
rect 43374 32786 43426 32798
rect 42130 32734 42142 32786
rect 42194 32734 42206 32786
rect 37326 32722 37378 32734
rect 43374 32722 43426 32734
rect 46398 32786 46450 32798
rect 46398 32722 46450 32734
rect 46846 32786 46898 32798
rect 46846 32722 46898 32734
rect 47182 32786 47234 32798
rect 56702 32786 56754 32798
rect 52210 32734 52222 32786
rect 52274 32734 52286 32786
rect 47182 32722 47234 32734
rect 56702 32722 56754 32734
rect 33742 32674 33794 32686
rect 29362 32622 29374 32674
rect 29426 32622 29438 32674
rect 33742 32610 33794 32622
rect 34302 32674 34354 32686
rect 34302 32610 34354 32622
rect 36878 32674 36930 32686
rect 36878 32610 36930 32622
rect 46958 32674 47010 32686
rect 46958 32610 47010 32622
rect 50094 32674 50146 32686
rect 50094 32610 50146 32622
rect 50206 32674 50258 32686
rect 50206 32610 50258 32622
rect 51662 32674 51714 32686
rect 51662 32610 51714 32622
rect 52782 32674 52834 32686
rect 52782 32610 52834 32622
rect 54798 32674 54850 32686
rect 54798 32610 54850 32622
rect 31278 32562 31330 32574
rect 12450 32510 12462 32562
rect 12514 32510 12526 32562
rect 18274 32510 18286 32562
rect 18338 32510 18350 32562
rect 23650 32510 23662 32562
rect 23714 32510 23726 32562
rect 24434 32510 24446 32562
rect 24498 32510 24510 32562
rect 30146 32510 30158 32562
rect 30210 32510 30222 32562
rect 30818 32510 30830 32562
rect 30882 32510 30894 32562
rect 31278 32498 31330 32510
rect 33966 32562 34018 32574
rect 33966 32498 34018 32510
rect 37102 32562 37154 32574
rect 37102 32498 37154 32510
rect 37438 32562 37490 32574
rect 37438 32498 37490 32510
rect 41806 32562 41858 32574
rect 41806 32498 41858 32510
rect 43710 32562 43762 32574
rect 43710 32498 43762 32510
rect 43934 32562 43986 32574
rect 43934 32498 43986 32510
rect 44382 32562 44434 32574
rect 46062 32562 46114 32574
rect 45826 32510 45838 32562
rect 45890 32510 45902 32562
rect 44382 32498 44434 32510
rect 46062 32498 46114 32510
rect 47518 32562 47570 32574
rect 49758 32562 49810 32574
rect 49298 32510 49310 32562
rect 49362 32510 49374 32562
rect 47518 32498 47570 32510
rect 49758 32498 49810 32510
rect 50766 32562 50818 32574
rect 50766 32498 50818 32510
rect 51774 32562 51826 32574
rect 54238 32562 54290 32574
rect 52098 32510 52110 32562
rect 52162 32510 52174 32562
rect 51774 32498 51826 32510
rect 54238 32498 54290 32510
rect 15822 32450 15874 32462
rect 33182 32450 33234 32462
rect 13122 32398 13134 32450
rect 13186 32398 13198 32450
rect 15250 32398 15262 32450
rect 15314 32398 15326 32450
rect 18946 32398 18958 32450
rect 19010 32398 19022 32450
rect 21074 32398 21086 32450
rect 21138 32398 21150 32450
rect 21522 32398 21534 32450
rect 21586 32398 21598 32450
rect 27234 32398 27246 32450
rect 27298 32398 27310 32450
rect 32386 32398 32398 32450
rect 32450 32398 32462 32450
rect 15822 32386 15874 32398
rect 33182 32386 33234 32398
rect 41582 32450 41634 32462
rect 41582 32386 41634 32398
rect 42926 32450 42978 32462
rect 42926 32386 42978 32398
rect 43822 32450 43874 32462
rect 43822 32386 43874 32398
rect 48862 32450 48914 32462
rect 48862 32386 48914 32398
rect 51326 32450 51378 32462
rect 51326 32386 51378 32398
rect 15934 32338 15986 32350
rect 15934 32274 15986 32286
rect 46286 32338 46338 32350
rect 46286 32274 46338 32286
rect 46510 32338 46562 32350
rect 46510 32274 46562 32286
rect 50206 32338 50258 32350
rect 50206 32274 50258 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 25342 32002 25394 32014
rect 38110 32002 38162 32014
rect 37538 31950 37550 32002
rect 37602 31950 37614 32002
rect 25342 31938 25394 31950
rect 38110 31938 38162 31950
rect 46958 32002 47010 32014
rect 50978 31950 50990 32002
rect 51042 31950 51054 32002
rect 46958 31938 47010 31950
rect 13918 31890 13970 31902
rect 14814 31890 14866 31902
rect 24894 31890 24946 31902
rect 26462 31890 26514 31902
rect 14466 31838 14478 31890
rect 14530 31838 14542 31890
rect 15586 31838 15598 31890
rect 15650 31838 15662 31890
rect 18946 31838 18958 31890
rect 19010 31838 19022 31890
rect 21858 31838 21870 31890
rect 21922 31838 21934 31890
rect 25666 31838 25678 31890
rect 25730 31838 25742 31890
rect 13918 31826 13970 31838
rect 14814 31826 14866 31838
rect 24894 31826 24946 31838
rect 26462 31826 26514 31838
rect 27358 31890 27410 31902
rect 27358 31826 27410 31838
rect 33630 31890 33682 31902
rect 33630 31826 33682 31838
rect 36206 31890 36258 31902
rect 44942 31890 44994 31902
rect 44258 31838 44270 31890
rect 44322 31838 44334 31890
rect 36206 31826 36258 31838
rect 44942 31826 44994 31838
rect 51998 31890 52050 31902
rect 53106 31838 53118 31890
rect 53170 31838 53182 31890
rect 55234 31838 55246 31890
rect 55298 31838 55310 31890
rect 57362 31838 57374 31890
rect 57426 31838 57438 31890
rect 51998 31826 52050 31838
rect 13806 31778 13858 31790
rect 15710 31778 15762 31790
rect 20526 31778 20578 31790
rect 30382 31778 30434 31790
rect 14130 31726 14142 31778
rect 14194 31726 14206 31778
rect 16482 31726 16494 31778
rect 16546 31726 16558 31778
rect 17490 31726 17502 31778
rect 17554 31726 17566 31778
rect 19058 31726 19070 31778
rect 19122 31726 19134 31778
rect 20066 31726 20078 31778
rect 20130 31726 20142 31778
rect 21298 31726 21310 31778
rect 21362 31726 21374 31778
rect 22642 31726 22654 31778
rect 22706 31726 22718 31778
rect 26674 31726 26686 31778
rect 26738 31726 26750 31778
rect 13806 31714 13858 31726
rect 15710 31714 15762 31726
rect 20526 31714 20578 31726
rect 30382 31714 30434 31726
rect 32174 31778 32226 31790
rect 33854 31778 33906 31790
rect 32722 31726 32734 31778
rect 32786 31726 32798 31778
rect 32174 31714 32226 31726
rect 33854 31714 33906 31726
rect 37326 31778 37378 31790
rect 46734 31778 46786 31790
rect 37538 31726 37550 31778
rect 37602 31726 37614 31778
rect 41458 31726 41470 31778
rect 41522 31726 41534 31778
rect 37326 31714 37378 31726
rect 46734 31714 46786 31726
rect 47182 31778 47234 31790
rect 47182 31714 47234 31726
rect 49086 31778 49138 31790
rect 52670 31778 52722 31790
rect 50978 31726 50990 31778
rect 51042 31726 51054 31778
rect 51314 31726 51326 31778
rect 51378 31726 51390 31778
rect 54002 31726 54014 31778
rect 54066 31726 54078 31778
rect 54786 31726 54798 31778
rect 54850 31726 54862 31778
rect 58034 31726 58046 31778
rect 58098 31726 58110 31778
rect 49086 31714 49138 31726
rect 52670 31714 52722 31726
rect 14590 31666 14642 31678
rect 14590 31602 14642 31614
rect 16158 31666 16210 31678
rect 18734 31666 18786 31678
rect 16594 31614 16606 31666
rect 16658 31614 16670 31666
rect 16158 31602 16210 31614
rect 18734 31602 18786 31614
rect 20414 31666 20466 31678
rect 20414 31602 20466 31614
rect 20750 31666 20802 31678
rect 22542 31666 22594 31678
rect 21522 31614 21534 31666
rect 21586 31614 21598 31666
rect 20750 31602 20802 31614
rect 22542 31602 22594 31614
rect 25006 31666 25058 31678
rect 25006 31602 25058 31614
rect 25566 31666 25618 31678
rect 25566 31602 25618 31614
rect 26014 31666 26066 31678
rect 31614 31666 31666 31678
rect 33182 31666 33234 31678
rect 34078 31666 34130 31678
rect 26226 31614 26238 31666
rect 26290 31614 26302 31666
rect 30034 31614 30046 31666
rect 30098 31614 30110 31666
rect 32498 31614 32510 31666
rect 32562 31614 32574 31666
rect 33394 31614 33406 31666
rect 33458 31614 33470 31666
rect 26014 31602 26066 31614
rect 31614 31602 31666 31614
rect 33182 31602 33234 31614
rect 34078 31602 34130 31614
rect 36990 31666 37042 31678
rect 36990 31602 37042 31614
rect 38222 31666 38274 31678
rect 38222 31602 38274 31614
rect 39678 31666 39730 31678
rect 39678 31602 39730 31614
rect 40014 31666 40066 31678
rect 47966 31666 48018 31678
rect 42130 31614 42142 31666
rect 42194 31614 42206 31666
rect 40014 31602 40066 31614
rect 47966 31602 48018 31614
rect 48190 31666 48242 31678
rect 48190 31602 48242 31614
rect 48414 31666 48466 31678
rect 48414 31602 48466 31614
rect 51550 31666 51602 31678
rect 51550 31602 51602 31614
rect 51886 31666 51938 31678
rect 54226 31614 54238 31666
rect 54290 31614 54302 31666
rect 51886 31602 51938 31614
rect 15598 31554 15650 31566
rect 15598 31490 15650 31502
rect 15934 31554 15986 31566
rect 17726 31554 17778 31566
rect 17602 31502 17614 31554
rect 17666 31502 17678 31554
rect 15934 31490 15986 31502
rect 17726 31490 17778 31502
rect 20302 31554 20354 31566
rect 33966 31554 34018 31566
rect 26450 31502 26462 31554
rect 26514 31502 26526 31554
rect 20302 31490 20354 31502
rect 33966 31490 34018 31502
rect 34526 31554 34578 31566
rect 34526 31490 34578 31502
rect 37102 31554 37154 31566
rect 37102 31490 37154 31502
rect 38670 31554 38722 31566
rect 38670 31490 38722 31502
rect 39342 31554 39394 31566
rect 39342 31490 39394 31502
rect 40350 31554 40402 31566
rect 40350 31490 40402 31502
rect 47630 31554 47682 31566
rect 47630 31490 47682 31502
rect 48302 31554 48354 31566
rect 49758 31554 49810 31566
rect 48738 31502 48750 31554
rect 48802 31502 48814 31554
rect 48302 31490 48354 31502
rect 49758 31490 49810 31502
rect 49982 31554 50034 31566
rect 49982 31490 50034 31502
rect 50094 31554 50146 31566
rect 50094 31490 50146 31502
rect 50206 31554 50258 31566
rect 50206 31490 50258 31502
rect 51438 31554 51490 31566
rect 54562 31502 54574 31554
rect 54626 31502 54638 31554
rect 51438 31490 51490 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 13246 31218 13298 31230
rect 13246 31154 13298 31166
rect 24670 31218 24722 31230
rect 24670 31154 24722 31166
rect 29710 31218 29762 31230
rect 29710 31154 29762 31166
rect 40014 31218 40066 31230
rect 40014 31154 40066 31166
rect 40910 31218 40962 31230
rect 40910 31154 40962 31166
rect 41806 31218 41858 31230
rect 41806 31154 41858 31166
rect 43150 31218 43202 31230
rect 44270 31218 44322 31230
rect 43474 31166 43486 31218
rect 43538 31166 43550 31218
rect 43150 31154 43202 31166
rect 44270 31154 44322 31166
rect 45502 31218 45554 31230
rect 45502 31154 45554 31166
rect 49422 31218 49474 31230
rect 49422 31154 49474 31166
rect 13470 31106 13522 31118
rect 13470 31042 13522 31054
rect 13806 31106 13858 31118
rect 13806 31042 13858 31054
rect 29150 31106 29202 31118
rect 29150 31042 29202 31054
rect 30158 31106 30210 31118
rect 39902 31106 39954 31118
rect 33842 31054 33854 31106
rect 33906 31054 33918 31106
rect 37090 31054 37102 31106
rect 37154 31054 37166 31106
rect 30158 31042 30210 31054
rect 39902 31042 39954 31054
rect 40126 31106 40178 31118
rect 42590 31106 42642 31118
rect 42130 31054 42142 31106
rect 42194 31054 42206 31106
rect 40126 31042 40178 31054
rect 42590 31042 42642 31054
rect 42814 31106 42866 31118
rect 42814 31042 42866 31054
rect 44158 31106 44210 31118
rect 44158 31042 44210 31054
rect 44718 31106 44770 31118
rect 44718 31042 44770 31054
rect 50542 31106 50594 31118
rect 50542 31042 50594 31054
rect 51886 31106 51938 31118
rect 51886 31042 51938 31054
rect 52110 31106 52162 31118
rect 52110 31042 52162 31054
rect 30046 30994 30098 31006
rect 44942 30994 44994 31006
rect 14130 30942 14142 30994
rect 14194 30942 14206 30994
rect 15810 30942 15822 30994
rect 15874 30942 15886 30994
rect 16146 30942 16158 30994
rect 16210 30942 16222 30994
rect 17826 30942 17838 30994
rect 17890 30942 17902 30994
rect 18722 30942 18734 30994
rect 18786 30942 18798 30994
rect 21410 30942 21422 30994
rect 21474 30942 21486 30994
rect 22978 30942 22990 30994
rect 23042 30942 23054 30994
rect 28018 30942 28030 30994
rect 28082 30942 28094 30994
rect 33058 30942 33070 30994
rect 33122 30942 33134 30994
rect 36418 30942 36430 30994
rect 36482 30942 36494 30994
rect 44370 30942 44382 30994
rect 44434 30942 44446 30994
rect 30046 30930 30098 30942
rect 44942 30930 44994 30942
rect 45278 30994 45330 31006
rect 45278 30930 45330 30942
rect 45614 30994 45666 31006
rect 47406 30994 47458 31006
rect 46498 30942 46510 30994
rect 46562 30942 46574 30994
rect 45614 30930 45666 30942
rect 47406 30930 47458 30942
rect 49198 30994 49250 31006
rect 49198 30930 49250 30942
rect 49422 30994 49474 31006
rect 49422 30930 49474 30942
rect 49758 30994 49810 31006
rect 49758 30930 49810 30942
rect 50094 30994 50146 31006
rect 50094 30930 50146 30942
rect 50206 30994 50258 31006
rect 50206 30930 50258 30942
rect 52558 30994 52610 31006
rect 54910 30994 54962 31006
rect 53778 30942 53790 30994
rect 53842 30942 53854 30994
rect 52558 30930 52610 30942
rect 54910 30930 54962 30942
rect 55358 30994 55410 31006
rect 55358 30930 55410 30942
rect 17390 30882 17442 30894
rect 19070 30882 19122 30894
rect 30718 30882 30770 30894
rect 46734 30882 46786 30894
rect 16818 30830 16830 30882
rect 16882 30830 16894 30882
rect 18274 30830 18286 30882
rect 18338 30830 18350 30882
rect 22082 30830 22094 30882
rect 22146 30830 22158 30882
rect 23314 30830 23326 30882
rect 23378 30830 23390 30882
rect 25218 30830 25230 30882
rect 25282 30830 25294 30882
rect 27346 30830 27358 30882
rect 27410 30830 27422 30882
rect 35970 30830 35982 30882
rect 36034 30830 36046 30882
rect 39218 30830 39230 30882
rect 39282 30830 39294 30882
rect 41346 30830 41358 30882
rect 41410 30830 41422 30882
rect 42466 30830 42478 30882
rect 42530 30830 42542 30882
rect 17390 30818 17442 30830
rect 19070 30818 19122 30830
rect 30718 30818 30770 30830
rect 46734 30818 46786 30830
rect 47966 30882 48018 30894
rect 47966 30818 48018 30830
rect 50430 30882 50482 30894
rect 50430 30818 50482 30830
rect 50990 30882 51042 30894
rect 50990 30818 51042 30830
rect 52334 30882 52386 30894
rect 52770 30830 52782 30882
rect 52834 30830 52846 30882
rect 53890 30830 53902 30882
rect 53954 30830 53966 30882
rect 52334 30818 52386 30830
rect 13134 30770 13186 30782
rect 13134 30706 13186 30718
rect 14142 30770 14194 30782
rect 14142 30706 14194 30718
rect 18734 30770 18786 30782
rect 24110 30770 24162 30782
rect 21970 30718 21982 30770
rect 22034 30718 22046 30770
rect 18734 30706 18786 30718
rect 24110 30706 24162 30718
rect 29262 30770 29314 30782
rect 29262 30706 29314 30718
rect 30158 30770 30210 30782
rect 30158 30706 30210 30718
rect 30606 30770 30658 30782
rect 30606 30706 30658 30718
rect 45054 30770 45106 30782
rect 45054 30706 45106 30718
rect 46958 30770 47010 30782
rect 46958 30706 47010 30718
rect 47070 30770 47122 30782
rect 47070 30706 47122 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 21310 30434 21362 30446
rect 18610 30382 18622 30434
rect 18674 30382 18686 30434
rect 21310 30370 21362 30382
rect 22766 30434 22818 30446
rect 39006 30434 39058 30446
rect 26338 30382 26350 30434
rect 26402 30382 26414 30434
rect 22766 30370 22818 30382
rect 39006 30370 39058 30382
rect 47742 30322 47794 30334
rect 11778 30270 11790 30322
rect 11842 30270 11854 30322
rect 47742 30258 47794 30270
rect 53454 30322 53506 30334
rect 53454 30258 53506 30270
rect 53678 30322 53730 30334
rect 54562 30270 54574 30322
rect 54626 30270 54638 30322
rect 53678 30258 53730 30270
rect 12238 30210 12290 30222
rect 8978 30158 8990 30210
rect 9042 30158 9054 30210
rect 12238 30146 12290 30158
rect 16718 30210 16770 30222
rect 16718 30146 16770 30158
rect 17166 30210 17218 30222
rect 22094 30210 22146 30222
rect 17378 30158 17390 30210
rect 17442 30158 17454 30210
rect 18610 30158 18622 30210
rect 18674 30158 18686 30210
rect 19506 30158 19518 30210
rect 19570 30158 19582 30210
rect 21634 30158 21646 30210
rect 21698 30158 21710 30210
rect 21858 30158 21870 30210
rect 21922 30158 21934 30210
rect 17166 30146 17218 30158
rect 22094 30146 22146 30158
rect 22430 30210 22482 30222
rect 22430 30146 22482 30158
rect 25790 30210 25842 30222
rect 25790 30146 25842 30158
rect 26126 30210 26178 30222
rect 28366 30210 28418 30222
rect 26562 30158 26574 30210
rect 26626 30158 26638 30210
rect 27122 30158 27134 30210
rect 27186 30158 27198 30210
rect 26126 30146 26178 30158
rect 28366 30146 28418 30158
rect 28702 30210 28754 30222
rect 28702 30146 28754 30158
rect 29038 30210 29090 30222
rect 29038 30146 29090 30158
rect 29486 30210 29538 30222
rect 29486 30146 29538 30158
rect 29598 30210 29650 30222
rect 35758 30210 35810 30222
rect 31042 30158 31054 30210
rect 31106 30158 31118 30210
rect 29598 30146 29650 30158
rect 35758 30146 35810 30158
rect 35870 30210 35922 30222
rect 39230 30210 39282 30222
rect 37426 30158 37438 30210
rect 37490 30158 37502 30210
rect 38210 30158 38222 30210
rect 38274 30158 38286 30210
rect 38658 30158 38670 30210
rect 38722 30158 38734 30210
rect 35870 30146 35922 30158
rect 39230 30146 39282 30158
rect 39790 30210 39842 30222
rect 39790 30146 39842 30158
rect 40238 30210 40290 30222
rect 40238 30146 40290 30158
rect 41134 30210 41186 30222
rect 41134 30146 41186 30158
rect 41694 30210 41746 30222
rect 41694 30146 41746 30158
rect 42030 30210 42082 30222
rect 42030 30146 42082 30158
rect 42590 30210 42642 30222
rect 46398 30210 46450 30222
rect 43026 30158 43038 30210
rect 43090 30158 43102 30210
rect 42590 30146 42642 30158
rect 46398 30146 46450 30158
rect 47070 30210 47122 30222
rect 47070 30146 47122 30158
rect 47854 30210 47906 30222
rect 47854 30146 47906 30158
rect 49534 30210 49586 30222
rect 49534 30146 49586 30158
rect 51886 30210 51938 30222
rect 56690 30158 56702 30210
rect 56754 30158 56766 30210
rect 57362 30158 57374 30210
rect 57426 30158 57438 30210
rect 51886 30146 51938 30158
rect 15710 30098 15762 30110
rect 9650 30046 9662 30098
rect 9714 30046 9726 30098
rect 15710 30034 15762 30046
rect 16606 30098 16658 30110
rect 21422 30098 21474 30110
rect 20066 30046 20078 30098
rect 20130 30046 20142 30098
rect 16606 30034 16658 30046
rect 21422 30034 21474 30046
rect 22318 30098 22370 30110
rect 22318 30034 22370 30046
rect 22878 30098 22930 30110
rect 28478 30098 28530 30110
rect 37662 30098 37714 30110
rect 47294 30098 47346 30110
rect 49870 30098 49922 30110
rect 26898 30046 26910 30098
rect 26962 30046 26974 30098
rect 34402 30046 34414 30098
rect 34466 30046 34478 30098
rect 46050 30046 46062 30098
rect 46114 30046 46126 30098
rect 48850 30046 48862 30098
rect 48914 30046 48926 30098
rect 22878 30034 22930 30046
rect 28478 30034 28530 30046
rect 37662 30034 37714 30046
rect 47294 30034 47346 30046
rect 49870 30034 49922 30046
rect 52110 30098 52162 30110
rect 52110 30034 52162 30046
rect 53006 30098 53058 30110
rect 53006 30034 53058 30046
rect 15934 29986 15986 29998
rect 15934 29922 15986 29934
rect 16046 29986 16098 29998
rect 16046 29922 16098 29934
rect 16158 29986 16210 29998
rect 16158 29922 16210 29934
rect 16494 29986 16546 29998
rect 16494 29922 16546 29934
rect 26574 29986 26626 29998
rect 26574 29922 26626 29934
rect 29262 29986 29314 29998
rect 29262 29922 29314 29934
rect 40574 29986 40626 29998
rect 45726 29986 45778 29998
rect 47630 29986 47682 29998
rect 43250 29934 43262 29986
rect 43314 29934 43326 29986
rect 46722 29934 46734 29986
rect 46786 29934 46798 29986
rect 40574 29922 40626 29934
rect 45726 29922 45778 29934
rect 47630 29922 47682 29934
rect 48078 29986 48130 29998
rect 48078 29922 48130 29934
rect 48526 29986 48578 29998
rect 48526 29922 48578 29934
rect 49422 29986 49474 29998
rect 49422 29922 49474 29934
rect 49646 29986 49698 29998
rect 52782 29986 52834 29998
rect 51538 29934 51550 29986
rect 51602 29934 51614 29986
rect 49646 29922 49698 29934
rect 52782 29922 52834 29934
rect 52894 29986 52946 29998
rect 54002 29934 54014 29986
rect 54066 29934 54078 29986
rect 52894 29922 52946 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 9774 29650 9826 29662
rect 9774 29586 9826 29598
rect 19406 29650 19458 29662
rect 19406 29586 19458 29598
rect 27694 29650 27746 29662
rect 35198 29650 35250 29662
rect 31938 29598 31950 29650
rect 32002 29598 32014 29650
rect 27694 29586 27746 29598
rect 35198 29586 35250 29598
rect 41022 29650 41074 29662
rect 41022 29586 41074 29598
rect 46958 29650 47010 29662
rect 46958 29586 47010 29598
rect 47406 29650 47458 29662
rect 47406 29586 47458 29598
rect 49310 29650 49362 29662
rect 49310 29586 49362 29598
rect 18846 29538 18898 29550
rect 12898 29486 12910 29538
rect 12962 29486 12974 29538
rect 18050 29486 18062 29538
rect 18114 29486 18126 29538
rect 18846 29474 18898 29486
rect 23662 29538 23714 29550
rect 34526 29538 34578 29550
rect 46062 29538 46114 29550
rect 28802 29486 28814 29538
rect 28866 29486 28878 29538
rect 39890 29486 39902 29538
rect 39954 29486 39966 29538
rect 50418 29486 50430 29538
rect 50482 29486 50494 29538
rect 23662 29474 23714 29486
rect 34526 29474 34578 29486
rect 46062 29474 46114 29486
rect 10110 29426 10162 29438
rect 23998 29426 24050 29438
rect 32286 29426 32338 29438
rect 5730 29374 5742 29426
rect 5794 29374 5806 29426
rect 12226 29374 12238 29426
rect 12290 29374 12302 29426
rect 17378 29374 17390 29426
rect 17442 29374 17454 29426
rect 17938 29374 17950 29426
rect 18002 29374 18014 29426
rect 22082 29374 22094 29426
rect 22146 29374 22158 29426
rect 24658 29374 24670 29426
rect 24722 29374 24734 29426
rect 25890 29374 25902 29426
rect 25954 29374 25966 29426
rect 28018 29374 28030 29426
rect 28082 29374 28094 29426
rect 10110 29362 10162 29374
rect 23998 29362 24050 29374
rect 32286 29362 32338 29374
rect 33070 29426 33122 29438
rect 33966 29426 34018 29438
rect 33730 29374 33742 29426
rect 33794 29374 33806 29426
rect 33070 29362 33122 29374
rect 33966 29362 34018 29374
rect 34750 29426 34802 29438
rect 34750 29362 34802 29374
rect 34974 29426 35026 29438
rect 34974 29362 35026 29374
rect 35310 29426 35362 29438
rect 45166 29426 45218 29438
rect 40114 29374 40126 29426
rect 40178 29374 40190 29426
rect 35310 29362 35362 29374
rect 45166 29362 45218 29374
rect 45390 29426 45442 29438
rect 45390 29362 45442 29374
rect 45838 29426 45890 29438
rect 45838 29362 45890 29374
rect 46398 29426 46450 29438
rect 46398 29362 46450 29374
rect 46622 29426 46674 29438
rect 46622 29362 46674 29374
rect 47070 29426 47122 29438
rect 47070 29362 47122 29374
rect 47182 29426 47234 29438
rect 47182 29362 47234 29374
rect 49086 29426 49138 29438
rect 49086 29362 49138 29374
rect 49198 29426 49250 29438
rect 49198 29362 49250 29374
rect 49534 29426 49586 29438
rect 53902 29426 53954 29438
rect 55358 29426 55410 29438
rect 50082 29374 50094 29426
rect 50146 29374 50158 29426
rect 51650 29374 51662 29426
rect 51714 29374 51726 29426
rect 53218 29374 53230 29426
rect 53282 29374 53294 29426
rect 54786 29374 54798 29426
rect 54850 29374 54862 29426
rect 49534 29362 49586 29374
rect 53902 29362 53954 29374
rect 55358 29362 55410 29374
rect 8990 29314 9042 29326
rect 15486 29314 15538 29326
rect 22766 29314 22818 29326
rect 6402 29262 6414 29314
rect 6466 29262 6478 29314
rect 8530 29262 8542 29314
rect 8594 29262 8606 29314
rect 15026 29262 15038 29314
rect 15090 29262 15102 29314
rect 18386 29262 18398 29314
rect 18450 29262 18462 29314
rect 21970 29262 21982 29314
rect 22034 29262 22046 29314
rect 8990 29250 9042 29262
rect 15486 29250 15538 29262
rect 22766 29250 22818 29262
rect 25230 29314 25282 29326
rect 32510 29314 32562 29326
rect 44494 29314 44546 29326
rect 25554 29262 25566 29314
rect 25618 29262 25630 29314
rect 30930 29262 30942 29314
rect 30994 29262 31006 29314
rect 34402 29262 34414 29314
rect 34466 29262 34478 29314
rect 25230 29250 25282 29262
rect 32510 29250 32562 29262
rect 44494 29250 44546 29262
rect 44830 29314 44882 29326
rect 44830 29250 44882 29262
rect 45614 29314 45666 29326
rect 45614 29250 45666 29262
rect 46174 29314 46226 29326
rect 50866 29262 50878 29314
rect 50930 29262 50942 29314
rect 54338 29262 54350 29314
rect 54402 29262 54414 29314
rect 46174 29250 46226 29262
rect 24334 29202 24386 29214
rect 24334 29138 24386 29150
rect 24670 29202 24722 29214
rect 24670 29138 24722 29150
rect 55134 29202 55186 29214
rect 55134 29138 55186 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 10558 28866 10610 28878
rect 10558 28802 10610 28814
rect 18286 28866 18338 28878
rect 18286 28802 18338 28814
rect 21310 28866 21362 28878
rect 21310 28802 21362 28814
rect 27582 28866 27634 28878
rect 27582 28802 27634 28814
rect 28254 28866 28306 28878
rect 28254 28802 28306 28814
rect 29150 28866 29202 28878
rect 29150 28802 29202 28814
rect 45166 28866 45218 28878
rect 53218 28814 53230 28866
rect 53282 28814 53294 28866
rect 45166 28802 45218 28814
rect 16830 28754 16882 28766
rect 30046 28754 30098 28766
rect 33406 28754 33458 28766
rect 36318 28754 36370 28766
rect 14242 28702 14254 28754
rect 14306 28702 14318 28754
rect 16370 28702 16382 28754
rect 16434 28702 16446 28754
rect 25330 28702 25342 28754
rect 25394 28702 25406 28754
rect 28578 28702 28590 28754
rect 28642 28702 28654 28754
rect 32162 28702 32174 28754
rect 32226 28702 32238 28754
rect 35074 28702 35086 28754
rect 35138 28702 35150 28754
rect 16830 28690 16882 28702
rect 30046 28690 30098 28702
rect 33406 28690 33458 28702
rect 36318 28690 36370 28702
rect 37662 28754 37714 28766
rect 37662 28690 37714 28702
rect 38110 28754 38162 28766
rect 41918 28754 41970 28766
rect 38546 28702 38558 28754
rect 38610 28702 38622 28754
rect 38110 28690 38162 28702
rect 41918 28690 41970 28702
rect 42366 28754 42418 28766
rect 42366 28690 42418 28702
rect 43374 28754 43426 28766
rect 43374 28690 43426 28702
rect 43822 28754 43874 28766
rect 43822 28690 43874 28702
rect 44270 28754 44322 28766
rect 49298 28702 49310 28754
rect 49362 28702 49374 28754
rect 51426 28702 51438 28754
rect 51490 28702 51502 28754
rect 52098 28702 52110 28754
rect 52162 28702 52174 28754
rect 53106 28702 53118 28754
rect 53170 28702 53182 28754
rect 54898 28702 54910 28754
rect 54962 28702 54974 28754
rect 44270 28690 44322 28702
rect 7086 28642 7138 28654
rect 7086 28578 7138 28590
rect 7534 28642 7586 28654
rect 7534 28578 7586 28590
rect 7870 28642 7922 28654
rect 7870 28578 7922 28590
rect 10894 28642 10946 28654
rect 21646 28642 21698 28654
rect 33294 28642 33346 28654
rect 11554 28590 11566 28642
rect 11618 28590 11630 28642
rect 13458 28590 13470 28642
rect 13522 28590 13534 28642
rect 23426 28590 23438 28642
rect 23490 28590 23502 28642
rect 24882 28590 24894 28642
rect 24946 28590 24958 28642
rect 25218 28590 25230 28642
rect 25282 28590 25294 28642
rect 27346 28590 27358 28642
rect 27410 28590 27422 28642
rect 27906 28590 27918 28642
rect 27970 28590 27982 28642
rect 29474 28590 29486 28642
rect 29538 28590 29550 28642
rect 32274 28590 32286 28642
rect 32338 28590 32350 28642
rect 10894 28578 10946 28590
rect 21646 28578 21698 28590
rect 33294 28578 33346 28590
rect 33630 28642 33682 28654
rect 33630 28578 33682 28590
rect 33854 28642 33906 28654
rect 33854 28578 33906 28590
rect 34078 28642 34130 28654
rect 34078 28578 34130 28590
rect 34414 28642 34466 28654
rect 34414 28578 34466 28590
rect 34750 28642 34802 28654
rect 42926 28642 42978 28654
rect 37202 28590 37214 28642
rect 37266 28590 37278 28642
rect 41458 28590 41470 28642
rect 41522 28590 41534 28642
rect 45602 28590 45614 28642
rect 45666 28590 45678 28642
rect 46834 28590 46846 28642
rect 46898 28590 46910 28642
rect 47618 28590 47630 28642
rect 47682 28590 47694 28642
rect 48514 28590 48526 28642
rect 48578 28590 48590 28642
rect 52994 28590 53006 28642
rect 53058 28590 53070 28642
rect 53778 28590 53790 28642
rect 53842 28590 53854 28642
rect 54226 28590 54238 28642
rect 54290 28590 54302 28642
rect 55346 28590 55358 28642
rect 55410 28590 55422 28642
rect 55682 28590 55694 28642
rect 55746 28590 55758 28642
rect 56466 28590 56478 28642
rect 56530 28590 56542 28642
rect 34750 28578 34802 28590
rect 42926 28578 42978 28590
rect 6750 28530 6802 28542
rect 18398 28530 18450 28542
rect 27134 28530 27186 28542
rect 8082 28478 8094 28530
rect 8146 28478 8158 28530
rect 8642 28478 8654 28530
rect 8706 28478 8718 28530
rect 11666 28478 11678 28530
rect 11730 28478 11742 28530
rect 26226 28478 26238 28530
rect 26290 28478 26302 28530
rect 6750 28466 6802 28478
rect 18398 28466 18450 28478
rect 27134 28466 27186 28478
rect 28478 28530 28530 28542
rect 28478 28466 28530 28478
rect 32958 28530 33010 28542
rect 32958 28466 33010 28478
rect 35534 28530 35586 28542
rect 45054 28530 45106 28542
rect 51774 28530 51826 28542
rect 40674 28478 40686 28530
rect 40738 28478 40750 28530
rect 46610 28478 46622 28530
rect 46674 28478 46686 28530
rect 47282 28478 47294 28530
rect 47346 28478 47358 28530
rect 55010 28478 55022 28530
rect 55074 28478 55086 28530
rect 56242 28478 56254 28530
rect 56306 28478 56318 28530
rect 35534 28466 35586 28478
rect 45054 28466 45106 28478
rect 51774 28466 51826 28478
rect 19630 28418 19682 28430
rect 19630 28354 19682 28366
rect 21422 28418 21474 28430
rect 21422 28354 21474 28366
rect 22878 28418 22930 28430
rect 29262 28418 29314 28430
rect 27570 28366 27582 28418
rect 27634 28366 27646 28418
rect 22878 28354 22930 28366
rect 29262 28354 29314 28366
rect 34302 28418 34354 28430
rect 34302 28354 34354 28366
rect 35086 28418 35138 28430
rect 35086 28354 35138 28366
rect 35310 28418 35362 28430
rect 35310 28354 35362 28366
rect 42254 28418 42306 28430
rect 42254 28354 42306 28366
rect 42478 28418 42530 28430
rect 48190 28418 48242 28430
rect 46946 28366 46958 28418
rect 47010 28366 47022 28418
rect 42478 28354 42530 28366
rect 48190 28354 48242 28366
rect 51998 28418 52050 28430
rect 51998 28354 52050 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 12910 28082 12962 28094
rect 12910 28018 12962 28030
rect 17502 28082 17554 28094
rect 17502 28018 17554 28030
rect 19070 28082 19122 28094
rect 32174 28082 32226 28094
rect 31826 28030 31838 28082
rect 31890 28030 31902 28082
rect 19070 28018 19122 28030
rect 32174 28018 32226 28030
rect 32398 28082 32450 28094
rect 32398 28018 32450 28030
rect 41022 28082 41074 28094
rect 41022 28018 41074 28030
rect 47742 28082 47794 28094
rect 47742 28018 47794 28030
rect 48862 28082 48914 28094
rect 48862 28018 48914 28030
rect 49534 28082 49586 28094
rect 49534 28018 49586 28030
rect 8878 27970 8930 27982
rect 38446 27970 38498 27982
rect 8194 27918 8206 27970
rect 8258 27918 8270 27970
rect 14466 27918 14478 27970
rect 14530 27918 14542 27970
rect 20402 27918 20414 27970
rect 20466 27918 20478 27970
rect 27682 27918 27694 27970
rect 27746 27918 27758 27970
rect 36530 27918 36542 27970
rect 36594 27918 36606 27970
rect 8878 27906 8930 27918
rect 38446 27906 38498 27918
rect 39678 27970 39730 27982
rect 49982 27970 50034 27982
rect 42354 27918 42366 27970
rect 42418 27918 42430 27970
rect 39678 27906 39730 27918
rect 49982 27906 50034 27918
rect 51774 27970 51826 27982
rect 51774 27906 51826 27918
rect 53902 27970 53954 27982
rect 54114 27918 54126 27970
rect 54178 27918 54190 27970
rect 56578 27918 56590 27970
rect 56642 27918 56654 27970
rect 53902 27906 53954 27918
rect 7646 27858 7698 27870
rect 32510 27858 32562 27870
rect 38558 27858 38610 27870
rect 47854 27858 47906 27870
rect 4050 27806 4062 27858
rect 4114 27806 4126 27858
rect 8082 27806 8094 27858
rect 8146 27806 8158 27858
rect 9538 27806 9550 27858
rect 9602 27806 9614 27858
rect 13794 27806 13806 27858
rect 13858 27806 13870 27858
rect 19730 27806 19742 27858
rect 19794 27806 19806 27858
rect 23986 27806 23998 27858
rect 24050 27806 24062 27858
rect 24322 27806 24334 27858
rect 24386 27806 24398 27858
rect 28354 27806 28366 27858
rect 28418 27806 28430 27858
rect 28802 27806 28814 27858
rect 28866 27806 28878 27858
rect 33170 27806 33182 27858
rect 33234 27806 33246 27858
rect 36418 27806 36430 27858
rect 36482 27806 36494 27858
rect 41682 27806 41694 27858
rect 41746 27806 41758 27858
rect 44818 27806 44830 27858
rect 44882 27806 44894 27858
rect 7646 27794 7698 27806
rect 32510 27794 32562 27806
rect 38558 27794 38610 27806
rect 47854 27794 47906 27806
rect 48974 27858 49026 27870
rect 53454 27858 53506 27870
rect 50418 27806 50430 27858
rect 50482 27806 50494 27858
rect 51650 27806 51662 27858
rect 51714 27806 51726 27858
rect 52322 27806 52334 27858
rect 52386 27806 52398 27858
rect 52770 27806 52782 27858
rect 52834 27806 52846 27858
rect 48974 27794 49026 27806
rect 53454 27794 53506 27806
rect 55022 27858 55074 27870
rect 55022 27794 55074 27806
rect 55582 27858 55634 27870
rect 56802 27806 56814 27858
rect 56866 27806 56878 27858
rect 55582 27794 55634 27806
rect 22990 27746 23042 27758
rect 54238 27746 54290 27758
rect 4722 27694 4734 27746
rect 4786 27694 4798 27746
rect 6850 27694 6862 27746
rect 6914 27694 6926 27746
rect 10322 27694 10334 27746
rect 10386 27694 10398 27746
rect 12450 27694 12462 27746
rect 12514 27694 12526 27746
rect 16594 27694 16606 27746
rect 16658 27694 16670 27746
rect 22530 27694 22542 27746
rect 22594 27694 22606 27746
rect 24098 27694 24110 27746
rect 24162 27694 24174 27746
rect 24546 27694 24558 27746
rect 24610 27694 24622 27746
rect 25554 27694 25566 27746
rect 25618 27694 25630 27746
rect 29586 27694 29598 27746
rect 29650 27694 29662 27746
rect 33954 27694 33966 27746
rect 34018 27694 34030 27746
rect 36082 27694 36094 27746
rect 36146 27694 36158 27746
rect 40898 27694 40910 27746
rect 40962 27694 40974 27746
rect 44482 27694 44494 27746
rect 44546 27694 44558 27746
rect 46274 27694 46286 27746
rect 46338 27694 46350 27746
rect 50754 27694 50766 27746
rect 50818 27694 50830 27746
rect 22990 27682 23042 27694
rect 54238 27682 54290 27694
rect 7310 27634 7362 27646
rect 7310 27570 7362 27582
rect 8990 27634 9042 27646
rect 8990 27570 9042 27582
rect 18958 27634 19010 27646
rect 18958 27570 19010 27582
rect 19294 27634 19346 27646
rect 19294 27570 19346 27582
rect 41246 27634 41298 27646
rect 41246 27570 41298 27582
rect 49086 27634 49138 27646
rect 53230 27634 53282 27646
rect 52210 27582 52222 27634
rect 52274 27582 52286 27634
rect 49086 27570 49138 27582
rect 53230 27570 53282 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 33742 27298 33794 27310
rect 33742 27234 33794 27246
rect 42366 27298 42418 27310
rect 42366 27234 42418 27246
rect 45054 27298 45106 27310
rect 53218 27246 53230 27298
rect 53282 27246 53294 27298
rect 45054 27234 45106 27246
rect 7534 27186 7586 27198
rect 7534 27122 7586 27134
rect 11118 27186 11170 27198
rect 19630 27186 19682 27198
rect 17154 27134 17166 27186
rect 17218 27134 17230 27186
rect 19282 27134 19294 27186
rect 19346 27134 19358 27186
rect 11118 27122 11170 27134
rect 19630 27122 19682 27134
rect 21310 27186 21362 27198
rect 28478 27186 28530 27198
rect 26338 27134 26350 27186
rect 26402 27134 26414 27186
rect 21310 27122 21362 27134
rect 28478 27122 28530 27134
rect 31502 27186 31554 27198
rect 32958 27186 33010 27198
rect 32162 27134 32174 27186
rect 32226 27134 32238 27186
rect 31502 27122 31554 27134
rect 32958 27122 33010 27134
rect 37326 27186 37378 27198
rect 37326 27122 37378 27134
rect 40014 27186 40066 27198
rect 40014 27122 40066 27134
rect 40462 27186 40514 27198
rect 40462 27122 40514 27134
rect 41806 27186 41858 27198
rect 41806 27122 41858 27134
rect 43598 27186 43650 27198
rect 43598 27122 43650 27134
rect 44830 27186 44882 27198
rect 44830 27122 44882 27134
rect 45390 27186 45442 27198
rect 52782 27186 52834 27198
rect 47394 27134 47406 27186
rect 47458 27134 47470 27186
rect 55570 27134 55582 27186
rect 55634 27134 55646 27186
rect 57698 27134 57710 27186
rect 57762 27134 57774 27186
rect 45390 27122 45442 27134
rect 52782 27122 52834 27134
rect 5966 27074 6018 27086
rect 5966 27010 6018 27022
rect 9998 27074 10050 27086
rect 9998 27010 10050 27022
rect 10782 27074 10834 27086
rect 20526 27074 20578 27086
rect 22206 27074 22258 27086
rect 11554 27022 11566 27074
rect 11618 27022 11630 27074
rect 16370 27022 16382 27074
rect 16434 27022 16446 27074
rect 20066 27022 20078 27074
rect 20130 27022 20142 27074
rect 21746 27022 21758 27074
rect 21810 27022 21822 27074
rect 10782 27010 10834 27022
rect 20526 27010 20578 27022
rect 22206 27010 22258 27022
rect 22542 27074 22594 27086
rect 31614 27074 31666 27086
rect 33294 27074 33346 27086
rect 23090 27022 23102 27074
rect 23154 27022 23166 27074
rect 23426 27022 23438 27074
rect 23490 27022 23502 27074
rect 32274 27022 32286 27074
rect 32338 27022 32350 27074
rect 22542 27010 22594 27022
rect 31614 27010 31666 27022
rect 33294 27010 33346 27022
rect 33518 27074 33570 27086
rect 34302 27074 34354 27086
rect 35982 27074 36034 27086
rect 33954 27022 33966 27074
rect 34018 27022 34030 27074
rect 34738 27022 34750 27074
rect 34802 27022 34814 27074
rect 35634 27022 35646 27074
rect 35698 27022 35710 27074
rect 33518 27010 33570 27022
rect 34302 27010 34354 27022
rect 35982 27010 36034 27022
rect 36430 27074 36482 27086
rect 38782 27074 38834 27086
rect 38322 27022 38334 27074
rect 38386 27022 38398 27074
rect 36430 27010 36482 27022
rect 38782 27010 38834 27022
rect 39230 27074 39282 27086
rect 39230 27010 39282 27022
rect 41918 27074 41970 27086
rect 41918 27010 41970 27022
rect 42142 27074 42194 27086
rect 42142 27010 42194 27022
rect 42814 27074 42866 27086
rect 42814 27010 42866 27022
rect 43262 27074 43314 27086
rect 43262 27010 43314 27022
rect 44158 27074 44210 27086
rect 51774 27074 51826 27086
rect 45714 27022 45726 27074
rect 45778 27022 45790 27074
rect 48738 27022 48750 27074
rect 48802 27022 48814 27074
rect 49634 27022 49646 27074
rect 49698 27022 49710 27074
rect 50530 27022 50542 27074
rect 50594 27022 50606 27074
rect 51426 27022 51438 27074
rect 51490 27022 51502 27074
rect 44158 27010 44210 27022
rect 51774 27010 51826 27022
rect 53678 27074 53730 27086
rect 53678 27010 53730 27022
rect 53790 27074 53842 27086
rect 54002 27022 54014 27074
rect 54066 27022 54078 27074
rect 54898 27022 54910 27074
rect 54962 27022 54974 27074
rect 53790 27010 53842 27022
rect 5630 26962 5682 26974
rect 5630 26898 5682 26910
rect 10334 26962 10386 26974
rect 13470 26962 13522 26974
rect 11890 26910 11902 26962
rect 11954 26910 11966 26962
rect 10334 26898 10386 26910
rect 13470 26898 13522 26910
rect 13806 26962 13858 26974
rect 41134 26962 41186 26974
rect 24210 26910 24222 26962
rect 24274 26910 24286 26962
rect 34514 26910 34526 26962
rect 34578 26910 34590 26962
rect 36194 26910 36206 26962
rect 36258 26910 36270 26962
rect 13806 26898 13858 26910
rect 41134 26898 41186 26910
rect 41694 26962 41746 26974
rect 41694 26898 41746 26910
rect 42702 26962 42754 26974
rect 42702 26898 42754 26910
rect 43038 26962 43090 26974
rect 51214 26962 51266 26974
rect 49746 26910 49758 26962
rect 49810 26910 49822 26962
rect 50418 26910 50430 26962
rect 50482 26910 50494 26962
rect 43038 26898 43090 26910
rect 51214 26898 51266 26910
rect 52110 26962 52162 26974
rect 52110 26898 52162 26910
rect 54462 26962 54514 26974
rect 54462 26898 54514 26910
rect 7086 26850 7138 26862
rect 7086 26786 7138 26798
rect 7646 26850 7698 26862
rect 7646 26786 7698 26798
rect 22654 26850 22706 26862
rect 22654 26786 22706 26798
rect 22878 26850 22930 26862
rect 22878 26786 22930 26798
rect 33182 26850 33234 26862
rect 33182 26786 33234 26798
rect 35646 26850 35698 26862
rect 35646 26786 35698 26798
rect 37214 26850 37266 26862
rect 37214 26786 37266 26798
rect 38670 26850 38722 26862
rect 38670 26786 38722 26798
rect 38894 26850 38946 26862
rect 38894 26786 38946 26798
rect 39342 26850 39394 26862
rect 39342 26786 39394 26798
rect 39454 26850 39506 26862
rect 39454 26786 39506 26798
rect 41246 26850 41298 26862
rect 41246 26786 41298 26798
rect 48526 26850 48578 26862
rect 48526 26786 48578 26798
rect 51102 26850 51154 26862
rect 51102 26786 51154 26798
rect 51998 26850 52050 26862
rect 51998 26786 52050 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 10110 26514 10162 26526
rect 10110 26450 10162 26462
rect 15710 26514 15762 26526
rect 15710 26450 15762 26462
rect 22766 26514 22818 26526
rect 22766 26450 22818 26462
rect 24222 26514 24274 26526
rect 36990 26514 37042 26526
rect 36082 26462 36094 26514
rect 36146 26462 36158 26514
rect 24222 26450 24274 26462
rect 36990 26450 37042 26462
rect 42702 26514 42754 26526
rect 42702 26450 42754 26462
rect 43598 26514 43650 26526
rect 43598 26450 43650 26462
rect 44046 26514 44098 26526
rect 48862 26514 48914 26526
rect 46722 26462 46734 26514
rect 46786 26462 46798 26514
rect 44046 26450 44098 26462
rect 48862 26450 48914 26462
rect 10558 26402 10610 26414
rect 21086 26402 21138 26414
rect 7522 26350 7534 26402
rect 7586 26350 7598 26402
rect 13122 26350 13134 26402
rect 13186 26350 13198 26402
rect 10558 26338 10610 26350
rect 21086 26338 21138 26350
rect 21870 26402 21922 26414
rect 22990 26402 23042 26414
rect 32398 26402 32450 26414
rect 22530 26350 22542 26402
rect 22594 26350 22606 26402
rect 29026 26350 29038 26402
rect 29090 26350 29102 26402
rect 29698 26350 29710 26402
rect 29762 26350 29774 26402
rect 21870 26338 21922 26350
rect 22990 26338 23042 26350
rect 32398 26338 32450 26350
rect 34526 26402 34578 26414
rect 47630 26402 47682 26414
rect 39330 26350 39342 26402
rect 39394 26350 39406 26402
rect 44482 26350 44494 26402
rect 44546 26350 44558 26402
rect 34526 26338 34578 26350
rect 47630 26338 47682 26350
rect 49422 26402 49474 26414
rect 53442 26350 53454 26402
rect 53506 26350 53518 26402
rect 53890 26350 53902 26402
rect 53954 26350 53966 26402
rect 49422 26338 49474 26350
rect 6974 26290 7026 26302
rect 10894 26290 10946 26302
rect 18958 26290 19010 26302
rect 7410 26238 7422 26290
rect 7474 26238 7486 26290
rect 12338 26238 12350 26290
rect 12402 26238 12414 26290
rect 6974 26226 7026 26238
rect 10894 26226 10946 26238
rect 18958 26226 19010 26238
rect 19518 26290 19570 26302
rect 20750 26290 20802 26302
rect 20402 26238 20414 26290
rect 20466 26238 20478 26290
rect 19518 26226 19570 26238
rect 20750 26226 20802 26238
rect 21198 26290 21250 26302
rect 21198 26226 21250 26238
rect 21422 26290 21474 26302
rect 21422 26226 21474 26238
rect 21646 26290 21698 26302
rect 23102 26290 23154 26302
rect 24334 26290 24386 26302
rect 22306 26238 22318 26290
rect 22370 26238 22382 26290
rect 23538 26238 23550 26290
rect 23602 26238 23614 26290
rect 24098 26238 24110 26290
rect 24162 26238 24174 26290
rect 21646 26226 21698 26238
rect 23102 26226 23154 26238
rect 24334 26226 24386 26238
rect 25118 26290 25170 26302
rect 25118 26226 25170 26238
rect 25454 26290 25506 26302
rect 25454 26226 25506 26238
rect 25678 26290 25730 26302
rect 25678 26226 25730 26238
rect 28702 26290 28754 26302
rect 31614 26290 31666 26302
rect 29474 26238 29486 26290
rect 29538 26238 29550 26290
rect 28702 26226 28754 26238
rect 31614 26226 31666 26238
rect 32062 26290 32114 26302
rect 32062 26226 32114 26238
rect 33070 26290 33122 26302
rect 33070 26226 33122 26238
rect 33294 26290 33346 26302
rect 33294 26226 33346 26238
rect 33518 26290 33570 26302
rect 33518 26226 33570 26238
rect 33630 26290 33682 26302
rect 33630 26226 33682 26238
rect 34078 26290 34130 26302
rect 34078 26226 34130 26238
rect 34414 26290 34466 26302
rect 34414 26226 34466 26238
rect 35310 26290 35362 26302
rect 35310 26226 35362 26238
rect 35534 26290 35586 26302
rect 35534 26226 35586 26238
rect 35982 26290 36034 26302
rect 36542 26290 36594 26302
rect 40910 26290 40962 26302
rect 36194 26238 36206 26290
rect 36258 26238 36270 26290
rect 40114 26238 40126 26290
rect 40178 26238 40190 26290
rect 35982 26226 36034 26238
rect 36542 26226 36594 26238
rect 40910 26226 40962 26238
rect 41246 26290 41298 26302
rect 41246 26226 41298 26238
rect 41470 26290 41522 26302
rect 41470 26226 41522 26238
rect 41918 26290 41970 26302
rect 49534 26290 49586 26302
rect 51550 26290 51602 26302
rect 54350 26290 54402 26302
rect 44370 26238 44382 26290
rect 44434 26238 44446 26290
rect 48178 26238 48190 26290
rect 48242 26238 48254 26290
rect 49858 26238 49870 26290
rect 49922 26238 49934 26290
rect 50978 26238 50990 26290
rect 51042 26238 51054 26290
rect 51314 26238 51326 26290
rect 51378 26238 51390 26290
rect 52322 26238 52334 26290
rect 52386 26238 52398 26290
rect 53330 26238 53342 26290
rect 53394 26238 53406 26290
rect 54786 26238 54798 26290
rect 54850 26238 54862 26290
rect 41918 26226 41970 26238
rect 49534 26226 49586 26238
rect 51550 26226 51602 26238
rect 54350 26226 54402 26238
rect 18622 26178 18674 26190
rect 15250 26126 15262 26178
rect 15314 26126 15326 26178
rect 18622 26114 18674 26126
rect 20862 26178 20914 26190
rect 20862 26114 20914 26126
rect 23886 26178 23938 26190
rect 23886 26114 23938 26126
rect 25342 26178 25394 26190
rect 25342 26114 25394 26126
rect 26686 26178 26738 26190
rect 26686 26114 26738 26126
rect 33182 26178 33234 26190
rect 33182 26114 33234 26126
rect 35758 26178 35810 26190
rect 41022 26178 41074 26190
rect 37202 26126 37214 26178
rect 37266 26126 37278 26178
rect 35758 26114 35810 26126
rect 41022 26114 41074 26126
rect 51438 26178 51490 26190
rect 52210 26126 52222 26178
rect 52274 26126 52286 26178
rect 51438 26114 51490 26126
rect 6638 26066 6690 26078
rect 26462 26066 26514 26078
rect 26114 26014 26126 26066
rect 26178 26014 26190 26066
rect 6638 26002 6690 26014
rect 26462 26002 26514 26014
rect 32510 26066 32562 26078
rect 32510 26002 32562 26014
rect 34526 26066 34578 26078
rect 50978 26014 50990 26066
rect 51042 26014 51054 26066
rect 52434 26014 52446 26066
rect 52498 26014 52510 26066
rect 34526 26002 34578 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 10670 25730 10722 25742
rect 10670 25666 10722 25678
rect 13582 25730 13634 25742
rect 13582 25666 13634 25678
rect 13918 25730 13970 25742
rect 53902 25730 53954 25742
rect 39554 25678 39566 25730
rect 39618 25678 39630 25730
rect 46498 25678 46510 25730
rect 46562 25678 46574 25730
rect 13918 25666 13970 25678
rect 53902 25666 53954 25678
rect 12798 25618 12850 25630
rect 46958 25618 47010 25630
rect 54014 25618 54066 25630
rect 9874 25566 9886 25618
rect 9938 25566 9950 25618
rect 18386 25566 18398 25618
rect 18450 25566 18462 25618
rect 25666 25566 25678 25618
rect 25730 25566 25742 25618
rect 27794 25566 27806 25618
rect 27858 25566 27870 25618
rect 30482 25566 30494 25618
rect 30546 25566 30558 25618
rect 32610 25566 32622 25618
rect 32674 25566 32686 25618
rect 33954 25566 33966 25618
rect 34018 25566 34030 25618
rect 40114 25566 40126 25618
rect 40178 25566 40190 25618
rect 41234 25566 41246 25618
rect 41298 25566 41310 25618
rect 45266 25566 45278 25618
rect 45330 25566 45342 25618
rect 47282 25566 47294 25618
rect 47346 25566 47358 25618
rect 50866 25566 50878 25618
rect 50930 25566 50942 25618
rect 52882 25566 52894 25618
rect 52946 25566 52958 25618
rect 12798 25554 12850 25566
rect 46958 25554 47010 25566
rect 54014 25554 54066 25566
rect 5966 25506 6018 25518
rect 12238 25506 12290 25518
rect 21646 25506 21698 25518
rect 23998 25506 24050 25518
rect 7074 25454 7086 25506
rect 7138 25454 7150 25506
rect 11442 25454 11454 25506
rect 11506 25454 11518 25506
rect 15586 25454 15598 25506
rect 15650 25454 15662 25506
rect 20290 25454 20302 25506
rect 20354 25454 20366 25506
rect 23538 25454 23550 25506
rect 23602 25454 23614 25506
rect 5966 25442 6018 25454
rect 12238 25442 12290 25454
rect 21646 25442 21698 25454
rect 23998 25442 24050 25454
rect 24334 25506 24386 25518
rect 24334 25442 24386 25454
rect 24894 25506 24946 25518
rect 40014 25506 40066 25518
rect 28578 25454 28590 25506
rect 28642 25454 28654 25506
rect 29698 25454 29710 25506
rect 29762 25454 29774 25506
rect 33058 25454 33070 25506
rect 33122 25454 33134 25506
rect 36194 25454 36206 25506
rect 36258 25454 36270 25506
rect 37090 25454 37102 25506
rect 37154 25454 37166 25506
rect 37986 25454 37998 25506
rect 38050 25454 38062 25506
rect 38210 25454 38222 25506
rect 38274 25454 38286 25506
rect 39890 25454 39902 25506
rect 39954 25454 39966 25506
rect 24894 25442 24946 25454
rect 40014 25442 40066 25454
rect 40798 25506 40850 25518
rect 45950 25506 46002 25518
rect 42242 25454 42254 25506
rect 42306 25454 42318 25506
rect 42802 25454 42814 25506
rect 42866 25454 42878 25506
rect 43138 25454 43150 25506
rect 43202 25454 43214 25506
rect 44930 25454 44942 25506
rect 44994 25454 45006 25506
rect 45714 25454 45726 25506
rect 45778 25454 45790 25506
rect 40798 25442 40850 25454
rect 45950 25442 46002 25454
rect 46062 25506 46114 25518
rect 47394 25454 47406 25506
rect 47458 25454 47470 25506
rect 47618 25454 47630 25506
rect 47682 25454 47694 25506
rect 49186 25454 49198 25506
rect 49250 25454 49262 25506
rect 50642 25454 50654 25506
rect 50706 25454 50718 25506
rect 52770 25454 52782 25506
rect 52834 25454 52846 25506
rect 46062 25442 46114 25454
rect 19294 25394 19346 25406
rect 7746 25342 7758 25394
rect 7810 25342 7822 25394
rect 11218 25342 11230 25394
rect 11282 25342 11294 25394
rect 11890 25342 11902 25394
rect 11954 25342 11966 25394
rect 14130 25342 14142 25394
rect 14194 25342 14206 25394
rect 14690 25342 14702 25394
rect 14754 25342 14766 25394
rect 16258 25342 16270 25394
rect 16322 25342 16334 25394
rect 19294 25330 19346 25342
rect 19854 25394 19906 25406
rect 19854 25330 19906 25342
rect 20750 25394 20802 25406
rect 20750 25330 20802 25342
rect 29374 25394 29426 25406
rect 44158 25394 44210 25406
rect 54462 25394 54514 25406
rect 33842 25342 33854 25394
rect 33906 25342 33918 25394
rect 34626 25342 34638 25394
rect 34690 25342 34702 25394
rect 37762 25342 37774 25394
rect 37826 25342 37838 25394
rect 42578 25342 42590 25394
rect 42642 25342 42654 25394
rect 53330 25342 53342 25394
rect 53394 25342 53406 25394
rect 29374 25330 29426 25342
rect 44158 25330 44210 25342
rect 54462 25330 54514 25342
rect 5630 25282 5682 25294
rect 5630 25218 5682 25230
rect 10334 25282 10386 25294
rect 10334 25218 10386 25230
rect 18734 25282 18786 25294
rect 22654 25282 22706 25294
rect 21970 25230 21982 25282
rect 22034 25230 22046 25282
rect 18734 25218 18786 25230
rect 22654 25218 22706 25230
rect 23102 25282 23154 25294
rect 23102 25218 23154 25230
rect 25342 25282 25394 25294
rect 25342 25218 25394 25230
rect 44270 25282 44322 25294
rect 44270 25218 44322 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 7758 24946 7810 24958
rect 7758 24882 7810 24894
rect 13022 24946 13074 24958
rect 20638 24946 20690 24958
rect 15474 24894 15486 24946
rect 15538 24894 15550 24946
rect 13022 24882 13074 24894
rect 20638 24882 20690 24894
rect 20750 24946 20802 24958
rect 20750 24882 20802 24894
rect 22318 24946 22370 24958
rect 22318 24882 22370 24894
rect 22766 24946 22818 24958
rect 22766 24882 22818 24894
rect 24670 24946 24722 24958
rect 24670 24882 24722 24894
rect 26350 24946 26402 24958
rect 26350 24882 26402 24894
rect 28478 24946 28530 24958
rect 28478 24882 28530 24894
rect 29374 24946 29426 24958
rect 29374 24882 29426 24894
rect 32510 24946 32562 24958
rect 32510 24882 32562 24894
rect 32622 24946 32674 24958
rect 32622 24882 32674 24894
rect 36990 24946 37042 24958
rect 41682 24894 41694 24946
rect 41746 24894 41758 24946
rect 49522 24894 49534 24946
rect 49586 24894 49598 24946
rect 36990 24882 37042 24894
rect 8094 24834 8146 24846
rect 4946 24782 4958 24834
rect 5010 24782 5022 24834
rect 8094 24770 8146 24782
rect 8878 24834 8930 24846
rect 18510 24834 18562 24846
rect 10434 24782 10446 24834
rect 10498 24782 10510 24834
rect 8878 24770 8930 24782
rect 18510 24770 18562 24782
rect 20862 24834 20914 24846
rect 23550 24834 23602 24846
rect 23090 24782 23102 24834
rect 23154 24782 23166 24834
rect 20862 24770 20914 24782
rect 23550 24770 23602 24782
rect 23662 24834 23714 24846
rect 32062 24834 32114 24846
rect 35422 24834 35474 24846
rect 26674 24782 26686 24834
rect 26738 24782 26750 24834
rect 28130 24782 28142 24834
rect 28194 24782 28206 24834
rect 33058 24782 33070 24834
rect 33122 24782 33134 24834
rect 23662 24770 23714 24782
rect 32062 24770 32114 24782
rect 35422 24770 35474 24782
rect 35646 24834 35698 24846
rect 35646 24770 35698 24782
rect 37438 24834 37490 24846
rect 37438 24770 37490 24782
rect 38894 24834 38946 24846
rect 47182 24834 47234 24846
rect 42690 24782 42702 24834
rect 42754 24782 42766 24834
rect 38894 24770 38946 24782
rect 47182 24770 47234 24782
rect 47518 24834 47570 24846
rect 47518 24770 47570 24782
rect 48974 24834 49026 24846
rect 51090 24782 51102 24834
rect 51154 24782 51166 24834
rect 52658 24782 52670 24834
rect 52722 24782 52734 24834
rect 48974 24770 49026 24782
rect 15822 24722 15874 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 9650 24670 9662 24722
rect 9714 24670 9726 24722
rect 15822 24658 15874 24670
rect 16270 24722 16322 24734
rect 19630 24722 19682 24734
rect 25566 24722 25618 24734
rect 41022 24722 41074 24734
rect 18162 24670 18174 24722
rect 18226 24670 18238 24722
rect 19058 24670 19070 24722
rect 19122 24670 19134 24722
rect 21634 24670 21646 24722
rect 21698 24670 21710 24722
rect 32274 24670 32286 24722
rect 32338 24670 32350 24722
rect 33842 24670 33854 24722
rect 33906 24670 33918 24722
rect 34066 24670 34078 24722
rect 34130 24670 34142 24722
rect 36194 24670 36206 24722
rect 36258 24670 36270 24722
rect 40002 24670 40014 24722
rect 40066 24670 40078 24722
rect 16270 24658 16322 24670
rect 19630 24658 19682 24670
rect 25566 24658 25618 24670
rect 41022 24658 41074 24670
rect 41134 24722 41186 24734
rect 41134 24658 41186 24670
rect 41246 24722 41298 24734
rect 47854 24722 47906 24734
rect 43474 24670 43486 24722
rect 43538 24670 43550 24722
rect 43922 24670 43934 24722
rect 43986 24670 43998 24722
rect 45378 24670 45390 24722
rect 45442 24670 45454 24722
rect 46498 24670 46510 24722
rect 46562 24670 46574 24722
rect 41246 24658 41298 24670
rect 47854 24658 47906 24670
rect 48190 24722 48242 24734
rect 48190 24658 48242 24670
rect 49198 24722 49250 24734
rect 49198 24658 49250 24670
rect 49534 24722 49586 24734
rect 49858 24670 49870 24722
rect 49922 24670 49934 24722
rect 51314 24670 51326 24722
rect 51378 24670 51390 24722
rect 51986 24670 51998 24722
rect 52050 24670 52062 24722
rect 49534 24658 49586 24670
rect 25230 24610 25282 24622
rect 47966 24610 48018 24622
rect 7074 24558 7086 24610
rect 7138 24558 7150 24610
rect 12562 24558 12574 24610
rect 12626 24558 12638 24610
rect 17826 24558 17838 24610
rect 17890 24558 17902 24610
rect 19170 24558 19182 24610
rect 19234 24558 19246 24610
rect 20066 24558 20078 24610
rect 20130 24558 20142 24610
rect 21298 24558 21310 24610
rect 21362 24558 21374 24610
rect 24210 24558 24222 24610
rect 24274 24558 24286 24610
rect 25778 24558 25790 24610
rect 25842 24558 25854 24610
rect 28914 24558 28926 24610
rect 28978 24558 28990 24610
rect 42466 24558 42478 24610
rect 42530 24558 42542 24610
rect 46722 24558 46734 24610
rect 46786 24558 46798 24610
rect 25230 24546 25282 24558
rect 47966 24546 48018 24558
rect 50206 24610 50258 24622
rect 54786 24558 54798 24610
rect 54850 24558 54862 24610
rect 50206 24546 50258 24558
rect 8990 24498 9042 24510
rect 8990 24434 9042 24446
rect 22094 24498 22146 24510
rect 22094 24434 22146 24446
rect 22430 24498 22482 24510
rect 22430 24434 22482 24446
rect 23662 24498 23714 24510
rect 23662 24434 23714 24446
rect 35758 24498 35810 24510
rect 35758 24434 35810 24446
rect 49422 24498 49474 24510
rect 49422 24434 49474 24446
rect 50430 24498 50482 24510
rect 50430 24434 50482 24446
rect 50766 24498 50818 24510
rect 50766 24434 50818 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 11230 24162 11282 24174
rect 11230 24098 11282 24110
rect 11566 24162 11618 24174
rect 11566 24098 11618 24110
rect 14926 24162 14978 24174
rect 14926 24098 14978 24110
rect 35422 24162 35474 24174
rect 35422 24098 35474 24110
rect 43934 24162 43986 24174
rect 49198 24162 49250 24174
rect 47170 24110 47182 24162
rect 47234 24110 47246 24162
rect 43934 24098 43986 24110
rect 49198 24098 49250 24110
rect 7422 24050 7474 24062
rect 8654 24050 8706 24062
rect 8306 23998 8318 24050
rect 8370 23998 8382 24050
rect 7422 23986 7474 23998
rect 8654 23986 8706 23998
rect 9214 24050 9266 24062
rect 32510 24050 32562 24062
rect 23538 23998 23550 24050
rect 23602 23998 23614 24050
rect 29138 23998 29150 24050
rect 29202 23998 29214 24050
rect 9214 23986 9266 23998
rect 32510 23986 32562 23998
rect 33630 24050 33682 24062
rect 33630 23986 33682 23998
rect 34078 24050 34130 24062
rect 34078 23986 34130 23998
rect 34190 24050 34242 24062
rect 34190 23986 34242 23998
rect 36318 24050 36370 24062
rect 43710 24050 43762 24062
rect 37314 23998 37326 24050
rect 37378 23998 37390 24050
rect 36318 23986 36370 23998
rect 43710 23986 43762 23998
rect 53230 24050 53282 24062
rect 53230 23986 53282 23998
rect 53678 24050 53730 24062
rect 53678 23986 53730 23998
rect 17278 23938 17330 23950
rect 7970 23886 7982 23938
rect 8034 23886 8046 23938
rect 12114 23886 12126 23938
rect 12178 23886 12190 23938
rect 17278 23874 17330 23886
rect 17502 23938 17554 23950
rect 17502 23874 17554 23886
rect 19630 23938 19682 23950
rect 19630 23874 19682 23886
rect 19966 23938 20018 23950
rect 23102 23938 23154 23950
rect 33182 23938 33234 23950
rect 35646 23938 35698 23950
rect 38334 23938 38386 23950
rect 44942 23938 44994 23950
rect 21970 23886 21982 23938
rect 22034 23886 22046 23938
rect 22530 23886 22542 23938
rect 22594 23886 22606 23938
rect 24882 23886 24894 23938
rect 24946 23886 24958 23938
rect 25554 23886 25566 23938
rect 25618 23886 25630 23938
rect 32050 23886 32062 23938
rect 32114 23886 32126 23938
rect 35186 23886 35198 23938
rect 35250 23886 35262 23938
rect 37202 23886 37214 23938
rect 37266 23886 37278 23938
rect 37874 23886 37886 23938
rect 37938 23886 37950 23938
rect 40002 23886 40014 23938
rect 40066 23886 40078 23938
rect 41682 23886 41694 23938
rect 41746 23886 41758 23938
rect 42018 23886 42030 23938
rect 42082 23886 42094 23938
rect 19966 23874 20018 23886
rect 23102 23874 23154 23886
rect 33182 23874 33234 23886
rect 35646 23874 35698 23886
rect 38334 23874 38386 23886
rect 44942 23874 44994 23886
rect 45166 23938 45218 23950
rect 45166 23874 45218 23886
rect 45390 23938 45442 23950
rect 45950 23938 46002 23950
rect 45602 23886 45614 23938
rect 45666 23886 45678 23938
rect 45390 23874 45442 23886
rect 45950 23874 46002 23886
rect 46174 23938 46226 23950
rect 46174 23874 46226 23886
rect 46734 23938 46786 23950
rect 50878 23938 50930 23950
rect 47954 23886 47966 23938
rect 48018 23886 48030 23938
rect 50418 23886 50430 23938
rect 50482 23886 50494 23938
rect 46734 23874 46786 23886
rect 50878 23874 50930 23886
rect 51214 23938 51266 23950
rect 51214 23874 51266 23886
rect 51438 23938 51490 23950
rect 51438 23874 51490 23886
rect 4622 23826 4674 23838
rect 17614 23826 17666 23838
rect 7746 23774 7758 23826
rect 7810 23774 7822 23826
rect 12226 23774 12238 23826
rect 12290 23774 12302 23826
rect 15138 23774 15150 23826
rect 15202 23774 15214 23826
rect 15474 23774 15486 23826
rect 15538 23774 15550 23826
rect 4622 23762 4674 23774
rect 17614 23762 17666 23774
rect 17838 23826 17890 23838
rect 17838 23762 17890 23774
rect 18734 23826 18786 23838
rect 18734 23762 18786 23774
rect 21534 23826 21586 23838
rect 33406 23826 33458 23838
rect 23986 23774 23998 23826
rect 24050 23774 24062 23826
rect 31266 23774 31278 23826
rect 31330 23774 31342 23826
rect 21534 23762 21586 23774
rect 33406 23762 33458 23774
rect 33742 23826 33794 23838
rect 33742 23762 33794 23774
rect 34302 23826 34354 23838
rect 34302 23762 34354 23774
rect 34974 23826 35026 23838
rect 34974 23762 35026 23774
rect 35870 23826 35922 23838
rect 46510 23826 46562 23838
rect 37426 23774 37438 23826
rect 37490 23774 37502 23826
rect 39890 23774 39902 23826
rect 39954 23774 39966 23826
rect 41122 23774 41134 23826
rect 41186 23774 41198 23826
rect 42130 23774 42142 23826
rect 42194 23774 42206 23826
rect 42578 23774 42590 23826
rect 42642 23774 42654 23826
rect 35870 23762 35922 23774
rect 46510 23762 46562 23774
rect 47630 23826 47682 23838
rect 47630 23762 47682 23774
rect 47742 23826 47794 23838
rect 47742 23762 47794 23774
rect 48750 23826 48802 23838
rect 48750 23762 48802 23774
rect 49422 23826 49474 23838
rect 49422 23762 49474 23774
rect 50990 23826 51042 23838
rect 50990 23762 51042 23774
rect 51662 23826 51714 23838
rect 51662 23762 51714 23774
rect 51886 23826 51938 23838
rect 51886 23762 51938 23774
rect 52782 23826 52834 23838
rect 52782 23762 52834 23774
rect 4286 23714 4338 23726
rect 4286 23650 4338 23662
rect 6414 23714 6466 23726
rect 6414 23650 6466 23662
rect 8766 23714 8818 23726
rect 8766 23650 8818 23662
rect 13806 23714 13858 23726
rect 13806 23650 13858 23662
rect 14254 23714 14306 23726
rect 14254 23650 14306 23662
rect 14590 23714 14642 23726
rect 18286 23714 18338 23726
rect 16818 23662 16830 23714
rect 16882 23662 16894 23714
rect 14590 23650 14642 23662
rect 18286 23650 18338 23662
rect 22878 23714 22930 23726
rect 22878 23650 22930 23662
rect 22990 23714 23042 23726
rect 22990 23650 23042 23662
rect 35982 23714 36034 23726
rect 46398 23714 46450 23726
rect 43026 23662 43038 23714
rect 43090 23662 43102 23714
rect 44258 23662 44270 23714
rect 44322 23662 44334 23714
rect 45490 23662 45502 23714
rect 45554 23662 45566 23714
rect 35982 23650 36034 23662
rect 46398 23650 46450 23662
rect 48302 23714 48354 23726
rect 48302 23650 48354 23662
rect 48414 23714 48466 23726
rect 48414 23650 48466 23662
rect 48526 23714 48578 23726
rect 48526 23650 48578 23662
rect 49310 23714 49362 23726
rect 49310 23650 49362 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 6526 23378 6578 23390
rect 17726 23378 17778 23390
rect 12898 23326 12910 23378
rect 12962 23326 12974 23378
rect 6526 23314 6578 23326
rect 17726 23314 17778 23326
rect 17950 23378 18002 23390
rect 17950 23314 18002 23326
rect 24446 23378 24498 23390
rect 24446 23314 24498 23326
rect 29374 23378 29426 23390
rect 29374 23314 29426 23326
rect 33966 23378 34018 23390
rect 33966 23314 34018 23326
rect 34302 23378 34354 23390
rect 34302 23314 34354 23326
rect 34526 23378 34578 23390
rect 41806 23378 41858 23390
rect 38546 23326 38558 23378
rect 38610 23326 38622 23378
rect 34526 23314 34578 23326
rect 41806 23314 41858 23326
rect 49198 23378 49250 23390
rect 51886 23378 51938 23390
rect 50866 23326 50878 23378
rect 50930 23326 50942 23378
rect 49198 23314 49250 23326
rect 51886 23314 51938 23326
rect 52334 23378 52386 23390
rect 52334 23314 52386 23326
rect 2382 23266 2434 23278
rect 24334 23266 24386 23278
rect 3938 23214 3950 23266
rect 4002 23214 4014 23266
rect 7410 23214 7422 23266
rect 7474 23214 7486 23266
rect 20066 23214 20078 23266
rect 20130 23214 20142 23266
rect 22194 23214 22206 23266
rect 22258 23214 22270 23266
rect 23090 23214 23102 23266
rect 23154 23214 23166 23266
rect 2382 23202 2434 23214
rect 24334 23202 24386 23214
rect 34190 23266 34242 23278
rect 39678 23266 39730 23278
rect 34738 23214 34750 23266
rect 34802 23214 34814 23266
rect 36418 23214 36430 23266
rect 36482 23214 36494 23266
rect 38770 23214 38782 23266
rect 38834 23214 38846 23266
rect 34190 23202 34242 23214
rect 39678 23202 39730 23214
rect 39790 23266 39842 23278
rect 46062 23266 46114 23278
rect 42578 23214 42590 23266
rect 42642 23214 42654 23266
rect 39790 23202 39842 23214
rect 46062 23202 46114 23214
rect 46510 23266 46562 23278
rect 49646 23266 49698 23278
rect 52446 23266 52498 23278
rect 47506 23214 47518 23266
rect 47570 23214 47582 23266
rect 50754 23214 50766 23266
rect 50818 23214 50830 23266
rect 46510 23202 46562 23214
rect 49646 23202 49698 23214
rect 52446 23202 52498 23214
rect 53006 23266 53058 23278
rect 53006 23202 53058 23214
rect 2718 23154 2770 23166
rect 9662 23154 9714 23166
rect 3266 23102 3278 23154
rect 3330 23102 3342 23154
rect 7634 23102 7646 23154
rect 7698 23102 7710 23154
rect 2718 23090 2770 23102
rect 9662 23090 9714 23102
rect 13246 23154 13298 23166
rect 18062 23154 18114 23166
rect 13794 23102 13806 23154
rect 13858 23102 13870 23154
rect 13246 23090 13298 23102
rect 18062 23090 18114 23102
rect 18622 23154 18674 23166
rect 24670 23154 24722 23166
rect 35086 23154 35138 23166
rect 39454 23154 39506 23166
rect 20738 23102 20750 23154
rect 20802 23102 20814 23154
rect 22642 23102 22654 23154
rect 22706 23102 22718 23154
rect 28578 23102 28590 23154
rect 28642 23102 28654 23154
rect 29138 23102 29150 23154
rect 29202 23102 29214 23154
rect 35634 23102 35646 23154
rect 35698 23102 35710 23154
rect 36530 23102 36542 23154
rect 36594 23102 36606 23154
rect 37762 23102 37774 23154
rect 37826 23102 37838 23154
rect 38994 23102 39006 23154
rect 39058 23102 39070 23154
rect 18622 23090 18674 23102
rect 24670 23090 24722 23102
rect 35086 23090 35138 23102
rect 39454 23090 39506 23102
rect 40238 23154 40290 23166
rect 46286 23154 46338 23166
rect 48638 23154 48690 23166
rect 43586 23102 43598 23154
rect 43650 23102 43662 23154
rect 43810 23102 43822 23154
rect 43874 23102 43886 23154
rect 45378 23102 45390 23154
rect 45442 23102 45454 23154
rect 47058 23102 47070 23154
rect 47122 23102 47134 23154
rect 47954 23102 47966 23154
rect 48018 23102 48030 23154
rect 40238 23090 40290 23102
rect 46286 23090 46338 23102
rect 48638 23090 48690 23102
rect 49086 23154 49138 23166
rect 49086 23090 49138 23102
rect 49310 23154 49362 23166
rect 49310 23090 49362 23102
rect 50094 23154 50146 23166
rect 50094 23090 50146 23102
rect 50542 23154 50594 23166
rect 51314 23102 51326 23154
rect 51378 23102 51390 23154
rect 50542 23090 50594 23102
rect 12574 23042 12626 23054
rect 6066 22990 6078 23042
rect 6130 22990 6142 23042
rect 12574 22978 12626 22990
rect 13470 23042 13522 23054
rect 25342 23042 25394 23054
rect 46174 23042 46226 23054
rect 49758 23042 49810 23054
rect 14578 22990 14590 23042
rect 14642 22990 14654 23042
rect 16706 22990 16718 23042
rect 16770 22990 16782 23042
rect 19842 22990 19854 23042
rect 19906 22990 19918 23042
rect 23426 22990 23438 23042
rect 23490 22990 23502 23042
rect 25666 22990 25678 23042
rect 25730 22990 25742 23042
rect 27794 22990 27806 23042
rect 27858 22990 27870 23042
rect 42130 22990 42142 23042
rect 42194 22990 42206 23042
rect 47394 22990 47406 23042
rect 47458 22990 47470 23042
rect 13470 22978 13522 22990
rect 25342 22978 25394 22990
rect 46174 22978 46226 22990
rect 49758 22978 49810 22990
rect 49982 23042 50034 23054
rect 49982 22978 50034 22990
rect 51774 23042 51826 23054
rect 51774 22978 51826 22990
rect 6862 22930 6914 22942
rect 6862 22866 6914 22878
rect 18510 22930 18562 22942
rect 40462 22930 40514 22942
rect 51662 22930 51714 22942
rect 19618 22878 19630 22930
rect 19682 22878 19694 22930
rect 51090 22878 51102 22930
rect 51154 22878 51166 22930
rect 18510 22866 18562 22878
rect 40462 22866 40514 22878
rect 51662 22866 51714 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 5742 22594 5794 22606
rect 5742 22530 5794 22542
rect 8654 22594 8706 22606
rect 8654 22530 8706 22542
rect 13582 22594 13634 22606
rect 13582 22530 13634 22542
rect 15150 22594 15202 22606
rect 15150 22530 15202 22542
rect 25790 22594 25842 22606
rect 25790 22530 25842 22542
rect 29262 22594 29314 22606
rect 29262 22530 29314 22542
rect 29598 22594 29650 22606
rect 29598 22530 29650 22542
rect 36094 22594 36146 22606
rect 36094 22530 36146 22542
rect 38222 22594 38274 22606
rect 38222 22530 38274 22542
rect 38334 22594 38386 22606
rect 38334 22530 38386 22542
rect 38558 22594 38610 22606
rect 38558 22530 38610 22542
rect 38670 22594 38722 22606
rect 48750 22594 48802 22606
rect 40898 22542 40910 22594
rect 40962 22542 40974 22594
rect 44818 22542 44830 22594
rect 44882 22542 44894 22594
rect 50978 22542 50990 22594
rect 51042 22591 51054 22594
rect 51650 22591 51662 22594
rect 51042 22545 51662 22591
rect 51042 22542 51054 22545
rect 51650 22542 51662 22545
rect 51714 22542 51726 22594
rect 38670 22530 38722 22542
rect 48750 22530 48802 22542
rect 23102 22482 23154 22494
rect 2482 22430 2494 22482
rect 2546 22430 2558 22482
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 12562 22430 12574 22482
rect 12626 22430 12638 22482
rect 19170 22430 19182 22482
rect 19234 22430 19246 22482
rect 23102 22418 23154 22430
rect 24446 22482 24498 22494
rect 36206 22482 36258 22494
rect 37326 22482 37378 22494
rect 24882 22430 24894 22482
rect 24946 22430 24958 22482
rect 34178 22430 34190 22482
rect 34242 22430 34254 22482
rect 37090 22430 37102 22482
rect 37154 22430 37166 22482
rect 24446 22418 24498 22430
rect 36206 22418 36258 22430
rect 37326 22418 37378 22430
rect 39118 22482 39170 22494
rect 46510 22482 46562 22494
rect 40114 22430 40126 22482
rect 40178 22430 40190 22482
rect 40562 22430 40574 22482
rect 40626 22430 40638 22482
rect 42018 22430 42030 22482
rect 42082 22430 42094 22482
rect 39118 22418 39170 22430
rect 46510 22418 46562 22430
rect 48078 22482 48130 22494
rect 48078 22418 48130 22430
rect 49870 22482 49922 22494
rect 49870 22418 49922 22430
rect 51214 22482 51266 22494
rect 51214 22418 51266 22430
rect 52110 22482 52162 22494
rect 52110 22418 52162 22430
rect 6078 22370 6130 22382
rect 7646 22370 7698 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 6850 22318 6862 22370
rect 6914 22318 6926 22370
rect 6078 22306 6130 22318
rect 7646 22306 7698 22318
rect 7982 22370 8034 22382
rect 20638 22370 20690 22382
rect 8978 22318 8990 22370
rect 9042 22318 9054 22370
rect 9650 22318 9662 22370
rect 9714 22318 9726 22370
rect 14130 22318 14142 22370
rect 14194 22318 14206 22370
rect 18722 22318 18734 22370
rect 18786 22318 18798 22370
rect 7982 22306 8034 22318
rect 20638 22306 20690 22318
rect 22766 22370 22818 22382
rect 22766 22306 22818 22318
rect 24782 22370 24834 22382
rect 24782 22306 24834 22318
rect 25566 22370 25618 22382
rect 25566 22306 25618 22318
rect 27694 22370 27746 22382
rect 50766 22370 50818 22382
rect 28466 22318 28478 22370
rect 28530 22318 28542 22370
rect 33282 22318 33294 22370
rect 33346 22318 33358 22370
rect 36418 22318 36430 22370
rect 36482 22318 36494 22370
rect 39778 22318 39790 22370
rect 39842 22318 39854 22370
rect 40674 22318 40686 22370
rect 40738 22318 40750 22370
rect 42578 22318 42590 22370
rect 42642 22318 42654 22370
rect 42802 22318 42814 22370
rect 42866 22318 42878 22370
rect 46050 22318 46062 22370
rect 46114 22318 46126 22370
rect 47506 22318 47518 22370
rect 47570 22318 47582 22370
rect 47842 22318 47854 22370
rect 47906 22318 47918 22370
rect 48402 22318 48414 22370
rect 48466 22318 48478 22370
rect 27694 22306 27746 22318
rect 50766 22306 50818 22318
rect 51662 22370 51714 22382
rect 51662 22306 51714 22318
rect 13582 22258 13634 22270
rect 6738 22206 6750 22258
rect 6802 22206 6814 22258
rect 10434 22206 10446 22258
rect 10498 22206 10510 22258
rect 14366 22258 14418 22270
rect 21870 22258 21922 22270
rect 13582 22194 13634 22206
rect 13694 22202 13746 22214
rect 5070 22146 5122 22158
rect 5070 22082 5122 22094
rect 7534 22146 7586 22158
rect 7534 22082 7586 22094
rect 7870 22146 7922 22158
rect 7870 22082 7922 22094
rect 8766 22146 8818 22158
rect 15362 22206 15374 22258
rect 15426 22206 15438 22258
rect 15922 22206 15934 22258
rect 15986 22206 15998 22258
rect 18162 22206 18174 22258
rect 18226 22206 18238 22258
rect 19058 22206 19070 22258
rect 19122 22206 19134 22258
rect 14366 22194 14418 22206
rect 21870 22194 21922 22206
rect 26686 22258 26738 22270
rect 26686 22194 26738 22206
rect 26798 22258 26850 22270
rect 26798 22194 26850 22206
rect 27022 22258 27074 22270
rect 45278 22258 45330 22270
rect 28242 22206 28254 22258
rect 28306 22206 28318 22258
rect 29810 22206 29822 22258
rect 29874 22206 29886 22258
rect 30370 22206 30382 22258
rect 30434 22206 30446 22258
rect 43362 22206 43374 22258
rect 43426 22206 43438 22258
rect 27022 22194 27074 22206
rect 45278 22194 45330 22206
rect 45390 22258 45442 22270
rect 45390 22194 45442 22206
rect 45502 22258 45554 22270
rect 49758 22258 49810 22270
rect 49410 22206 49422 22258
rect 49474 22206 49486 22258
rect 45502 22194 45554 22206
rect 49758 22194 49810 22206
rect 49982 22258 50034 22270
rect 50418 22206 50430 22258
rect 50482 22206 50494 22258
rect 49982 22194 50034 22206
rect 13694 22138 13746 22150
rect 14814 22146 14866 22158
rect 26126 22146 26178 22158
rect 8766 22082 8818 22094
rect 23314 22094 23326 22146
rect 23378 22094 23390 22146
rect 14814 22082 14866 22094
rect 26126 22082 26178 22094
rect 27358 22146 27410 22158
rect 27358 22082 27410 22094
rect 37774 22146 37826 22158
rect 37774 22082 37826 22094
rect 48638 22146 48690 22158
rect 48638 22082 48690 22094
rect 49086 22146 49138 22158
rect 49086 22082 49138 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 8990 21810 9042 21822
rect 8990 21746 9042 21758
rect 10894 21810 10946 21822
rect 10894 21746 10946 21758
rect 27134 21810 27186 21822
rect 27134 21746 27186 21758
rect 29710 21810 29762 21822
rect 29710 21746 29762 21758
rect 30494 21810 30546 21822
rect 30494 21746 30546 21758
rect 35534 21810 35586 21822
rect 47630 21810 47682 21822
rect 49534 21810 49586 21822
rect 38882 21758 38894 21810
rect 38946 21758 38958 21810
rect 48738 21758 48750 21810
rect 48802 21758 48814 21810
rect 35534 21746 35586 21758
rect 47630 21746 47682 21758
rect 49534 21746 49586 21758
rect 7534 21698 7586 21710
rect 7534 21634 7586 21646
rect 7758 21698 7810 21710
rect 7758 21634 7810 21646
rect 8206 21698 8258 21710
rect 8206 21634 8258 21646
rect 9550 21698 9602 21710
rect 9550 21634 9602 21646
rect 11230 21698 11282 21710
rect 11230 21634 11282 21646
rect 11902 21698 11954 21710
rect 19854 21698 19906 21710
rect 12786 21646 12798 21698
rect 12850 21646 12862 21698
rect 14466 21646 14478 21698
rect 14530 21646 14542 21698
rect 11902 21634 11954 21646
rect 19854 21634 19906 21646
rect 19966 21698 20018 21710
rect 19966 21634 20018 21646
rect 21982 21698 22034 21710
rect 25230 21698 25282 21710
rect 23202 21646 23214 21698
rect 23266 21646 23278 21698
rect 23986 21646 23998 21698
rect 24050 21646 24062 21698
rect 24658 21646 24670 21698
rect 24722 21646 24734 21698
rect 21982 21634 22034 21646
rect 25230 21634 25282 21646
rect 26462 21698 26514 21710
rect 26462 21634 26514 21646
rect 29150 21698 29202 21710
rect 31950 21698 32002 21710
rect 34750 21698 34802 21710
rect 47406 21698 47458 21710
rect 30034 21646 30046 21698
rect 30098 21646 30110 21698
rect 33730 21646 33742 21698
rect 33794 21646 33806 21698
rect 34066 21646 34078 21698
rect 34130 21646 34142 21698
rect 36642 21646 36654 21698
rect 36706 21646 36718 21698
rect 41010 21646 41022 21698
rect 41074 21646 41086 21698
rect 46050 21646 46062 21698
rect 46114 21646 46126 21698
rect 50978 21646 50990 21698
rect 51042 21646 51054 21698
rect 29150 21634 29202 21646
rect 31950 21634 32002 21646
rect 34750 21634 34802 21646
rect 47406 21634 47458 21646
rect 8542 21586 8594 21598
rect 9998 21586 10050 21598
rect 12238 21586 12290 21598
rect 13918 21586 13970 21598
rect 16158 21586 16210 21598
rect 1810 21534 1822 21586
rect 1874 21534 1886 21586
rect 8866 21534 8878 21586
rect 8930 21534 8942 21586
rect 9762 21534 9774 21586
rect 9826 21534 9838 21586
rect 10098 21534 10110 21586
rect 10162 21534 10174 21586
rect 12898 21534 12910 21586
rect 12962 21534 12974 21586
rect 14690 21534 14702 21586
rect 14754 21534 14766 21586
rect 8542 21522 8594 21534
rect 9998 21522 10050 21534
rect 12238 21522 12290 21534
rect 13918 21522 13970 21534
rect 16158 21522 16210 21534
rect 16718 21586 16770 21598
rect 16718 21522 16770 21534
rect 20190 21586 20242 21598
rect 20190 21522 20242 21534
rect 20526 21586 20578 21598
rect 20526 21522 20578 21534
rect 20862 21586 20914 21598
rect 20862 21522 20914 21534
rect 22206 21586 22258 21598
rect 23550 21586 23602 21598
rect 25454 21586 25506 21598
rect 32286 21586 32338 21598
rect 22978 21534 22990 21586
rect 23042 21534 23054 21586
rect 24546 21534 24558 21586
rect 24610 21534 24622 21586
rect 26898 21534 26910 21586
rect 26962 21534 26974 21586
rect 22206 21522 22258 21534
rect 23550 21522 23602 21534
rect 25454 21522 25506 21534
rect 32286 21522 32338 21534
rect 33182 21586 33234 21598
rect 33182 21522 33234 21534
rect 35086 21586 35138 21598
rect 39902 21586 39954 21598
rect 35858 21534 35870 21586
rect 35922 21534 35934 21586
rect 35086 21522 35138 21534
rect 39902 21522 39954 21534
rect 40126 21586 40178 21598
rect 40126 21522 40178 21534
rect 40462 21586 40514 21598
rect 43038 21586 43090 21598
rect 47294 21586 47346 21598
rect 42018 21534 42030 21586
rect 42082 21534 42094 21586
rect 46834 21534 46846 21586
rect 46898 21534 46910 21586
rect 40462 21522 40514 21534
rect 43038 21522 43090 21534
rect 47294 21522 47346 21534
rect 47854 21586 47906 21598
rect 49646 21586 49698 21598
rect 48962 21534 48974 21586
rect 49026 21534 49038 21586
rect 50194 21534 50206 21586
rect 50258 21534 50270 21586
rect 47854 21522 47906 21534
rect 49646 21522 49698 21534
rect 5070 21474 5122 21486
rect 8654 21474 8706 21486
rect 2482 21422 2494 21474
rect 2546 21422 2558 21474
rect 4610 21422 4622 21474
rect 4674 21422 4686 21474
rect 7858 21422 7870 21474
rect 7922 21422 7934 21474
rect 5070 21410 5122 21422
rect 8654 21410 8706 21422
rect 9662 21474 9714 21486
rect 9662 21410 9714 21422
rect 15262 21474 15314 21486
rect 15262 21410 15314 21422
rect 17502 21474 17554 21486
rect 17502 21410 17554 21422
rect 18510 21474 18562 21486
rect 18510 21410 18562 21422
rect 26350 21474 26402 21486
rect 26350 21410 26402 21422
rect 40238 21474 40290 21486
rect 48302 21474 48354 21486
rect 42130 21422 42142 21474
rect 42194 21422 42206 21474
rect 43474 21422 43486 21474
rect 43538 21422 43550 21474
rect 43922 21422 43934 21474
rect 43986 21422 43998 21474
rect 53106 21422 53118 21474
rect 53170 21422 53182 21474
rect 40238 21410 40290 21422
rect 48302 21410 48354 21422
rect 13582 21362 13634 21374
rect 13582 21298 13634 21310
rect 20638 21362 20690 21374
rect 20638 21298 20690 21310
rect 21310 21362 21362 21374
rect 21310 21298 21362 21310
rect 22542 21362 22594 21374
rect 22542 21298 22594 21310
rect 23662 21362 23714 21374
rect 23662 21298 23714 21310
rect 25790 21362 25842 21374
rect 25790 21298 25842 21310
rect 29038 21362 29090 21374
rect 29038 21298 29090 21310
rect 33518 21362 33570 21374
rect 33518 21298 33570 21310
rect 49534 21362 49586 21374
rect 49534 21298 49586 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 4174 21026 4226 21038
rect 4174 20962 4226 20974
rect 7646 21026 7698 21038
rect 7646 20962 7698 20974
rect 7982 21026 8034 21038
rect 11790 21026 11842 21038
rect 18958 21026 19010 21038
rect 8530 20974 8542 21026
rect 8594 20974 8606 21026
rect 12338 20974 12350 21026
rect 12402 20974 12414 21026
rect 14354 20974 14366 21026
rect 14418 20974 14430 21026
rect 7982 20962 8034 20974
rect 11790 20962 11842 20974
rect 18958 20962 19010 20974
rect 20526 21026 20578 21038
rect 20526 20962 20578 20974
rect 21646 21026 21698 21038
rect 21646 20962 21698 20974
rect 23326 21026 23378 21038
rect 23326 20962 23378 20974
rect 35086 21026 35138 21038
rect 41794 20974 41806 21026
rect 41858 20974 41870 21026
rect 35086 20962 35138 20974
rect 11230 20914 11282 20926
rect 11230 20850 11282 20862
rect 20414 20914 20466 20926
rect 20414 20850 20466 20862
rect 24222 20914 24274 20926
rect 26350 20914 26402 20926
rect 24994 20862 25006 20914
rect 25058 20862 25070 20914
rect 24222 20850 24274 20862
rect 26350 20850 26402 20862
rect 27470 20914 27522 20926
rect 27470 20850 27522 20862
rect 28590 20914 28642 20926
rect 37214 20914 37266 20926
rect 42814 20914 42866 20926
rect 44270 20914 44322 20926
rect 48302 20914 48354 20926
rect 31826 20862 31838 20914
rect 31890 20862 31902 20914
rect 33954 20862 33966 20914
rect 34018 20862 34030 20914
rect 41234 20862 41246 20914
rect 41298 20862 41310 20914
rect 44034 20862 44046 20914
rect 44098 20862 44110 20914
rect 45602 20862 45614 20914
rect 45666 20862 45678 20914
rect 47730 20862 47742 20914
rect 47794 20862 47806 20914
rect 28590 20850 28642 20862
rect 37214 20850 37266 20862
rect 42814 20850 42866 20862
rect 44270 20850 44322 20862
rect 48302 20850 48354 20862
rect 48638 20914 48690 20926
rect 48638 20850 48690 20862
rect 49870 20914 49922 20926
rect 49870 20850 49922 20862
rect 9102 20802 9154 20814
rect 12910 20802 12962 20814
rect 14926 20802 14978 20814
rect 4946 20750 4958 20802
rect 5010 20750 5022 20802
rect 7970 20750 7982 20802
rect 8034 20750 8046 20802
rect 8530 20750 8542 20802
rect 8594 20750 8606 20802
rect 12338 20750 12350 20802
rect 12402 20750 12414 20802
rect 14354 20750 14366 20802
rect 14418 20750 14430 20802
rect 9102 20738 9154 20750
rect 12910 20738 12962 20750
rect 14926 20738 14978 20750
rect 15598 20802 15650 20814
rect 22318 20802 22370 20814
rect 29150 20802 29202 20814
rect 17378 20750 17390 20802
rect 17442 20750 17454 20802
rect 18050 20750 18062 20802
rect 18114 20750 18126 20802
rect 21522 20750 21534 20802
rect 21586 20750 21598 20802
rect 21746 20750 21758 20802
rect 21810 20750 21822 20802
rect 24546 20750 24558 20802
rect 24610 20750 24622 20802
rect 25666 20750 25678 20802
rect 25730 20750 25742 20802
rect 15598 20738 15650 20750
rect 22318 20738 22370 20750
rect 29150 20738 29202 20750
rect 30718 20802 30770 20814
rect 35422 20802 35474 20814
rect 42030 20802 42082 20814
rect 31042 20750 31054 20802
rect 31106 20750 31118 20802
rect 38434 20750 38446 20802
rect 38498 20750 38510 20802
rect 41570 20750 41582 20802
rect 41634 20750 41646 20802
rect 30718 20738 30770 20750
rect 35422 20738 35474 20750
rect 42030 20738 42082 20750
rect 42366 20802 42418 20814
rect 44930 20750 44942 20802
rect 44994 20750 45006 20802
rect 42366 20738 42418 20750
rect 2382 20690 2434 20702
rect 2382 20626 2434 20638
rect 2718 20690 2770 20702
rect 2718 20626 2770 20638
rect 3838 20690 3890 20702
rect 5966 20690 6018 20702
rect 11566 20690 11618 20702
rect 15262 20690 15314 20702
rect 4722 20638 4734 20690
rect 4786 20638 4798 20690
rect 8866 20638 8878 20690
rect 8930 20638 8942 20690
rect 12674 20638 12686 20690
rect 12738 20638 12750 20690
rect 14690 20638 14702 20690
rect 14754 20638 14766 20690
rect 3838 20626 3890 20638
rect 5966 20626 6018 20638
rect 11566 20626 11618 20638
rect 15262 20626 15314 20638
rect 19182 20690 19234 20702
rect 19182 20626 19234 20638
rect 21310 20690 21362 20702
rect 21310 20626 21362 20638
rect 23214 20690 23266 20702
rect 27022 20690 27074 20702
rect 25442 20638 25454 20690
rect 25506 20638 25518 20690
rect 35634 20638 35646 20690
rect 35698 20638 35710 20690
rect 35970 20638 35982 20690
rect 36034 20638 36046 20690
rect 39106 20638 39118 20690
rect 39170 20638 39182 20690
rect 23214 20626 23266 20638
rect 27022 20626 27074 20638
rect 5630 20578 5682 20590
rect 5630 20514 5682 20526
rect 8990 20578 9042 20590
rect 8990 20514 9042 20526
rect 11678 20578 11730 20590
rect 11678 20514 11730 20526
rect 12798 20578 12850 20590
rect 12798 20514 12850 20526
rect 14814 20578 14866 20590
rect 21982 20578 22034 20590
rect 17602 20526 17614 20578
rect 17666 20526 17678 20578
rect 18274 20526 18286 20578
rect 18338 20526 18350 20578
rect 18610 20526 18622 20578
rect 18674 20526 18686 20578
rect 14814 20514 14866 20526
rect 21982 20514 22034 20526
rect 22206 20578 22258 20590
rect 22206 20514 22258 20526
rect 22766 20578 22818 20590
rect 22766 20514 22818 20526
rect 23774 20578 23826 20590
rect 23774 20514 23826 20526
rect 26686 20578 26738 20590
rect 41582 20578 41634 20590
rect 29474 20526 29486 20578
rect 29538 20526 29550 20578
rect 26686 20514 26738 20526
rect 41582 20514 41634 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 17838 20242 17890 20254
rect 17838 20178 17890 20190
rect 23214 20242 23266 20254
rect 23214 20178 23266 20190
rect 41134 20242 41186 20254
rect 41134 20178 41186 20190
rect 45838 20242 45890 20254
rect 45838 20178 45890 20190
rect 47182 20242 47234 20254
rect 47182 20178 47234 20190
rect 9774 20130 9826 20142
rect 18286 20130 18338 20142
rect 22430 20130 22482 20142
rect 5506 20078 5518 20130
rect 5570 20078 5582 20130
rect 16370 20078 16382 20130
rect 16434 20078 16446 20130
rect 19954 20078 19966 20130
rect 20018 20078 20030 20130
rect 20850 20078 20862 20130
rect 20914 20078 20926 20130
rect 21298 20078 21310 20130
rect 21362 20078 21374 20130
rect 9774 20066 9826 20078
rect 18286 20066 18338 20078
rect 22430 20066 22482 20078
rect 23102 20130 23154 20142
rect 23102 20066 23154 20078
rect 23774 20130 23826 20142
rect 28926 20130 28978 20142
rect 30830 20130 30882 20142
rect 26338 20078 26350 20130
rect 26402 20078 26414 20130
rect 29474 20078 29486 20130
rect 29538 20078 29550 20130
rect 30034 20078 30046 20130
rect 30098 20078 30110 20130
rect 23774 20066 23826 20078
rect 28926 20066 28978 20078
rect 30830 20066 30882 20078
rect 33070 20130 33122 20142
rect 41582 20130 41634 20142
rect 34962 20078 34974 20130
rect 35026 20078 35038 20130
rect 33070 20066 33122 20078
rect 41582 20066 41634 20078
rect 41694 20130 41746 20142
rect 41694 20066 41746 20078
rect 15038 20018 15090 20030
rect 4834 19966 4846 20018
rect 4898 19966 4910 20018
rect 11890 19966 11902 20018
rect 11954 19966 11966 20018
rect 14354 19966 14366 20018
rect 14418 19966 14430 20018
rect 14914 19966 14926 20018
rect 14978 19966 14990 20018
rect 15038 19954 15090 19966
rect 15150 20018 15202 20030
rect 15710 20018 15762 20030
rect 18622 20018 18674 20030
rect 15474 19966 15486 20018
rect 15538 19966 15550 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 15150 19954 15202 19966
rect 15710 19954 15762 19966
rect 18622 19954 18674 19966
rect 19070 20018 19122 20030
rect 23438 20018 23490 20030
rect 33406 20018 33458 20030
rect 20178 19966 20190 20018
rect 20242 19966 20254 20018
rect 22642 19966 22654 20018
rect 22706 19966 22718 20018
rect 25554 19966 25566 20018
rect 25618 19966 25630 20018
rect 30594 19966 30606 20018
rect 30658 19966 30670 20018
rect 34290 19966 34302 20018
rect 34354 19966 34366 20018
rect 37426 19966 37438 20018
rect 37490 19966 37502 20018
rect 19070 19954 19122 19966
rect 23438 19954 23490 19966
rect 33406 19954 33458 19966
rect 8094 19906 8146 19918
rect 7634 19854 7646 19906
rect 7698 19854 7710 19906
rect 8094 19842 8146 19854
rect 8766 19906 8818 19918
rect 8766 19842 8818 19854
rect 9550 19906 9602 19918
rect 9550 19842 9602 19854
rect 21982 19906 22034 19918
rect 21982 19842 22034 19854
rect 24670 19906 24722 19918
rect 42142 19906 42194 19918
rect 28466 19854 28478 19906
rect 28530 19854 28542 19906
rect 37090 19854 37102 19906
rect 37154 19854 37166 19906
rect 39778 19854 39790 19906
rect 39842 19854 39854 19906
rect 24670 19842 24722 19854
rect 42142 19842 42194 19854
rect 9886 19794 9938 19806
rect 9886 19730 9938 19742
rect 11566 19794 11618 19806
rect 11566 19730 11618 19742
rect 11902 19794 11954 19806
rect 15934 19794 15986 19806
rect 14578 19742 14590 19794
rect 14642 19742 14654 19794
rect 11902 19730 11954 19742
rect 15934 19730 15986 19742
rect 16046 19794 16098 19806
rect 16046 19730 16098 19742
rect 19406 19794 19458 19806
rect 19406 19730 19458 19742
rect 21646 19794 21698 19806
rect 21646 19730 21698 19742
rect 29262 19794 29314 19806
rect 29262 19730 29314 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 6526 19458 6578 19470
rect 6526 19394 6578 19406
rect 6862 19458 6914 19470
rect 6862 19394 6914 19406
rect 10334 19458 10386 19470
rect 10334 19394 10386 19406
rect 14926 19458 14978 19470
rect 30718 19458 30770 19470
rect 16706 19406 16718 19458
rect 16770 19406 16782 19458
rect 14926 19394 14978 19406
rect 30718 19394 30770 19406
rect 37102 19346 37154 19358
rect 18274 19294 18286 19346
rect 18338 19294 18350 19346
rect 20402 19294 20414 19346
rect 20466 19294 20478 19346
rect 24210 19294 24222 19346
rect 24274 19294 24286 19346
rect 25442 19294 25454 19346
rect 25506 19294 25518 19346
rect 32498 19294 32510 19346
rect 32562 19294 32574 19346
rect 34626 19294 34638 19346
rect 34690 19294 34702 19346
rect 37102 19282 37154 19294
rect 10222 19234 10274 19246
rect 11566 19234 11618 19246
rect 14702 19234 14754 19246
rect 7634 19182 7646 19234
rect 7698 19182 7710 19234
rect 9314 19182 9326 19234
rect 9378 19182 9390 19234
rect 10658 19182 10670 19234
rect 10722 19182 10734 19234
rect 11890 19182 11902 19234
rect 11954 19182 11966 19234
rect 14466 19182 14478 19234
rect 14530 19182 14542 19234
rect 10222 19170 10274 19182
rect 11566 19170 11618 19182
rect 14702 19170 14754 19182
rect 15038 19234 15090 19246
rect 30382 19234 30434 19246
rect 35982 19234 36034 19246
rect 15698 19182 15710 19234
rect 15762 19182 15774 19234
rect 16146 19182 16158 19234
rect 16210 19182 16222 19234
rect 16482 19182 16494 19234
rect 16546 19182 16558 19234
rect 17490 19182 17502 19234
rect 17554 19182 17566 19234
rect 21298 19182 21310 19234
rect 21362 19182 21374 19234
rect 24994 19182 25006 19234
rect 25058 19182 25070 19234
rect 26002 19182 26014 19234
rect 26066 19182 26078 19234
rect 26450 19182 26462 19234
rect 26514 19182 26526 19234
rect 29698 19182 29710 19234
rect 29762 19182 29774 19234
rect 31826 19182 31838 19234
rect 31890 19182 31902 19234
rect 35298 19182 35310 19234
rect 35362 19182 35374 19234
rect 15038 19170 15090 19182
rect 30382 19170 30434 19182
rect 35982 19170 36034 19182
rect 2830 19122 2882 19134
rect 2830 19058 2882 19070
rect 3614 19122 3666 19134
rect 8206 19122 8258 19134
rect 7410 19070 7422 19122
rect 7474 19070 7486 19122
rect 3614 19058 3666 19070
rect 8206 19058 8258 19070
rect 8318 19122 8370 19134
rect 8318 19058 8370 19070
rect 8990 19122 9042 19134
rect 8990 19058 9042 19070
rect 9886 19122 9938 19134
rect 9886 19058 9938 19070
rect 11118 19122 11170 19134
rect 11330 19070 11342 19122
rect 11394 19070 11406 19122
rect 22082 19070 22094 19122
rect 22146 19070 22158 19122
rect 25666 19070 25678 19122
rect 25730 19070 25742 19122
rect 26786 19070 26798 19122
rect 26850 19070 26862 19122
rect 29810 19070 29822 19122
rect 29874 19070 29886 19122
rect 35410 19070 35422 19122
rect 35474 19070 35486 19122
rect 11118 19058 11170 19070
rect 2494 19010 2546 19022
rect 2494 18946 2546 18958
rect 3278 19010 3330 19022
rect 3278 18946 3330 18958
rect 5742 19010 5794 19022
rect 5742 18946 5794 18958
rect 7982 19010 8034 19022
rect 7982 18946 8034 18958
rect 9102 19010 9154 19022
rect 11902 19010 11954 19022
rect 10098 18958 10110 19010
rect 10162 18958 10174 19010
rect 9102 18946 9154 18958
rect 11902 18946 11954 18958
rect 24670 19010 24722 19022
rect 36318 19010 36370 19022
rect 27010 18958 27022 19010
rect 27074 18958 27086 19010
rect 24670 18946 24722 18958
rect 36318 18946 36370 18958
rect 37550 19010 37602 19022
rect 37550 18946 37602 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 8654 18674 8706 18686
rect 14142 18674 14194 18686
rect 25566 18674 25618 18686
rect 11442 18622 11454 18674
rect 11506 18622 11518 18674
rect 16370 18622 16382 18674
rect 16434 18622 16446 18674
rect 8654 18610 8706 18622
rect 14142 18610 14194 18622
rect 25566 18610 25618 18622
rect 26350 18674 26402 18686
rect 26350 18610 26402 18622
rect 38670 18674 38722 18686
rect 38670 18610 38722 18622
rect 9550 18562 9602 18574
rect 12910 18562 12962 18574
rect 20862 18562 20914 18574
rect 3042 18510 3054 18562
rect 3106 18510 3118 18562
rect 6514 18510 6526 18562
rect 6578 18510 6590 18562
rect 11218 18510 11230 18562
rect 11282 18510 11294 18562
rect 13570 18510 13582 18562
rect 13634 18510 13646 18562
rect 9550 18498 9602 18510
rect 12910 18498 12962 18510
rect 20862 18498 20914 18510
rect 27246 18562 27298 18574
rect 27246 18498 27298 18510
rect 27694 18562 27746 18574
rect 27694 18498 27746 18510
rect 27918 18562 27970 18574
rect 31042 18510 31054 18562
rect 31106 18510 31118 18562
rect 33730 18510 33742 18562
rect 33794 18510 33806 18562
rect 34066 18510 34078 18562
rect 34130 18510 34142 18562
rect 27918 18498 27970 18510
rect 5630 18450 5682 18462
rect 2258 18398 2270 18450
rect 2322 18398 2334 18450
rect 5630 18386 5682 18398
rect 5966 18450 6018 18462
rect 8430 18450 8482 18462
rect 6626 18398 6638 18450
rect 6690 18398 6702 18450
rect 5966 18386 6018 18398
rect 8430 18386 8482 18398
rect 8990 18450 9042 18462
rect 8990 18386 9042 18398
rect 9886 18450 9938 18462
rect 9886 18386 9938 18398
rect 9998 18450 10050 18462
rect 11006 18450 11058 18462
rect 13022 18450 13074 18462
rect 10322 18398 10334 18450
rect 10386 18398 10398 18450
rect 11554 18398 11566 18450
rect 11618 18398 11630 18450
rect 12338 18398 12350 18450
rect 12402 18398 12414 18450
rect 12786 18398 12798 18450
rect 12850 18398 12862 18450
rect 9998 18386 10050 18398
rect 11006 18386 11058 18398
rect 13022 18386 13074 18398
rect 13358 18450 13410 18462
rect 13358 18386 13410 18398
rect 13806 18450 13858 18462
rect 17390 18450 17442 18462
rect 21646 18450 21698 18462
rect 14130 18398 14142 18450
rect 14194 18398 14206 18450
rect 15922 18398 15934 18450
rect 15986 18398 15998 18450
rect 16146 18398 16158 18450
rect 16210 18398 16222 18450
rect 21186 18398 21198 18450
rect 21250 18398 21262 18450
rect 13806 18386 13858 18398
rect 17390 18386 17442 18398
rect 21646 18386 21698 18398
rect 24334 18450 24386 18462
rect 24334 18386 24386 18398
rect 25454 18450 25506 18462
rect 31826 18398 31838 18450
rect 31890 18398 31902 18450
rect 38210 18398 38222 18450
rect 38274 18398 38286 18450
rect 25454 18386 25506 18398
rect 9662 18338 9714 18350
rect 17950 18338 18002 18350
rect 5170 18286 5182 18338
rect 5234 18286 5246 18338
rect 16034 18286 16046 18338
rect 16098 18286 16110 18338
rect 9662 18274 9714 18286
rect 17950 18274 18002 18286
rect 18398 18338 18450 18350
rect 18398 18274 18450 18286
rect 23774 18338 23826 18350
rect 23774 18274 23826 18286
rect 24110 18338 24162 18350
rect 26798 18338 26850 18350
rect 32286 18338 32338 18350
rect 24658 18286 24670 18338
rect 24722 18286 24734 18338
rect 28914 18286 28926 18338
rect 28978 18286 28990 18338
rect 24110 18274 24162 18286
rect 26798 18274 26850 18286
rect 32286 18274 32338 18286
rect 33182 18338 33234 18350
rect 33182 18274 33234 18286
rect 34862 18338 34914 18350
rect 35298 18286 35310 18338
rect 35362 18286 35374 18338
rect 37426 18286 37438 18338
rect 37490 18286 37502 18338
rect 34862 18274 34914 18286
rect 17502 18226 17554 18238
rect 11554 18174 11566 18226
rect 11618 18174 11630 18226
rect 12450 18174 12462 18226
rect 12514 18174 12526 18226
rect 17502 18162 17554 18174
rect 21198 18226 21250 18238
rect 21198 18162 21250 18174
rect 27582 18226 27634 18238
rect 27582 18162 27634 18174
rect 33518 18226 33570 18238
rect 33518 18162 33570 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 5742 17890 5794 17902
rect 12574 17890 12626 17902
rect 7186 17838 7198 17890
rect 7250 17887 7262 17890
rect 7634 17887 7646 17890
rect 7250 17841 7646 17887
rect 7250 17838 7262 17841
rect 7634 17838 7646 17841
rect 7698 17838 7710 17890
rect 5742 17826 5794 17838
rect 12574 17826 12626 17838
rect 15710 17890 15762 17902
rect 15710 17826 15762 17838
rect 24894 17890 24946 17902
rect 24894 17826 24946 17838
rect 25790 17890 25842 17902
rect 25790 17826 25842 17838
rect 27582 17890 27634 17902
rect 27582 17826 27634 17838
rect 30158 17890 30210 17902
rect 30158 17826 30210 17838
rect 7646 17778 7698 17790
rect 2482 17726 2494 17778
rect 2546 17726 2558 17778
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 7646 17714 7698 17726
rect 15374 17778 15426 17790
rect 15374 17714 15426 17726
rect 16158 17778 16210 17790
rect 16158 17714 16210 17726
rect 27134 17778 27186 17790
rect 27906 17726 27918 17778
rect 27970 17726 27982 17778
rect 27134 17714 27186 17726
rect 6078 17666 6130 17678
rect 8318 17666 8370 17678
rect 12462 17666 12514 17678
rect 14366 17666 14418 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 6514 17614 6526 17666
rect 6578 17614 6590 17666
rect 8642 17614 8654 17666
rect 8706 17614 8718 17666
rect 9762 17614 9774 17666
rect 9826 17614 9838 17666
rect 12674 17614 12686 17666
rect 12738 17614 12750 17666
rect 14130 17614 14142 17666
rect 14194 17614 14206 17666
rect 6078 17602 6130 17614
rect 8318 17602 8370 17614
rect 12462 17602 12514 17614
rect 14366 17602 14418 17614
rect 14702 17666 14754 17678
rect 15598 17666 15650 17678
rect 17614 17666 17666 17678
rect 15138 17614 15150 17666
rect 15202 17614 15214 17666
rect 17154 17614 17166 17666
rect 17218 17614 17230 17666
rect 14702 17602 14754 17614
rect 15598 17602 15650 17614
rect 17614 17602 17666 17614
rect 23214 17666 23266 17678
rect 23214 17602 23266 17614
rect 23886 17666 23938 17678
rect 25342 17666 25394 17678
rect 24658 17614 24670 17666
rect 24722 17614 24734 17666
rect 23886 17602 23938 17614
rect 25342 17602 25394 17614
rect 26574 17666 26626 17678
rect 29810 17614 29822 17666
rect 29874 17614 29886 17666
rect 33842 17614 33854 17666
rect 33906 17614 33918 17666
rect 35858 17614 35870 17666
rect 35922 17614 35934 17666
rect 26574 17602 26626 17614
rect 7870 17554 7922 17566
rect 10334 17554 10386 17566
rect 6850 17502 6862 17554
rect 6914 17502 6926 17554
rect 8082 17502 8094 17554
rect 8146 17502 8158 17554
rect 8978 17502 8990 17554
rect 9042 17502 9054 17554
rect 9986 17502 9998 17554
rect 10050 17502 10062 17554
rect 7870 17490 7922 17502
rect 10334 17490 10386 17502
rect 10670 17554 10722 17566
rect 10670 17490 10722 17502
rect 12126 17554 12178 17566
rect 14814 17554 14866 17566
rect 14578 17502 14590 17554
rect 14642 17502 14654 17554
rect 12126 17490 12178 17502
rect 14814 17490 14866 17502
rect 16942 17554 16994 17566
rect 19518 17554 19570 17566
rect 16942 17490 16994 17502
rect 17950 17498 18002 17510
rect 5070 17442 5122 17454
rect 9326 17442 9378 17454
rect 8306 17390 8318 17442
rect 8370 17390 8382 17442
rect 5070 17378 5122 17390
rect 9326 17378 9378 17390
rect 11118 17442 11170 17454
rect 11118 17378 11170 17390
rect 12910 17442 12962 17454
rect 12910 17378 12962 17390
rect 16606 17442 16658 17454
rect 19518 17490 19570 17502
rect 23550 17554 23602 17566
rect 25678 17554 25730 17566
rect 25106 17502 25118 17554
rect 25170 17502 25182 17554
rect 23550 17490 23602 17502
rect 25678 17490 25730 17502
rect 36094 17554 36146 17566
rect 36094 17490 36146 17502
rect 17950 17434 18002 17446
rect 19182 17442 19234 17454
rect 25790 17442 25842 17454
rect 16606 17378 16658 17390
rect 24210 17390 24222 17442
rect 24274 17390 24286 17442
rect 24994 17390 25006 17442
rect 25058 17390 25070 17442
rect 19182 17378 19234 17390
rect 25790 17378 25842 17390
rect 27022 17442 27074 17454
rect 27022 17378 27074 17390
rect 27246 17442 27298 17454
rect 27246 17378 27298 17390
rect 27806 17442 27858 17454
rect 27806 17378 27858 17390
rect 30046 17442 30098 17454
rect 30046 17378 30098 17390
rect 34078 17442 34130 17454
rect 34078 17378 34130 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 6414 17106 6466 17118
rect 6414 17042 6466 17054
rect 6862 17106 6914 17118
rect 6862 17042 6914 17054
rect 7646 17106 7698 17118
rect 7646 17042 7698 17054
rect 8430 17106 8482 17118
rect 8430 17042 8482 17054
rect 8990 17106 9042 17118
rect 9886 17106 9938 17118
rect 9538 17054 9550 17106
rect 9602 17054 9614 17106
rect 8990 17042 9042 17054
rect 9886 17042 9938 17054
rect 10334 17106 10386 17118
rect 10334 17042 10386 17054
rect 11342 17106 11394 17118
rect 11342 17042 11394 17054
rect 16158 17106 16210 17118
rect 16158 17042 16210 17054
rect 21646 17106 21698 17118
rect 21646 17042 21698 17054
rect 25230 17106 25282 17118
rect 25230 17042 25282 17054
rect 26462 17106 26514 17118
rect 27918 17106 27970 17118
rect 27122 17054 27134 17106
rect 27186 17054 27198 17106
rect 26462 17042 26514 17054
rect 27918 17042 27970 17054
rect 36878 17106 36930 17118
rect 36878 17042 36930 17054
rect 2382 16994 2434 17006
rect 14814 16994 14866 17006
rect 16830 16994 16882 17006
rect 8082 16942 8094 16994
rect 8146 16942 8158 16994
rect 15138 16942 15150 16994
rect 15202 16942 15214 16994
rect 15810 16942 15822 16994
rect 15874 16942 15886 16994
rect 2382 16930 2434 16942
rect 14814 16930 14866 16942
rect 16830 16930 16882 16942
rect 17390 16994 17442 17006
rect 21758 16994 21810 17006
rect 26014 16994 26066 17006
rect 28702 16994 28754 17006
rect 19058 16942 19070 16994
rect 19122 16942 19134 16994
rect 23874 16942 23886 16994
rect 23938 16942 23950 16994
rect 27346 16942 27358 16994
rect 27410 16942 27422 16994
rect 17390 16930 17442 16942
rect 21758 16930 21810 16942
rect 26014 16930 26066 16942
rect 28702 16930 28754 16942
rect 30830 16994 30882 17006
rect 30830 16930 30882 16942
rect 31278 16994 31330 17006
rect 31938 16942 31950 16994
rect 32002 16942 32014 16994
rect 32386 16942 32398 16994
rect 32450 16942 32462 16994
rect 34290 16942 34302 16994
rect 34354 16942 34366 16994
rect 31278 16930 31330 16942
rect 2718 16882 2770 16894
rect 2718 16818 2770 16830
rect 6078 16882 6130 16894
rect 6078 16818 6130 16830
rect 6302 16882 6354 16894
rect 6302 16818 6354 16830
rect 6750 16882 6802 16894
rect 6750 16818 6802 16830
rect 11790 16882 11842 16894
rect 11790 16818 11842 16830
rect 12798 16882 12850 16894
rect 14478 16882 14530 16894
rect 13010 16830 13022 16882
rect 13074 16830 13086 16882
rect 13570 16830 13582 16882
rect 13634 16830 13646 16882
rect 12798 16818 12850 16830
rect 14478 16818 14530 16830
rect 15486 16882 15538 16894
rect 21422 16882 21474 16894
rect 27582 16882 27634 16894
rect 28366 16882 28418 16894
rect 16594 16830 16606 16882
rect 16658 16830 16670 16882
rect 17602 16830 17614 16882
rect 17666 16830 17678 16882
rect 18274 16830 18286 16882
rect 18338 16830 18350 16882
rect 22642 16830 22654 16882
rect 22706 16830 22718 16882
rect 25218 16830 25230 16882
rect 25282 16830 25294 16882
rect 25778 16830 25790 16882
rect 25842 16830 25854 16882
rect 26898 16830 26910 16882
rect 26962 16830 26974 16882
rect 28018 16830 28030 16882
rect 28082 16830 28094 16882
rect 30594 16830 30606 16882
rect 30658 16830 30670 16882
rect 33618 16830 33630 16882
rect 33682 16830 33694 16882
rect 15486 16818 15538 16830
rect 21422 16818 21474 16830
rect 27582 16818 27634 16830
rect 28366 16818 28418 16830
rect 7422 16770 7474 16782
rect 10894 16770 10946 16782
rect 7746 16718 7758 16770
rect 7810 16718 7822 16770
rect 7422 16706 7474 16718
rect 10894 16706 10946 16718
rect 11230 16770 11282 16782
rect 11230 16706 11282 16718
rect 12910 16770 12962 16782
rect 12910 16706 12962 16718
rect 13246 16770 13298 16782
rect 13246 16706 13298 16718
rect 14702 16770 14754 16782
rect 27134 16770 27186 16782
rect 21186 16718 21198 16770
rect 21250 16718 21262 16770
rect 36418 16718 36430 16770
rect 36482 16718 36494 16770
rect 14702 16706 14754 16718
rect 27134 16706 27186 16718
rect 14366 16658 14418 16670
rect 14366 16594 14418 16606
rect 25566 16658 25618 16670
rect 31614 16658 31666 16670
rect 28130 16606 28142 16658
rect 28194 16606 28206 16658
rect 25566 16594 25618 16606
rect 31614 16594 31666 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 5742 16322 5794 16334
rect 5742 16258 5794 16270
rect 6078 16322 6130 16334
rect 6078 16258 6130 16270
rect 19518 16322 19570 16334
rect 19518 16258 19570 16270
rect 19854 16322 19906 16334
rect 19854 16258 19906 16270
rect 28142 16322 28194 16334
rect 28142 16258 28194 16270
rect 29598 16322 29650 16334
rect 29598 16258 29650 16270
rect 34190 16322 34242 16334
rect 34190 16258 34242 16270
rect 16046 16210 16098 16222
rect 2482 16158 2494 16210
rect 2546 16158 2558 16210
rect 4610 16158 4622 16210
rect 4674 16158 4686 16210
rect 11106 16158 11118 16210
rect 11170 16158 11182 16210
rect 16046 16146 16098 16158
rect 21534 16210 21586 16222
rect 21534 16146 21586 16158
rect 24222 16210 24274 16222
rect 24222 16146 24274 16158
rect 26238 16210 26290 16222
rect 30818 16158 30830 16210
rect 30882 16158 30894 16210
rect 32946 16158 32958 16210
rect 33010 16158 33022 16210
rect 26238 16146 26290 16158
rect 11902 16098 11954 16110
rect 1810 16046 1822 16098
rect 1874 16046 1886 16098
rect 6850 16046 6862 16098
rect 6914 16046 6926 16098
rect 8194 16046 8206 16098
rect 8258 16046 8270 16098
rect 11902 16034 11954 16046
rect 14254 16098 14306 16110
rect 16382 16098 16434 16110
rect 14802 16046 14814 16098
rect 14866 16046 14878 16098
rect 14254 16034 14306 16046
rect 16382 16034 16434 16046
rect 17502 16098 17554 16110
rect 19070 16098 19122 16110
rect 22766 16098 22818 16110
rect 18050 16046 18062 16098
rect 18114 16046 18126 16098
rect 20514 16046 20526 16098
rect 20578 16046 20590 16098
rect 17502 16034 17554 16046
rect 19070 16034 19122 16046
rect 22766 16034 22818 16046
rect 23438 16098 23490 16110
rect 23438 16034 23490 16046
rect 24334 16098 24386 16110
rect 24334 16034 24386 16046
rect 25678 16098 25730 16110
rect 27022 16098 27074 16110
rect 34526 16098 34578 16110
rect 26674 16046 26686 16098
rect 26738 16046 26750 16098
rect 27234 16046 27246 16098
rect 27298 16046 27310 16098
rect 27906 16046 27918 16098
rect 27970 16046 27982 16098
rect 33618 16046 33630 16098
rect 33682 16046 33694 16098
rect 35858 16046 35870 16098
rect 35922 16046 35934 16098
rect 25678 16034 25730 16046
rect 27022 16034 27074 16046
rect 34526 16034 34578 16046
rect 7422 15986 7474 15998
rect 6738 15934 6750 15986
rect 6802 15934 6814 15986
rect 7422 15922 7474 15934
rect 7646 15986 7698 15998
rect 7646 15922 7698 15934
rect 7758 15986 7810 15998
rect 15262 15986 15314 15998
rect 8978 15934 8990 15986
rect 9042 15934 9054 15986
rect 12226 15934 12238 15986
rect 12290 15934 12302 15986
rect 12450 15934 12462 15986
rect 12514 15934 12526 15986
rect 13906 15934 13918 15986
rect 13970 15934 13982 15986
rect 14578 15934 14590 15986
rect 14642 15934 14654 15986
rect 7758 15922 7810 15934
rect 15262 15922 15314 15934
rect 15598 15986 15650 15998
rect 24558 15986 24610 15998
rect 16706 15934 16718 15986
rect 16770 15934 16782 15986
rect 18274 15934 18286 15986
rect 18338 15934 18350 15986
rect 20402 15934 20414 15986
rect 20466 15934 20478 15986
rect 15598 15922 15650 15934
rect 24558 15922 24610 15934
rect 27470 15986 27522 15998
rect 28590 15986 28642 15998
rect 28354 15934 28366 15986
rect 28418 15934 28430 15986
rect 29810 15934 29822 15986
rect 29874 15934 29886 15986
rect 30370 15934 30382 15986
rect 30434 15934 30446 15986
rect 34738 15934 34750 15986
rect 34802 15934 34814 15986
rect 35074 15934 35086 15986
rect 35138 15934 35150 15986
rect 27470 15922 27522 15934
rect 28590 15922 28642 15934
rect 5070 15874 5122 15886
rect 5070 15810 5122 15822
rect 11566 15874 11618 15886
rect 11566 15810 11618 15822
rect 15934 15874 15986 15886
rect 21982 15874 22034 15886
rect 24110 15874 24162 15886
rect 17154 15822 17166 15874
rect 17218 15822 17230 15874
rect 18722 15822 18734 15874
rect 18786 15822 18798 15874
rect 23090 15822 23102 15874
rect 23154 15822 23166 15874
rect 23762 15822 23774 15874
rect 23826 15822 23838 15874
rect 15934 15810 15986 15822
rect 21982 15810 22034 15822
rect 24110 15810 24162 15822
rect 25006 15874 25058 15886
rect 26126 15874 26178 15886
rect 25330 15822 25342 15874
rect 25394 15822 25406 15874
rect 25006 15810 25058 15822
rect 26126 15810 26178 15822
rect 26350 15874 26402 15886
rect 26350 15810 26402 15822
rect 26686 15874 26738 15886
rect 29262 15874 29314 15886
rect 28130 15822 28142 15874
rect 28194 15822 28206 15874
rect 26686 15810 26738 15822
rect 29262 15810 29314 15822
rect 36094 15874 36146 15886
rect 36094 15810 36146 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 12574 15538 12626 15550
rect 12574 15474 12626 15486
rect 12798 15538 12850 15550
rect 12798 15474 12850 15486
rect 13470 15538 13522 15550
rect 13470 15474 13522 15486
rect 14478 15538 14530 15550
rect 14478 15474 14530 15486
rect 14926 15538 14978 15550
rect 14926 15474 14978 15486
rect 17838 15538 17890 15550
rect 17838 15474 17890 15486
rect 19406 15538 19458 15550
rect 23662 15538 23714 15550
rect 23314 15486 23326 15538
rect 23378 15486 23390 15538
rect 19406 15474 19458 15486
rect 23662 15474 23714 15486
rect 24222 15538 24274 15550
rect 24222 15474 24274 15486
rect 24446 15538 24498 15550
rect 24446 15474 24498 15486
rect 25342 15538 25394 15550
rect 25342 15474 25394 15486
rect 25566 15538 25618 15550
rect 25566 15474 25618 15486
rect 26686 15538 26738 15550
rect 30942 15538 30994 15550
rect 28242 15486 28254 15538
rect 28306 15486 28318 15538
rect 26686 15474 26738 15486
rect 30942 15474 30994 15486
rect 33406 15538 33458 15550
rect 33406 15474 33458 15486
rect 33854 15538 33906 15550
rect 33854 15474 33906 15486
rect 38782 15538 38834 15550
rect 38782 15474 38834 15486
rect 20078 15426 20130 15438
rect 25790 15426 25842 15438
rect 10322 15374 10334 15426
rect 10386 15374 10398 15426
rect 12002 15374 12014 15426
rect 12066 15374 12078 15426
rect 20514 15374 20526 15426
rect 20578 15374 20590 15426
rect 20078 15362 20130 15374
rect 25790 15362 25842 15374
rect 27470 15426 27522 15438
rect 28018 15374 28030 15426
rect 28082 15374 28094 15426
rect 31490 15374 31502 15426
rect 31554 15374 31566 15426
rect 31826 15374 31838 15426
rect 31890 15374 31902 15426
rect 34850 15374 34862 15426
rect 34914 15374 34926 15426
rect 37538 15374 37550 15426
rect 37602 15374 37614 15426
rect 27470 15362 27522 15374
rect 11454 15314 11506 15326
rect 12910 15314 12962 15326
rect 21646 15314 21698 15326
rect 2930 15262 2942 15314
rect 2994 15262 3006 15314
rect 6962 15262 6974 15314
rect 7026 15262 7038 15314
rect 10434 15262 10446 15314
rect 10498 15262 10510 15314
rect 12226 15262 12238 15314
rect 12290 15262 12302 15314
rect 19842 15262 19854 15314
rect 19906 15262 19918 15314
rect 20626 15262 20638 15314
rect 20690 15262 20702 15314
rect 11454 15250 11506 15262
rect 12910 15250 12962 15262
rect 21646 15250 21698 15262
rect 24558 15314 24610 15326
rect 24558 15250 24610 15262
rect 24670 15314 24722 15326
rect 24670 15250 24722 15262
rect 25230 15314 25282 15326
rect 25230 15250 25282 15262
rect 26350 15314 26402 15326
rect 27134 15314 27186 15326
rect 26674 15262 26686 15314
rect 26738 15262 26750 15314
rect 26350 15250 26402 15262
rect 27134 15250 27186 15262
rect 27806 15314 27858 15326
rect 27806 15250 27858 15262
rect 28254 15314 28306 15326
rect 28354 15262 28366 15314
rect 28418 15262 28430 15314
rect 34962 15262 34974 15314
rect 35026 15262 35038 15314
rect 38322 15262 38334 15314
rect 38386 15262 38398 15314
rect 28254 15250 28306 15262
rect 13918 15202 13970 15214
rect 3602 15150 3614 15202
rect 3666 15150 3678 15202
rect 5730 15150 5742 15202
rect 5794 15150 5806 15202
rect 8194 15150 8206 15202
rect 8258 15150 8270 15202
rect 9762 15150 9774 15202
rect 9826 15150 9838 15202
rect 13918 15138 13970 15150
rect 15598 15202 15650 15214
rect 15598 15138 15650 15150
rect 31278 15202 31330 15214
rect 31278 15138 31330 15150
rect 34190 15202 34242 15214
rect 35410 15150 35422 15202
rect 35474 15150 35486 15202
rect 34190 15138 34242 15150
rect 11118 15090 11170 15102
rect 11118 15026 11170 15038
rect 21310 15090 21362 15102
rect 26898 15038 26910 15090
rect 26962 15038 26974 15090
rect 21310 15026 21362 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 11006 14754 11058 14766
rect 11006 14690 11058 14702
rect 11678 14754 11730 14766
rect 11678 14690 11730 14702
rect 15150 14754 15202 14766
rect 27358 14754 27410 14766
rect 26786 14702 26798 14754
rect 26850 14702 26862 14754
rect 15150 14690 15202 14702
rect 27358 14690 27410 14702
rect 36206 14754 36258 14766
rect 36206 14690 36258 14702
rect 10894 14642 10946 14654
rect 9874 14590 9886 14642
rect 9938 14590 9950 14642
rect 10894 14578 10946 14590
rect 15374 14642 15426 14654
rect 24670 14642 24722 14654
rect 22082 14590 22094 14642
rect 22146 14590 22158 14642
rect 24210 14590 24222 14642
rect 24274 14590 24286 14642
rect 15374 14578 15426 14590
rect 24670 14578 24722 14590
rect 5966 14530 6018 14542
rect 12014 14530 12066 14542
rect 16494 14530 16546 14542
rect 7074 14478 7086 14530
rect 7138 14478 7150 14530
rect 13794 14478 13806 14530
rect 13858 14478 13870 14530
rect 5966 14466 6018 14478
rect 12014 14466 12066 14478
rect 16494 14466 16546 14478
rect 16830 14530 16882 14542
rect 25006 14530 25058 14542
rect 21410 14478 21422 14530
rect 21474 14478 21486 14530
rect 16830 14466 16882 14478
rect 25006 14466 25058 14478
rect 26126 14530 26178 14542
rect 27694 14530 27746 14542
rect 35870 14530 35922 14542
rect 26338 14478 26350 14530
rect 26402 14478 26414 14530
rect 28354 14478 28366 14530
rect 28418 14478 28430 14530
rect 30370 14478 30382 14530
rect 30434 14478 30446 14530
rect 26126 14466 26178 14478
rect 27694 14466 27746 14478
rect 35870 14466 35922 14478
rect 3838 14418 3890 14430
rect 3838 14354 3890 14366
rect 4174 14418 4226 14430
rect 10222 14418 10274 14430
rect 7746 14366 7758 14418
rect 7810 14366 7822 14418
rect 4174 14354 4226 14366
rect 10222 14354 10274 14366
rect 10558 14418 10610 14430
rect 15934 14418 15986 14430
rect 12226 14366 12238 14418
rect 12290 14366 12302 14418
rect 12562 14366 12574 14418
rect 12626 14366 12638 14418
rect 14130 14366 14142 14418
rect 14194 14366 14206 14418
rect 10558 14354 10610 14366
rect 15934 14354 15986 14366
rect 25566 14418 25618 14430
rect 28466 14366 28478 14418
rect 28530 14366 28542 14418
rect 35074 14366 35086 14418
rect 35138 14366 35150 14418
rect 35522 14366 35534 14418
rect 35586 14366 35598 14418
rect 25566 14354 25618 14366
rect 30606 14306 30658 14318
rect 13570 14254 13582 14306
rect 13634 14254 13646 14306
rect 14802 14254 14814 14306
rect 14866 14254 14878 14306
rect 17154 14254 17166 14306
rect 17218 14254 17230 14306
rect 30606 14242 30658 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 6190 13970 6242 13982
rect 6190 13906 6242 13918
rect 7982 13970 8034 13982
rect 7982 13906 8034 13918
rect 9102 13970 9154 13982
rect 9102 13906 9154 13918
rect 12798 13970 12850 13982
rect 12798 13906 12850 13918
rect 13470 13970 13522 13982
rect 13470 13906 13522 13918
rect 13806 13970 13858 13982
rect 13806 13906 13858 13918
rect 15934 13970 15986 13982
rect 15934 13906 15986 13918
rect 25342 13970 25394 13982
rect 27134 13970 27186 13982
rect 26562 13918 26574 13970
rect 26626 13918 26638 13970
rect 25342 13906 25394 13918
rect 27134 13906 27186 13918
rect 3054 13858 3106 13870
rect 3054 13794 3106 13806
rect 3726 13858 3778 13870
rect 8318 13858 8370 13870
rect 7186 13806 7198 13858
rect 7250 13806 7262 13858
rect 3726 13794 3778 13806
rect 8318 13794 8370 13806
rect 12910 13858 12962 13870
rect 17390 13858 17442 13870
rect 14466 13806 14478 13858
rect 14530 13806 14542 13858
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 19170 13806 19182 13858
rect 19234 13806 19246 13858
rect 27682 13806 27694 13858
rect 27746 13806 27758 13858
rect 31714 13806 31726 13858
rect 31778 13806 31790 13858
rect 34290 13806 34302 13858
rect 34354 13806 34366 13858
rect 12910 13794 12962 13806
rect 17390 13794 17442 13806
rect 4062 13746 4114 13758
rect 3266 13694 3278 13746
rect 3330 13694 3342 13746
rect 4062 13682 4114 13694
rect 6526 13746 6578 13758
rect 17726 13746 17778 13758
rect 26462 13746 26514 13758
rect 7298 13694 7310 13746
rect 7362 13694 7374 13746
rect 9986 13694 9998 13746
rect 10050 13694 10062 13746
rect 19394 13694 19406 13746
rect 19458 13694 19470 13746
rect 20850 13694 20862 13746
rect 20914 13694 20926 13746
rect 21186 13694 21198 13746
rect 21250 13694 21262 13746
rect 26002 13694 26014 13746
rect 26066 13694 26078 13746
rect 6526 13682 6578 13694
rect 17726 13682 17778 13694
rect 26462 13682 26514 13694
rect 26798 13746 26850 13758
rect 27918 13746 27970 13758
rect 33182 13746 33234 13758
rect 27122 13694 27134 13746
rect 27186 13694 27198 13746
rect 32498 13694 32510 13746
rect 32562 13694 32574 13746
rect 26798 13682 26850 13694
rect 27918 13682 27970 13694
rect 33182 13682 33234 13694
rect 33518 13746 33570 13758
rect 33954 13694 33966 13746
rect 34018 13694 34030 13746
rect 33518 13682 33570 13694
rect 5294 13634 5346 13646
rect 18286 13634 18338 13646
rect 24446 13634 24498 13646
rect 10658 13582 10670 13634
rect 10722 13582 10734 13634
rect 22306 13582 22318 13634
rect 22370 13582 22382 13634
rect 5294 13570 5346 13582
rect 18286 13570 18338 13582
rect 24446 13570 24498 13582
rect 27470 13634 27522 13646
rect 29586 13582 29598 13634
rect 29650 13582 29662 13634
rect 27470 13570 27522 13582
rect 12798 13522 12850 13534
rect 12798 13458 12850 13470
rect 14142 13522 14194 13534
rect 14142 13458 14194 13470
rect 18622 13522 18674 13534
rect 18622 13458 18674 13470
rect 20526 13522 20578 13534
rect 20526 13458 20578 13470
rect 20862 13522 20914 13534
rect 20862 13458 20914 13470
rect 26350 13522 26402 13534
rect 26350 13458 26402 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 5742 13186 5794 13198
rect 5742 13122 5794 13134
rect 19742 13186 19794 13198
rect 19742 13122 19794 13134
rect 22094 13186 22146 13198
rect 27918 13186 27970 13198
rect 22978 13134 22990 13186
rect 23042 13134 23054 13186
rect 25554 13134 25566 13186
rect 25618 13134 25630 13186
rect 27346 13134 27358 13186
rect 27410 13134 27422 13186
rect 22094 13122 22146 13134
rect 27918 13122 27970 13134
rect 30382 13186 30434 13198
rect 30382 13122 30434 13134
rect 35198 13186 35250 13198
rect 35198 13122 35250 13134
rect 35534 13186 35586 13198
rect 35534 13122 35586 13134
rect 8542 13074 8594 13086
rect 12462 13074 12514 13086
rect 23438 13074 23490 13086
rect 2818 13022 2830 13074
rect 2882 13022 2894 13074
rect 4946 13022 4958 13074
rect 5010 13022 5022 13074
rect 11666 13022 11678 13074
rect 11730 13022 11742 13074
rect 19394 13022 19406 13074
rect 19458 13022 19470 13074
rect 8542 13010 8594 13022
rect 12462 13010 12514 13022
rect 23438 13010 23490 13022
rect 26238 13074 26290 13086
rect 26238 13010 26290 13022
rect 26910 13074 26962 13086
rect 26910 13010 26962 13022
rect 32734 13074 32786 13086
rect 32734 13010 32786 13022
rect 6078 12962 6130 12974
rect 13918 12962 13970 12974
rect 20078 12962 20130 12974
rect 2034 12910 2046 12962
rect 2098 12910 2110 12962
rect 8866 12910 8878 12962
rect 8930 12910 8942 12962
rect 16594 12910 16606 12962
rect 16658 12910 16670 12962
rect 6078 12898 6130 12910
rect 13918 12898 13970 12910
rect 20078 12898 20130 12910
rect 21982 12962 22034 12974
rect 24222 12962 24274 12974
rect 22306 12910 22318 12962
rect 22370 12910 22382 12962
rect 22754 12910 22766 12962
rect 22818 12910 22830 12962
rect 23314 12910 23326 12962
rect 23378 12910 23390 12962
rect 21982 12898 22034 12910
rect 24222 12898 24274 12910
rect 24334 12962 24386 12974
rect 25118 12962 25170 12974
rect 24434 12910 24446 12962
rect 24498 12910 24510 12962
rect 24334 12898 24386 12910
rect 25118 12898 25170 12910
rect 25342 12962 25394 12974
rect 29598 12962 29650 12974
rect 30718 12962 30770 12974
rect 25666 12910 25678 12962
rect 25730 12910 25742 12962
rect 26450 12910 26462 12962
rect 26514 12910 26526 12962
rect 27346 12910 27358 12962
rect 27410 12910 27422 12962
rect 29362 12910 29374 12962
rect 29426 12910 29438 12962
rect 29698 12910 29710 12962
rect 29762 12910 29774 12962
rect 31490 12910 31502 12962
rect 31554 12910 31566 12962
rect 33170 12910 33182 12962
rect 33234 12910 33246 12962
rect 25342 12898 25394 12910
rect 29598 12898 29650 12910
rect 30718 12898 30770 12910
rect 20302 12850 20354 12862
rect 6402 12798 6414 12850
rect 6466 12798 6478 12850
rect 6850 12798 6862 12850
rect 6914 12798 6926 12850
rect 9538 12798 9550 12850
rect 9602 12798 9614 12850
rect 14130 12798 14142 12850
rect 14194 12798 14206 12850
rect 14466 12798 14478 12850
rect 14530 12798 14542 12850
rect 17266 12798 17278 12850
rect 17330 12798 17342 12850
rect 20302 12786 20354 12798
rect 21646 12850 21698 12862
rect 21646 12786 21698 12798
rect 23550 12850 23602 12862
rect 23550 12786 23602 12798
rect 23886 12850 23938 12862
rect 23886 12786 23938 12798
rect 25006 12850 25058 12862
rect 25006 12786 25058 12798
rect 26126 12850 26178 12862
rect 26126 12786 26178 12798
rect 26798 12850 26850 12862
rect 28030 12850 28082 12862
rect 27010 12798 27022 12850
rect 27074 12798 27086 12850
rect 26798 12786 26850 12798
rect 28030 12786 28082 12798
rect 28254 12850 28306 12862
rect 28254 12786 28306 12798
rect 29150 12850 29202 12862
rect 31266 12798 31278 12850
rect 31330 12798 31342 12850
rect 35746 12798 35758 12850
rect 35810 12798 35822 12850
rect 36306 12798 36318 12850
rect 36370 12798 36382 12850
rect 29150 12786 29202 12798
rect 12798 12738 12850 12750
rect 12798 12674 12850 12686
rect 13582 12738 13634 12750
rect 13582 12674 13634 12686
rect 20750 12738 20802 12750
rect 20750 12674 20802 12686
rect 22430 12738 22482 12750
rect 22430 12674 22482 12686
rect 24670 12738 24722 12750
rect 24670 12674 24722 12686
rect 29934 12738 29986 12750
rect 29934 12674 29986 12686
rect 33406 12738 33458 12750
rect 33406 12674 33458 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 5070 12402 5122 12414
rect 5070 12338 5122 12350
rect 9886 12402 9938 12414
rect 9886 12338 9938 12350
rect 16830 12402 16882 12414
rect 16830 12338 16882 12350
rect 18062 12402 18114 12414
rect 18062 12338 18114 12350
rect 21646 12402 21698 12414
rect 21646 12338 21698 12350
rect 22990 12402 23042 12414
rect 22990 12338 23042 12350
rect 23438 12402 23490 12414
rect 23438 12338 23490 12350
rect 25790 12402 25842 12414
rect 25790 12338 25842 12350
rect 29262 12402 29314 12414
rect 39678 12402 39730 12414
rect 29922 12350 29934 12402
rect 29986 12350 29998 12402
rect 29262 12338 29314 12350
rect 39678 12338 39730 12350
rect 10558 12290 10610 12302
rect 2482 12238 2494 12290
rect 2546 12238 2558 12290
rect 6066 12238 6078 12290
rect 6130 12238 6142 12290
rect 10558 12226 10610 12238
rect 10894 12290 10946 12302
rect 16494 12290 16546 12302
rect 29598 12290 29650 12302
rect 12898 12238 12910 12290
rect 12962 12238 12974 12290
rect 13346 12238 13358 12290
rect 13410 12238 13422 12290
rect 18946 12238 18958 12290
rect 19010 12238 19022 12290
rect 24098 12238 24110 12290
rect 24162 12238 24174 12290
rect 24434 12238 24446 12290
rect 24498 12238 24510 12290
rect 33842 12238 33854 12290
rect 33906 12238 33918 12290
rect 10894 12226 10946 12238
rect 16494 12226 16546 12238
rect 29598 12226 29650 12238
rect 5406 12178 5458 12190
rect 10222 12178 10274 12190
rect 1810 12126 1822 12178
rect 1874 12126 1886 12178
rect 6178 12126 6190 12178
rect 6242 12126 6254 12178
rect 5406 12114 5458 12126
rect 10222 12114 10274 12126
rect 12350 12178 12402 12190
rect 12350 12114 12402 12126
rect 18398 12178 18450 12190
rect 27918 12178 27970 12190
rect 19170 12126 19182 12178
rect 19234 12126 19246 12178
rect 27010 12126 27022 12178
rect 27074 12126 27086 12178
rect 33058 12126 33070 12178
rect 33122 12126 33134 12178
rect 39106 12126 39118 12178
rect 39170 12126 39182 12178
rect 18398 12114 18450 12126
rect 27918 12114 27970 12126
rect 12686 12066 12738 12078
rect 4610 12014 4622 12066
rect 4674 12014 4686 12066
rect 12686 12002 12738 12014
rect 19742 12066 19794 12078
rect 19742 12002 19794 12014
rect 21534 12066 21586 12078
rect 21534 12002 21586 12014
rect 22878 12066 22930 12078
rect 26350 12066 26402 12078
rect 27470 12066 27522 12078
rect 25330 12014 25342 12066
rect 25394 12014 25406 12066
rect 26898 12014 26910 12066
rect 26962 12014 26974 12066
rect 35970 12014 35982 12066
rect 36034 12014 36046 12066
rect 36306 12014 36318 12066
rect 36370 12014 36382 12066
rect 38434 12014 38446 12066
rect 38498 12014 38510 12066
rect 22878 12002 22930 12014
rect 26350 12002 26402 12014
rect 27470 12002 27522 12014
rect 23774 11954 23826 11966
rect 23774 11890 23826 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 15150 11618 15202 11630
rect 15150 11554 15202 11566
rect 19854 11618 19906 11630
rect 19854 11554 19906 11566
rect 27582 11618 27634 11630
rect 27582 11554 27634 11566
rect 30382 11618 30434 11630
rect 30382 11554 30434 11566
rect 33294 11618 33346 11630
rect 33294 11554 33346 11566
rect 33630 11618 33682 11630
rect 33630 11554 33682 11566
rect 35534 11618 35586 11630
rect 35534 11554 35586 11566
rect 4846 11506 4898 11518
rect 8990 11506 9042 11518
rect 12910 11506 12962 11518
rect 23438 11506 23490 11518
rect 8530 11454 8542 11506
rect 8594 11454 8606 11506
rect 10322 11454 10334 11506
rect 10386 11454 10398 11506
rect 12450 11454 12462 11506
rect 12514 11454 12526 11506
rect 16370 11454 16382 11506
rect 16434 11454 16446 11506
rect 18498 11454 18510 11506
rect 18562 11454 18574 11506
rect 4846 11442 4898 11454
rect 8990 11442 9042 11454
rect 12910 11442 12962 11454
rect 23438 11442 23490 11454
rect 24334 11506 24386 11518
rect 24334 11442 24386 11454
rect 24558 11506 24610 11518
rect 24558 11442 24610 11454
rect 37102 11506 37154 11518
rect 37102 11442 37154 11454
rect 14814 11394 14866 11406
rect 25454 11394 25506 11406
rect 26462 11394 26514 11406
rect 5618 11342 5630 11394
rect 5682 11342 5694 11394
rect 9538 11342 9550 11394
rect 9602 11342 9614 11394
rect 15698 11342 15710 11394
rect 15762 11342 15774 11394
rect 20290 11342 20302 11394
rect 20354 11342 20366 11394
rect 23986 11342 23998 11394
rect 24050 11342 24062 11394
rect 25890 11342 25902 11394
rect 25954 11342 25966 11394
rect 26674 11342 26686 11394
rect 26738 11342 26750 11394
rect 29586 11342 29598 11394
rect 29650 11342 29662 11394
rect 14814 11330 14866 11342
rect 25454 11330 25506 11342
rect 26462 11330 26514 11342
rect 27246 11282 27298 11294
rect 6402 11230 6414 11282
rect 6466 11230 6478 11282
rect 14018 11230 14030 11282
rect 14082 11230 14094 11282
rect 14578 11230 14590 11282
rect 14642 11230 14654 11282
rect 20626 11230 20638 11282
rect 20690 11230 20702 11282
rect 27246 11218 27298 11230
rect 27694 11282 27746 11294
rect 27694 11218 27746 11230
rect 29262 11282 29314 11294
rect 30594 11230 30606 11282
rect 30658 11230 30670 11282
rect 30930 11230 30942 11282
rect 30994 11230 31006 11282
rect 33842 11230 33854 11282
rect 33906 11230 33918 11282
rect 34290 11230 34302 11282
rect 34354 11230 34366 11282
rect 35746 11230 35758 11282
rect 35810 11230 35822 11282
rect 36306 11230 36318 11282
rect 36370 11230 36382 11282
rect 29262 11218 29314 11230
rect 19070 11170 19122 11182
rect 19070 11106 19122 11118
rect 19518 11170 19570 11182
rect 19518 11106 19570 11118
rect 26126 11170 26178 11182
rect 26126 11106 26178 11118
rect 29374 11170 29426 11182
rect 29374 11106 29426 11118
rect 30046 11170 30098 11182
rect 30046 11106 30098 11118
rect 35198 11170 35250 11182
rect 35198 11106 35250 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 6302 10834 6354 10846
rect 6302 10770 6354 10782
rect 13134 10834 13186 10846
rect 13134 10770 13186 10782
rect 17838 10834 17890 10846
rect 17838 10770 17890 10782
rect 18958 10834 19010 10846
rect 18958 10770 19010 10782
rect 29598 10834 29650 10846
rect 29598 10770 29650 10782
rect 29934 10834 29986 10846
rect 35982 10834 36034 10846
rect 30258 10782 30270 10834
rect 30322 10782 30334 10834
rect 29934 10770 29986 10782
rect 35982 10770 36034 10782
rect 14030 10722 14082 10734
rect 18174 10722 18226 10734
rect 35646 10722 35698 10734
rect 7970 10670 7982 10722
rect 8034 10670 8046 10722
rect 12450 10670 12462 10722
rect 12514 10670 12526 10722
rect 16258 10670 16270 10722
rect 16322 10670 16334 10722
rect 24322 10670 24334 10722
rect 24386 10670 24398 10722
rect 26450 10670 26462 10722
rect 26514 10670 26526 10722
rect 30818 10670 30830 10722
rect 30882 10670 30894 10722
rect 14030 10658 14082 10670
rect 18174 10658 18226 10670
rect 35646 10658 35698 10670
rect 6638 10610 6690 10622
rect 6638 10546 6690 10558
rect 7086 10610 7138 10622
rect 7086 10546 7138 10558
rect 7422 10610 7474 10622
rect 14366 10610 14418 10622
rect 8194 10558 8206 10610
rect 8258 10558 8270 10610
rect 12562 10558 12574 10610
rect 12626 10558 12638 10610
rect 7422 10546 7474 10558
rect 14366 10546 14418 10558
rect 16606 10610 16658 10622
rect 24670 10610 24722 10622
rect 31502 10610 31554 10622
rect 18386 10558 18398 10610
rect 18450 10558 18462 10610
rect 19058 10558 19070 10610
rect 19122 10558 19134 10610
rect 20066 10558 20078 10610
rect 20130 10558 20142 10610
rect 25666 10558 25678 10610
rect 25730 10558 25742 10610
rect 30706 10558 30718 10610
rect 30770 10558 30782 10610
rect 16606 10546 16658 10558
rect 24670 10546 24722 10558
rect 31502 10546 31554 10558
rect 15486 10498 15538 10510
rect 23326 10498 23378 10510
rect 19282 10446 19294 10498
rect 19346 10446 19358 10498
rect 20738 10446 20750 10498
rect 20802 10446 20814 10498
rect 22866 10446 22878 10498
rect 22930 10446 22942 10498
rect 15486 10434 15538 10446
rect 23326 10434 23378 10446
rect 25342 10498 25394 10510
rect 28578 10446 28590 10498
rect 28642 10446 28654 10498
rect 25342 10434 25394 10446
rect 11454 10386 11506 10398
rect 11454 10322 11506 10334
rect 11790 10386 11842 10398
rect 11790 10322 11842 10334
rect 31838 10386 31890 10398
rect 31838 10322 31890 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 12462 10050 12514 10062
rect 12462 9986 12514 9998
rect 12798 10050 12850 10062
rect 12798 9986 12850 9998
rect 26462 10050 26514 10062
rect 26462 9986 26514 9998
rect 16942 9938 16994 9950
rect 25006 9938 25058 9950
rect 14242 9886 14254 9938
rect 14306 9886 14318 9938
rect 16370 9886 16382 9938
rect 16434 9886 16446 9938
rect 17938 9886 17950 9938
rect 18002 9886 18014 9938
rect 20066 9886 20078 9938
rect 20130 9886 20142 9938
rect 16942 9874 16994 9886
rect 25006 9874 25058 9886
rect 26014 9938 26066 9950
rect 26014 9874 26066 9886
rect 7646 9826 7698 9838
rect 20414 9826 20466 9838
rect 6626 9774 6638 9826
rect 6690 9774 6702 9826
rect 8082 9774 8094 9826
rect 8146 9774 8158 9826
rect 13458 9774 13470 9826
rect 13522 9774 13534 9826
rect 17266 9774 17278 9826
rect 17330 9774 17342 9826
rect 7646 9762 7698 9774
rect 20414 9762 20466 9774
rect 22318 9826 22370 9838
rect 22318 9762 22370 9774
rect 26798 9826 26850 9838
rect 27346 9774 27358 9826
rect 27410 9774 27422 9826
rect 29922 9774 29934 9826
rect 29986 9774 29998 9826
rect 31042 9774 31054 9826
rect 31106 9774 31118 9826
rect 26798 9762 26850 9774
rect 7310 9714 7362 9726
rect 20750 9714 20802 9726
rect 8306 9662 8318 9714
rect 8370 9662 8382 9714
rect 11890 9662 11902 9714
rect 11954 9662 11966 9714
rect 12226 9662 12238 9714
rect 12290 9662 12302 9714
rect 22530 9662 22542 9714
rect 22594 9662 22606 9714
rect 23090 9662 23102 9714
rect 23154 9662 23166 9714
rect 27570 9662 27582 9714
rect 27634 9662 27646 9714
rect 7310 9650 7362 9662
rect 20750 9650 20802 9662
rect 6862 9602 6914 9614
rect 6862 9538 6914 9550
rect 21982 9602 22034 9614
rect 21982 9538 22034 9550
rect 25566 9602 25618 9614
rect 25566 9538 25618 9550
rect 30158 9602 30210 9614
rect 30158 9538 30210 9550
rect 31278 9602 31330 9614
rect 31278 9538 31330 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 14366 9266 14418 9278
rect 14366 9202 14418 9214
rect 18398 9266 18450 9278
rect 18398 9202 18450 9214
rect 20526 9266 20578 9278
rect 20526 9202 20578 9214
rect 28590 9266 28642 9278
rect 28590 9202 28642 9214
rect 33182 9266 33234 9278
rect 33182 9202 33234 9214
rect 27582 9154 27634 9166
rect 6850 9102 6862 9154
rect 6914 9102 6926 9154
rect 13122 9102 13134 9154
rect 13186 9102 13198 9154
rect 15474 9102 15486 9154
rect 15538 9102 15550 9154
rect 18946 9102 18958 9154
rect 19010 9102 19022 9154
rect 19506 9102 19518 9154
rect 19570 9102 19582 9154
rect 25778 9102 25790 9154
rect 25842 9102 25854 9154
rect 31378 9102 31390 9154
rect 31442 9102 31454 9154
rect 27582 9090 27634 9102
rect 27022 9042 27074 9054
rect 6066 8990 6078 9042
rect 6130 8990 6142 9042
rect 9538 8990 9550 9042
rect 9602 8990 9614 9042
rect 12898 8990 12910 9042
rect 12962 8990 12974 9042
rect 15362 8990 15374 9042
rect 15426 8990 15438 9042
rect 24546 8990 24558 9042
rect 24610 8990 24622 9042
rect 26002 8990 26014 9042
rect 26066 8990 26078 9042
rect 26674 8990 26686 9042
rect 26738 8990 26750 9042
rect 27794 8990 27806 9042
rect 27858 8990 27870 9042
rect 32162 8990 32174 9042
rect 32226 8990 32238 9042
rect 27022 8978 27074 8990
rect 13694 8930 13746 8942
rect 8978 8878 8990 8930
rect 9042 8878 9054 8930
rect 10322 8878 10334 8930
rect 10386 8878 10398 8930
rect 12450 8878 12462 8930
rect 12514 8878 12526 8930
rect 13694 8866 13746 8878
rect 20078 8930 20130 8942
rect 20078 8866 20130 8878
rect 21310 8930 21362 8942
rect 25566 8930 25618 8942
rect 21746 8878 21758 8930
rect 21810 8878 21822 8930
rect 23874 8878 23886 8930
rect 23938 8878 23950 8930
rect 21310 8866 21362 8878
rect 25566 8866 25618 8878
rect 27246 8930 27298 8942
rect 27246 8866 27298 8878
rect 28478 8930 28530 8942
rect 29250 8878 29262 8930
rect 29314 8878 29326 8930
rect 28478 8866 28530 8878
rect 14702 8818 14754 8830
rect 14702 8754 14754 8766
rect 18734 8818 18786 8830
rect 18734 8754 18786 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 9214 8370 9266 8382
rect 9214 8306 9266 8318
rect 13582 8370 13634 8382
rect 13582 8306 13634 8318
rect 22430 8370 22482 8382
rect 22430 8306 22482 8318
rect 25230 8370 25282 8382
rect 26450 8318 26462 8370
rect 26514 8318 26526 8370
rect 28578 8318 28590 8370
rect 28642 8318 28654 8370
rect 30706 8318 30718 8370
rect 30770 8318 30782 8370
rect 32834 8318 32846 8370
rect 32898 8318 32910 8370
rect 25230 8306 25282 8318
rect 10670 8258 10722 8270
rect 10670 8194 10722 8206
rect 13918 8258 13970 8270
rect 18510 8258 18562 8270
rect 18274 8206 18286 8258
rect 18338 8206 18350 8258
rect 13918 8194 13970 8206
rect 18510 8194 18562 8206
rect 19182 8258 19234 8270
rect 19182 8194 19234 8206
rect 19630 8258 19682 8270
rect 19630 8194 19682 8206
rect 20078 8258 20130 8270
rect 20078 8194 20130 8206
rect 20414 8258 20466 8270
rect 23662 8258 23714 8270
rect 21858 8206 21870 8258
rect 21922 8206 21934 8258
rect 22306 8206 22318 8258
rect 22370 8206 22382 8258
rect 22978 8206 22990 8258
rect 23042 8206 23054 8258
rect 20414 8194 20466 8206
rect 23662 8194 23714 8206
rect 23998 8258 24050 8270
rect 34190 8258 34242 8270
rect 24658 8206 24670 8258
rect 24722 8206 24734 8258
rect 25666 8206 25678 8258
rect 25730 8206 25742 8258
rect 33618 8206 33630 8258
rect 33682 8206 33694 8258
rect 23998 8194 24050 8206
rect 34190 8194 34242 8206
rect 10334 8146 10386 8158
rect 17726 8146 17778 8158
rect 14130 8094 14142 8146
rect 14194 8094 14206 8146
rect 14690 8094 14702 8146
rect 14754 8094 14766 8146
rect 10334 8082 10386 8094
rect 17726 8082 17778 8094
rect 18846 8146 18898 8158
rect 24446 8146 24498 8158
rect 22866 8094 22878 8146
rect 22930 8094 22942 8146
rect 18846 8082 18898 8094
rect 24446 8082 24498 8094
rect 12686 8034 12738 8046
rect 12686 7970 12738 7982
rect 20750 8034 20802 8046
rect 20750 7970 20802 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 19182 7698 19234 7710
rect 19182 7634 19234 7646
rect 24110 7698 24162 7710
rect 24110 7634 24162 7646
rect 24670 7698 24722 7710
rect 24670 7634 24722 7646
rect 25342 7698 25394 7710
rect 25342 7634 25394 7646
rect 26798 7698 26850 7710
rect 26798 7634 26850 7646
rect 16494 7586 16546 7598
rect 13346 7534 13358 7586
rect 13410 7534 13422 7586
rect 18498 7534 18510 7586
rect 18562 7534 18574 7586
rect 20962 7534 20974 7586
rect 21026 7534 21038 7586
rect 27346 7534 27358 7586
rect 27410 7534 27422 7586
rect 27906 7534 27918 7586
rect 27970 7534 27982 7586
rect 16494 7522 16546 7534
rect 12574 7474 12626 7486
rect 16830 7474 16882 7486
rect 13234 7422 13246 7474
rect 13298 7422 13310 7474
rect 12574 7410 12626 7422
rect 16830 7410 16882 7422
rect 17502 7474 17554 7486
rect 17502 7410 17554 7422
rect 17838 7474 17890 7486
rect 24222 7474 24274 7486
rect 18274 7422 18286 7474
rect 18338 7422 18350 7474
rect 20290 7422 20302 7474
rect 20354 7422 20366 7474
rect 23986 7422 23998 7474
rect 24050 7422 24062 7474
rect 17838 7410 17890 7422
rect 24222 7410 24274 7422
rect 27134 7474 27186 7486
rect 27134 7410 27186 7422
rect 23090 7310 23102 7362
rect 23154 7310 23166 7362
rect 12238 7250 12290 7262
rect 12238 7186 12290 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 14366 6914 14418 6926
rect 14366 6850 14418 6862
rect 23550 6914 23602 6926
rect 23550 6850 23602 6862
rect 22766 6802 22818 6814
rect 12898 6750 12910 6802
rect 12962 6750 12974 6802
rect 16370 6750 16382 6802
rect 16434 6750 16446 6802
rect 18498 6750 18510 6802
rect 18562 6750 18574 6802
rect 22766 6738 22818 6750
rect 24894 6802 24946 6814
rect 24894 6738 24946 6750
rect 13582 6690 13634 6702
rect 18958 6690 19010 6702
rect 10098 6638 10110 6690
rect 10162 6638 10174 6690
rect 14802 6638 14814 6690
rect 14866 6638 14878 6690
rect 15698 6638 15710 6690
rect 15762 6638 15774 6690
rect 13582 6626 13634 6638
rect 18958 6626 19010 6638
rect 23214 6690 23266 6702
rect 28590 6690 28642 6702
rect 23986 6638 23998 6690
rect 24050 6638 24062 6690
rect 23214 6626 23266 6638
rect 28590 6626 28642 6638
rect 26910 6578 26962 6590
rect 10770 6526 10782 6578
rect 10834 6526 10846 6578
rect 15026 6526 15038 6578
rect 15090 6526 15102 6578
rect 24322 6526 24334 6578
rect 24386 6526 24398 6578
rect 26910 6514 26962 6526
rect 28478 6578 28530 6590
rect 28478 6514 28530 6526
rect 14030 6466 14082 6478
rect 14030 6402 14082 6414
rect 22206 6466 22258 6478
rect 22206 6402 22258 6414
rect 27246 6466 27298 6478
rect 27246 6402 27298 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 11230 6130 11282 6142
rect 11230 6066 11282 6078
rect 14926 6130 14978 6142
rect 14926 6066 14978 6078
rect 26350 6130 26402 6142
rect 26350 6066 26402 6078
rect 26798 6130 26850 6142
rect 26798 6066 26850 6078
rect 13470 6018 13522 6030
rect 13470 5954 13522 5966
rect 13806 6018 13858 6030
rect 16830 6018 16882 6030
rect 16034 5966 16046 6018
rect 16098 5966 16110 6018
rect 18274 5966 18286 6018
rect 18338 5966 18350 6018
rect 18498 5966 18510 6018
rect 18562 5966 18574 6018
rect 22530 5966 22542 6018
rect 22594 5966 22606 6018
rect 24322 5966 24334 6018
rect 24386 5966 24398 6018
rect 27906 5966 27918 6018
rect 27970 5966 27982 6018
rect 13806 5954 13858 5966
rect 16830 5954 16882 5966
rect 15262 5906 15314 5918
rect 16494 5906 16546 5918
rect 11442 5854 11454 5906
rect 11506 5854 11518 5906
rect 15922 5854 15934 5906
rect 15986 5854 15998 5906
rect 15262 5842 15314 5854
rect 16494 5842 16546 5854
rect 17614 5906 17666 5918
rect 17614 5842 17666 5854
rect 17950 5906 18002 5918
rect 17950 5842 18002 5854
rect 21870 5906 21922 5918
rect 23550 5906 23602 5918
rect 27134 5906 27186 5918
rect 22642 5854 22654 5906
rect 22706 5854 22718 5906
rect 24210 5854 24222 5906
rect 24274 5854 24286 5906
rect 27570 5854 27582 5906
rect 27634 5854 27646 5906
rect 21870 5842 21922 5854
rect 23550 5842 23602 5854
rect 27134 5842 27186 5854
rect 25342 5794 25394 5806
rect 25342 5730 25394 5742
rect 25790 5794 25842 5806
rect 25790 5730 25842 5742
rect 26238 5794 26290 5806
rect 26238 5730 26290 5742
rect 21534 5682 21586 5694
rect 21534 5618 21586 5630
rect 23214 5682 23266 5694
rect 23214 5618 23266 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 16270 5234 16322 5246
rect 19854 5234 19906 5246
rect 17266 5182 17278 5234
rect 17330 5182 17342 5234
rect 19394 5182 19406 5234
rect 19458 5182 19470 5234
rect 24994 5182 25006 5234
rect 25058 5182 25070 5234
rect 28242 5182 28254 5234
rect 28306 5182 28318 5234
rect 16270 5170 16322 5182
rect 19854 5170 19906 5182
rect 16594 5070 16606 5122
rect 16658 5070 16670 5122
rect 20514 5070 20526 5122
rect 20578 5070 20590 5122
rect 21522 5070 21534 5122
rect 21586 5070 21598 5122
rect 22082 5070 22094 5122
rect 22146 5070 22158 5122
rect 22866 5070 22878 5122
rect 22930 5070 22942 5122
rect 25330 5070 25342 5122
rect 25394 5070 25406 5122
rect 21758 5010 21810 5022
rect 26114 4958 26126 5010
rect 26178 4958 26190 5010
rect 21758 4946 21810 4958
rect 20750 4898 20802 4910
rect 20750 4834 20802 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 12238 4562 12290 4574
rect 12238 4498 12290 4510
rect 24222 4562 24274 4574
rect 24222 4498 24274 4510
rect 25678 4562 25730 4574
rect 25678 4498 25730 4510
rect 26014 4562 26066 4574
rect 26014 4498 26066 4510
rect 13346 4398 13358 4450
rect 13410 4398 13422 4450
rect 27458 4398 27470 4450
rect 27522 4398 27534 4450
rect 12562 4286 12574 4338
rect 12626 4286 12638 4338
rect 20850 4286 20862 4338
rect 20914 4286 20926 4338
rect 26226 4286 26238 4338
rect 26290 4286 26302 4338
rect 26674 4286 26686 4338
rect 26738 4286 26750 4338
rect 15474 4174 15486 4226
rect 15538 4174 15550 4226
rect 21634 4174 21646 4226
rect 21698 4174 21710 4226
rect 23762 4174 23774 4226
rect 23826 4174 23838 4226
rect 29586 4174 29598 4226
rect 29650 4174 29662 4226
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 26238 3778 26290 3790
rect 26238 3714 26290 3726
rect 26574 3778 26626 3790
rect 26574 3714 26626 3726
rect 27234 3502 27246 3554
rect 27298 3502 27310 3554
rect 27122 3390 27134 3442
rect 27186 3390 27198 3442
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 15150 57038 15202 57090
rect 16046 57038 16098 57090
rect 44382 57038 44434 57090
rect 44942 57038 44994 57090
rect 12574 56590 12626 56642
rect 13134 56590 13186 56642
rect 18510 56590 18562 56642
rect 18958 56590 19010 56642
rect 22094 56590 22146 56642
rect 22878 56590 22930 56642
rect 23662 56590 23714 56642
rect 24222 56590 24274 56642
rect 27358 56590 27410 56642
rect 28366 56590 28418 56642
rect 29486 56590 29538 56642
rect 30046 56590 30098 56642
rect 39230 56590 39282 56642
rect 39902 56590 39954 56642
rect 54238 56590 54290 56642
rect 55022 56590 55074 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4622 56254 4674 56306
rect 4958 56254 5010 56306
rect 6974 56254 7026 56306
rect 8206 56254 8258 56306
rect 9662 56254 9714 56306
rect 11006 56254 11058 56306
rect 12350 56254 12402 56306
rect 13694 56254 13746 56306
rect 14702 56254 14754 56306
rect 15150 56254 15202 56306
rect 15598 56254 15650 56306
rect 15934 56254 15986 56306
rect 18286 56254 18338 56306
rect 24670 56254 24722 56306
rect 27022 56254 27074 56306
rect 28366 56254 28418 56306
rect 28926 56254 28978 56306
rect 29486 56254 29538 56306
rect 31502 56254 31554 56306
rect 35310 56254 35362 56306
rect 39118 56254 39170 56306
rect 43598 56254 43650 56306
rect 44942 56254 44994 56306
rect 45950 56254 46002 56306
rect 47406 56254 47458 56306
rect 48638 56254 48690 56306
rect 49982 56254 50034 56306
rect 51326 56254 51378 56306
rect 52670 56254 52722 56306
rect 54014 56254 54066 56306
rect 55470 56254 55522 56306
rect 5518 56142 5570 56194
rect 5854 56142 5906 56194
rect 16270 56142 16322 56194
rect 17278 56142 17330 56194
rect 17614 56142 17666 56194
rect 18622 56142 18674 56194
rect 18958 56142 19010 56194
rect 19854 56142 19906 56194
rect 22094 56142 22146 56194
rect 23662 56142 23714 56194
rect 20078 56030 20130 56082
rect 21198 56030 21250 56082
rect 22766 56030 22818 56082
rect 26126 56030 26178 56082
rect 27806 56030 27858 56082
rect 30270 56030 30322 56082
rect 32174 56030 32226 56082
rect 33742 56030 33794 56082
rect 35982 56030 36034 56082
rect 37550 56030 37602 56082
rect 39790 56030 39842 56082
rect 42590 56030 42642 56082
rect 6190 55918 6242 55970
rect 7422 55918 7474 55970
rect 8654 55918 8706 55970
rect 10110 55918 10162 55970
rect 11454 55918 11506 55970
rect 13134 55918 13186 55970
rect 14142 55918 14194 55970
rect 19406 55918 19458 55970
rect 20750 55918 20802 55970
rect 25566 55918 25618 55970
rect 29934 55918 29986 55970
rect 30718 55918 30770 55970
rect 32622 55918 32674 55970
rect 34190 55918 34242 55970
rect 36430 55918 36482 55970
rect 37998 55918 38050 55970
rect 40462 55918 40514 55970
rect 42030 55918 42082 55970
rect 42926 55918 42978 55970
rect 44046 55918 44098 55970
rect 44494 55918 44546 55970
rect 46398 55918 46450 55970
rect 47854 55918 47906 55970
rect 49086 55918 49138 55970
rect 50430 55918 50482 55970
rect 51774 55918 51826 55970
rect 53118 55918 53170 55970
rect 55022 55918 55074 55970
rect 55918 55918 55970 55970
rect 45390 55806 45442 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 15486 55470 15538 55522
rect 16158 55470 16210 55522
rect 19182 55470 19234 55522
rect 4622 55358 4674 55410
rect 5854 55358 5906 55410
rect 14814 55358 14866 55410
rect 18510 55358 18562 55410
rect 20078 55358 20130 55410
rect 22430 55358 22482 55410
rect 28590 55358 28642 55410
rect 32062 55358 32114 55410
rect 35310 55358 35362 55410
rect 37438 55358 37490 55410
rect 39678 55358 39730 55410
rect 1822 55246 1874 55298
rect 8766 55246 8818 55298
rect 15262 55246 15314 55298
rect 16494 55246 16546 55298
rect 17166 55246 17218 55298
rect 17390 55246 17442 55298
rect 17838 55246 17890 55298
rect 25230 55246 25282 55298
rect 25790 55246 25842 55298
rect 29150 55246 29202 55298
rect 32510 55246 32562 55298
rect 38110 55246 38162 55298
rect 39118 55246 39170 55298
rect 42590 55246 42642 55298
rect 2494 55134 2546 55186
rect 7982 55134 8034 55186
rect 16606 55134 16658 55186
rect 16830 55134 16882 55186
rect 17950 55134 18002 55186
rect 18286 55134 18338 55186
rect 20414 55134 20466 55186
rect 21646 55134 21698 55186
rect 22094 55134 22146 55186
rect 24558 55134 24610 55186
rect 26462 55134 26514 55186
rect 29934 55134 29986 55186
rect 33182 55134 33234 55186
rect 35982 55134 36034 55186
rect 36318 55134 36370 55186
rect 38558 55134 38610 55186
rect 41806 55134 41858 55186
rect 42926 55134 42978 55186
rect 43038 55134 43090 55186
rect 43374 55134 43426 55186
rect 5070 55022 5122 55074
rect 9214 55022 9266 55074
rect 17054 55022 17106 55074
rect 18846 55022 18898 55074
rect 35646 55022 35698 55074
rect 39342 55022 39394 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 2494 54686 2546 54738
rect 16830 54686 16882 54738
rect 19182 54686 19234 54738
rect 19294 54686 19346 54738
rect 20190 54686 20242 54738
rect 26238 54686 26290 54738
rect 29262 54686 29314 54738
rect 30046 54686 30098 54738
rect 33070 54686 33122 54738
rect 39678 54686 39730 54738
rect 40238 54686 40290 54738
rect 40910 54686 40962 54738
rect 2382 54574 2434 54626
rect 7534 54574 7586 54626
rect 19742 54574 19794 54626
rect 24446 54574 24498 54626
rect 35646 54574 35698 54626
rect 2606 54462 2658 54514
rect 2942 54462 2994 54514
rect 3390 54462 3442 54514
rect 4398 54462 4450 54514
rect 6526 54462 6578 54514
rect 6974 54462 7026 54514
rect 7310 54462 7362 54514
rect 12126 54462 12178 54514
rect 12462 54462 12514 54514
rect 16270 54462 16322 54514
rect 17838 54462 17890 54514
rect 18286 54462 18338 54514
rect 18622 54462 18674 54514
rect 19070 54462 19122 54514
rect 19518 54462 19570 54514
rect 23102 54462 23154 54514
rect 23886 54462 23938 54514
rect 24334 54462 24386 54514
rect 28590 54462 28642 54514
rect 30382 54462 30434 54514
rect 34526 54462 34578 54514
rect 34862 54462 34914 54514
rect 39230 54462 39282 54514
rect 45502 54462 45554 54514
rect 3278 54350 3330 54402
rect 4958 54350 5010 54402
rect 6750 54350 6802 54402
rect 7646 54350 7698 54402
rect 13246 54350 13298 54402
rect 15374 54350 15426 54402
rect 20974 54350 21026 54402
rect 25342 54350 25394 54402
rect 25790 54350 25842 54402
rect 29710 54350 29762 54402
rect 32062 54350 32114 54402
rect 32510 54350 32562 54402
rect 37774 54350 37826 54402
rect 42702 54350 42754 54402
rect 44830 54350 44882 54402
rect 16494 54238 16546 54290
rect 24222 54238 24274 54290
rect 39118 54238 39170 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 13470 53902 13522 53954
rect 17166 53902 17218 53954
rect 24558 53902 24610 53954
rect 4622 53790 4674 53842
rect 9550 53790 9602 53842
rect 12798 53790 12850 53842
rect 13582 53790 13634 53842
rect 17390 53790 17442 53842
rect 20750 53790 20802 53842
rect 23774 53790 23826 53842
rect 33742 53790 33794 53842
rect 34190 53790 34242 53842
rect 35198 53790 35250 53842
rect 38558 53790 38610 53842
rect 39566 53790 39618 53842
rect 45950 53790 46002 53842
rect 51550 53790 51602 53842
rect 1822 53678 1874 53730
rect 9998 53678 10050 53730
rect 10670 53678 10722 53730
rect 17502 53678 17554 53730
rect 17838 53678 17890 53730
rect 22206 53678 22258 53730
rect 22878 53678 22930 53730
rect 24558 53678 24610 53730
rect 30942 53678 30994 53730
rect 38670 53678 38722 53730
rect 38782 53678 38834 53730
rect 39118 53678 39170 53730
rect 42254 53678 42306 53730
rect 42814 53678 42866 53730
rect 48750 53678 48802 53730
rect 2494 53566 2546 53618
rect 18622 53566 18674 53618
rect 23326 53566 23378 53618
rect 23550 53566 23602 53618
rect 23886 53566 23938 53618
rect 24222 53566 24274 53618
rect 31614 53566 31666 53618
rect 35534 53566 35586 53618
rect 35870 53566 35922 53618
rect 35982 53566 36034 53618
rect 37774 53566 37826 53618
rect 39454 53566 39506 53618
rect 39678 53566 39730 53618
rect 39790 53566 39842 53618
rect 39902 53566 39954 53618
rect 43374 53566 43426 53618
rect 43710 53566 43762 53618
rect 46286 53566 46338 53618
rect 49422 53566 49474 53618
rect 5070 53454 5122 53506
rect 13694 53454 13746 53506
rect 16830 53454 16882 53506
rect 25006 53454 25058 53506
rect 35310 53454 35362 53506
rect 36206 53454 36258 53506
rect 37886 53454 37938 53506
rect 38110 53454 38162 53506
rect 38446 53454 38498 53506
rect 46062 53454 46114 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 2718 53118 2770 53170
rect 3502 53118 3554 53170
rect 18846 53118 18898 53170
rect 19406 53118 19458 53170
rect 23886 53118 23938 53170
rect 24670 53118 24722 53170
rect 30830 53118 30882 53170
rect 31950 53118 32002 53170
rect 33966 53118 34018 53170
rect 34078 53118 34130 53170
rect 34302 53118 34354 53170
rect 34750 53118 34802 53170
rect 36878 53118 36930 53170
rect 39454 53118 39506 53170
rect 41022 53118 41074 53170
rect 42142 53118 42194 53170
rect 42590 53118 42642 53170
rect 49086 53118 49138 53170
rect 4398 53006 4450 53058
rect 8094 53006 8146 53058
rect 12910 53006 12962 53058
rect 18174 53006 18226 53058
rect 25454 53006 25506 53058
rect 26014 53006 26066 53058
rect 28254 53006 28306 53058
rect 38894 53006 38946 53058
rect 40238 53006 40290 53058
rect 41806 53006 41858 53058
rect 43038 53006 43090 53058
rect 45726 53006 45778 53058
rect 2942 52894 2994 52946
rect 3278 52894 3330 52946
rect 3614 52894 3666 52946
rect 3838 52894 3890 52946
rect 4286 52894 4338 52946
rect 4510 52894 4562 52946
rect 11454 52894 11506 52946
rect 12462 52894 12514 52946
rect 13470 52894 13522 52946
rect 13806 52894 13858 52946
rect 14030 52894 14082 52946
rect 18510 52894 18562 52946
rect 19182 52894 19234 52946
rect 19854 52894 19906 52946
rect 20078 52894 20130 52946
rect 23550 52894 23602 52946
rect 23774 52894 23826 52946
rect 23998 52894 24050 52946
rect 24222 52894 24274 52946
rect 27582 52894 27634 52946
rect 32286 52894 32338 52946
rect 34526 52894 34578 52946
rect 35198 52894 35250 52946
rect 35646 52894 35698 52946
rect 36206 52894 36258 52946
rect 37214 52894 37266 52946
rect 38110 52894 38162 52946
rect 38670 52894 38722 52946
rect 39006 52894 39058 52946
rect 41134 52894 41186 52946
rect 42478 52894 42530 52946
rect 43486 52894 43538 52946
rect 43934 52894 43986 52946
rect 45054 52894 45106 52946
rect 48862 52894 48914 52946
rect 49982 52894 50034 52946
rect 10334 52782 10386 52834
rect 10894 52782 10946 52834
rect 12014 52782 12066 52834
rect 13582 52782 13634 52834
rect 16606 52782 16658 52834
rect 17726 52782 17778 52834
rect 18734 52782 18786 52834
rect 19294 52782 19346 52834
rect 20862 52782 20914 52834
rect 22990 52782 23042 52834
rect 30382 52782 30434 52834
rect 35982 52782 36034 52834
rect 38446 52782 38498 52834
rect 39678 52782 39730 52834
rect 47854 52782 47906 52834
rect 49198 52782 49250 52834
rect 49534 52782 49586 52834
rect 49870 52782 49922 52834
rect 2606 52670 2658 52722
rect 4958 52670 5010 52722
rect 10558 52670 10610 52722
rect 11566 52670 11618 52722
rect 16494 52670 16546 52722
rect 17950 52670 18002 52722
rect 25230 52670 25282 52722
rect 25566 52670 25618 52722
rect 35422 52670 35474 52722
rect 36430 52670 36482 52722
rect 37662 52670 37714 52722
rect 37886 52670 37938 52722
rect 40014 52670 40066 52722
rect 41022 52670 41074 52722
rect 42590 52670 42642 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 4398 52334 4450 52386
rect 20638 52334 20690 52386
rect 37998 52334 38050 52386
rect 39342 52334 39394 52386
rect 40798 52334 40850 52386
rect 41246 52334 41298 52386
rect 49870 52334 49922 52386
rect 50542 52334 50594 52386
rect 7982 52222 8034 52274
rect 11342 52222 11394 52274
rect 18286 52222 18338 52274
rect 20190 52222 20242 52274
rect 24558 52222 24610 52274
rect 25006 52222 25058 52274
rect 27134 52222 27186 52274
rect 33294 52222 33346 52274
rect 33742 52222 33794 52274
rect 36094 52222 36146 52274
rect 38446 52222 38498 52274
rect 41806 52222 41858 52274
rect 46174 52222 46226 52274
rect 49422 52222 49474 52274
rect 4174 52110 4226 52162
rect 4622 52110 4674 52162
rect 6302 52110 6354 52162
rect 6414 52110 6466 52162
rect 6638 52110 6690 52162
rect 6862 52110 6914 52162
rect 7198 52110 7250 52162
rect 8542 52110 8594 52162
rect 12574 52110 12626 52162
rect 12798 52110 12850 52162
rect 12910 52110 12962 52162
rect 13694 52110 13746 52162
rect 13806 52110 13858 52162
rect 13918 52110 13970 52162
rect 14814 52110 14866 52162
rect 15486 52110 15538 52162
rect 18734 52110 18786 52162
rect 19182 52110 19234 52162
rect 19742 52110 19794 52162
rect 20750 52110 20802 52162
rect 23102 52110 23154 52162
rect 23550 52110 23602 52162
rect 24446 52110 24498 52162
rect 27918 52110 27970 52162
rect 30494 52110 30546 52162
rect 31166 52110 31218 52162
rect 39454 52110 39506 52162
rect 40126 52110 40178 52162
rect 40910 52110 40962 52162
rect 41246 52110 41298 52162
rect 42030 52110 42082 52162
rect 47406 52110 47458 52162
rect 47854 52110 47906 52162
rect 50542 52110 50594 52162
rect 50766 52110 50818 52162
rect 51886 52110 51938 52162
rect 7534 51998 7586 52050
rect 9214 51998 9266 52050
rect 16158 51998 16210 52050
rect 20638 51998 20690 52050
rect 23998 51998 24050 52050
rect 35758 51998 35810 52050
rect 36206 51998 36258 52050
rect 38110 51998 38162 52050
rect 38558 51998 38610 52050
rect 38782 51998 38834 52050
rect 39790 51998 39842 52050
rect 41582 51998 41634 52050
rect 42142 51998 42194 52050
rect 42702 51998 42754 52050
rect 49758 51998 49810 52050
rect 51102 51998 51154 52050
rect 51438 51998 51490 52050
rect 4286 51886 4338 51938
rect 5854 51886 5906 51938
rect 7086 51886 7138 51938
rect 14366 51886 14418 51938
rect 15038 51886 15090 51938
rect 24222 51886 24274 51938
rect 24558 51886 24610 51938
rect 28366 51886 28418 51938
rect 35982 51886 36034 51938
rect 37998 51886 38050 51938
rect 39006 51886 39058 51938
rect 40798 51886 40850 51938
rect 46734 51886 46786 51938
rect 47070 51886 47122 51938
rect 47742 51886 47794 51938
rect 49310 51886 49362 51938
rect 49870 51886 49922 51938
rect 50990 51886 51042 51938
rect 51326 51886 51378 51938
rect 51662 51886 51714 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 16270 51550 16322 51602
rect 22206 51550 22258 51602
rect 22318 51550 22370 51602
rect 23662 51550 23714 51602
rect 31838 51550 31890 51602
rect 33854 51550 33906 51602
rect 34862 51550 34914 51602
rect 35198 51550 35250 51602
rect 35982 51550 36034 51602
rect 38558 51550 38610 51602
rect 49086 51550 49138 51602
rect 4622 51438 4674 51490
rect 7198 51438 7250 51490
rect 11678 51438 11730 51490
rect 12798 51438 12850 51490
rect 13134 51438 13186 51490
rect 13470 51438 13522 51490
rect 15374 51438 15426 51490
rect 15822 51438 15874 51490
rect 17390 51438 17442 51490
rect 18286 51438 18338 51490
rect 19070 51438 19122 51490
rect 23102 51438 23154 51490
rect 34190 51438 34242 51490
rect 35422 51438 35474 51490
rect 37214 51438 37266 51490
rect 38446 51438 38498 51490
rect 38670 51438 38722 51490
rect 6190 51326 6242 51378
rect 6750 51326 6802 51378
rect 10558 51326 10610 51378
rect 11006 51326 11058 51378
rect 11342 51326 11394 51378
rect 12126 51326 12178 51378
rect 13806 51326 13858 51378
rect 14030 51326 14082 51378
rect 14478 51326 14530 51378
rect 15262 51326 15314 51378
rect 15598 51326 15650 51378
rect 16382 51326 16434 51378
rect 16830 51326 16882 51378
rect 18510 51326 18562 51378
rect 19854 51326 19906 51378
rect 20190 51326 20242 51378
rect 20526 51326 20578 51378
rect 22878 51326 22930 51378
rect 28142 51326 28194 51378
rect 28590 51326 28642 51378
rect 33966 51326 34018 51378
rect 34414 51326 34466 51378
rect 34638 51326 34690 51378
rect 34974 51326 35026 51378
rect 38782 51382 38834 51434
rect 40014 51438 40066 51490
rect 42030 51438 42082 51490
rect 42702 51438 42754 51490
rect 42926 51438 42978 51490
rect 43710 51438 43762 51490
rect 47630 51438 47682 51490
rect 49422 51438 49474 51490
rect 52446 51438 52498 51490
rect 35646 51326 35698 51378
rect 36206 51326 36258 51378
rect 36430 51326 36482 51378
rect 36654 51326 36706 51378
rect 36990 51326 37042 51378
rect 39230 51326 39282 51378
rect 39454 51326 39506 51378
rect 39790 51326 39842 51378
rect 41470 51326 41522 51378
rect 42254 51326 42306 51378
rect 43598 51326 43650 51378
rect 46398 51326 46450 51378
rect 46846 51326 46898 51378
rect 47070 51326 47122 51378
rect 47518 51326 47570 51378
rect 48862 51326 48914 51378
rect 49758 51326 49810 51378
rect 49982 51326 50034 51378
rect 50766 51326 50818 51378
rect 51662 51326 51714 51378
rect 6078 51214 6130 51266
rect 16046 51214 16098 51266
rect 17614 51214 17666 51266
rect 20078 51214 20130 51266
rect 22094 51214 22146 51266
rect 23774 51214 23826 51266
rect 25230 51214 25282 51266
rect 27358 51214 27410 51266
rect 29262 51214 29314 51266
rect 31390 51214 31442 51266
rect 36878 51214 36930 51266
rect 39678 51214 39730 51266
rect 41246 51214 41298 51266
rect 45614 51214 45666 51266
rect 46622 51214 46674 51266
rect 49870 51214 49922 51266
rect 50990 51214 51042 51266
rect 51326 51214 51378 51266
rect 54574 51214 54626 51266
rect 10110 51102 10162 51154
rect 10222 51102 10274 51154
rect 10446 51102 10498 51154
rect 11342 51102 11394 51154
rect 11790 51102 11842 51154
rect 12014 51102 12066 51154
rect 13582 51102 13634 51154
rect 14366 51102 14418 51154
rect 16270 51102 16322 51154
rect 17950 51102 18002 51154
rect 18958 51102 19010 51154
rect 23438 51102 23490 51154
rect 35870 51102 35922 51154
rect 41806 51102 41858 51154
rect 43710 51102 43762 51154
rect 45838 51102 45890 51154
rect 46174 51102 46226 51154
rect 47630 51102 47682 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 34638 50766 34690 50818
rect 34974 50766 35026 50818
rect 36206 50766 36258 50818
rect 42702 50766 42754 50818
rect 43038 50766 43090 50818
rect 45054 50766 45106 50818
rect 45390 50766 45442 50818
rect 49870 50766 49922 50818
rect 51102 50766 51154 50818
rect 2494 50654 2546 50706
rect 4622 50654 4674 50706
rect 6638 50654 6690 50706
rect 8766 50654 8818 50706
rect 10894 50654 10946 50706
rect 14702 50654 14754 50706
rect 24334 50654 24386 50706
rect 25006 50654 25058 50706
rect 28366 50654 28418 50706
rect 39230 50654 39282 50706
rect 42254 50654 42306 50706
rect 47070 50654 47122 50706
rect 48190 50654 48242 50706
rect 50206 50654 50258 50706
rect 55582 50654 55634 50706
rect 1822 50542 1874 50594
rect 5966 50542 6018 50594
rect 6190 50542 6242 50594
rect 6862 50542 6914 50594
rect 7086 50542 7138 50594
rect 8094 50542 8146 50594
rect 11230 50542 11282 50594
rect 12574 50542 12626 50594
rect 15038 50542 15090 50594
rect 15374 50542 15426 50594
rect 18398 50542 18450 50594
rect 19070 50542 19122 50594
rect 19406 50542 19458 50594
rect 19742 50542 19794 50594
rect 20190 50542 20242 50594
rect 20414 50542 20466 50594
rect 23550 50542 23602 50594
rect 24110 50542 24162 50594
rect 35422 50542 35474 50594
rect 35646 50542 35698 50594
rect 35982 50542 36034 50594
rect 36990 50542 37042 50594
rect 37662 50542 37714 50594
rect 38222 50542 38274 50594
rect 39118 50542 39170 50594
rect 39902 50542 39954 50594
rect 41694 50542 41746 50594
rect 42366 50542 42418 50594
rect 43598 50542 43650 50594
rect 46062 50542 46114 50594
rect 46622 50542 46674 50594
rect 47518 50542 47570 50594
rect 48078 50542 48130 50594
rect 48302 50542 48354 50594
rect 49310 50542 49362 50594
rect 49646 50542 49698 50594
rect 50542 50542 50594 50594
rect 50878 50542 50930 50594
rect 51214 50542 51266 50594
rect 52670 50542 52722 50594
rect 6526 50430 6578 50482
rect 7534 50430 7586 50482
rect 11790 50430 11842 50482
rect 12350 50430 12402 50482
rect 14926 50430 14978 50482
rect 15822 50430 15874 50482
rect 18510 50430 18562 50482
rect 18734 50430 18786 50482
rect 19182 50430 19234 50482
rect 19966 50430 20018 50482
rect 22542 50430 22594 50482
rect 22878 50430 22930 50482
rect 23886 50430 23938 50482
rect 24558 50430 24610 50482
rect 24894 50430 24946 50482
rect 25454 50430 25506 50482
rect 30718 50430 30770 50482
rect 34750 50430 34802 50482
rect 37102 50430 37154 50482
rect 38334 50430 38386 50482
rect 39006 50430 39058 50482
rect 39342 50430 39394 50482
rect 40126 50430 40178 50482
rect 40686 50430 40738 50482
rect 42030 50430 42082 50482
rect 42926 50430 42978 50482
rect 43374 50430 43426 50482
rect 46174 50430 46226 50482
rect 47294 50430 47346 50482
rect 48526 50430 48578 50482
rect 49422 50430 49474 50482
rect 50094 50430 50146 50482
rect 53454 50430 53506 50482
rect 5070 50318 5122 50370
rect 5630 50318 5682 50370
rect 7422 50318 7474 50370
rect 12910 50318 12962 50370
rect 24446 50318 24498 50370
rect 35310 50318 35362 50370
rect 39566 50318 39618 50370
rect 40014 50318 40066 50370
rect 41358 50318 41410 50370
rect 51326 50318 51378 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 10558 49982 10610 50034
rect 12350 49982 12402 50034
rect 16158 49982 16210 50034
rect 17838 49982 17890 50034
rect 18958 49982 19010 50034
rect 21982 49982 22034 50034
rect 22990 49982 23042 50034
rect 24222 49982 24274 50034
rect 34302 49982 34354 50034
rect 35086 49982 35138 50034
rect 37550 49982 37602 50034
rect 39790 49982 39842 50034
rect 40910 49982 40962 50034
rect 41918 49982 41970 50034
rect 43598 49982 43650 50034
rect 6190 49870 6242 49922
rect 12238 49870 12290 49922
rect 15934 49870 15986 49922
rect 18398 49870 18450 49922
rect 31502 49870 31554 49922
rect 31838 49870 31890 49922
rect 32174 49870 32226 49922
rect 36654 49870 36706 49922
rect 39118 49870 39170 49922
rect 43038 49870 43090 49922
rect 43262 49870 43314 49922
rect 48750 49870 48802 49922
rect 1822 49758 1874 49810
rect 5406 49758 5458 49810
rect 9998 49758 10050 49810
rect 11006 49758 11058 49810
rect 11230 49758 11282 49810
rect 12574 49758 12626 49810
rect 13246 49758 13298 49810
rect 13470 49758 13522 49810
rect 14142 49758 14194 49810
rect 14366 49758 14418 49810
rect 15038 49758 15090 49810
rect 16382 49758 16434 49810
rect 17278 49758 17330 49810
rect 17614 49758 17666 49810
rect 18622 49758 18674 49810
rect 19518 49758 19570 49810
rect 19742 49758 19794 49810
rect 20078 49758 20130 49810
rect 20526 49758 20578 49810
rect 21086 49758 21138 49810
rect 22206 49758 22258 49810
rect 22542 49758 22594 49810
rect 22878 49758 22930 49810
rect 23102 49758 23154 49810
rect 23662 49758 23714 49810
rect 24110 49758 24162 49810
rect 24334 49758 24386 49810
rect 27694 49758 27746 49810
rect 34190 49758 34242 49810
rect 34526 49758 34578 49810
rect 34862 49758 34914 49810
rect 35534 49758 35586 49810
rect 36206 49758 36258 49810
rect 36878 49758 36930 49810
rect 37326 49758 37378 49810
rect 37886 49758 37938 49810
rect 38670 49758 38722 49810
rect 39230 49758 39282 49810
rect 40014 49758 40066 49810
rect 41246 49758 41298 49810
rect 42142 49758 42194 49810
rect 43934 49758 43986 49810
rect 45390 49758 45442 49810
rect 48974 49758 49026 49810
rect 49870 49758 49922 49810
rect 2494 49646 2546 49698
rect 4622 49646 4674 49698
rect 5070 49646 5122 49698
rect 8318 49646 8370 49698
rect 8766 49646 8818 49698
rect 11678 49646 11730 49698
rect 13806 49646 13858 49698
rect 17726 49646 17778 49698
rect 19630 49646 19682 49698
rect 22990 49646 23042 49698
rect 28366 49646 28418 49698
rect 30494 49646 30546 49698
rect 31278 49646 31330 49698
rect 33966 49646 34018 49698
rect 34750 49646 34802 49698
rect 42926 49646 42978 49698
rect 44494 49646 44546 49698
rect 44942 49646 44994 49698
rect 47630 49646 47682 49698
rect 49086 49646 49138 49698
rect 49982 49646 50034 49698
rect 50990 49646 51042 49698
rect 10222 49534 10274 49586
rect 10894 49534 10946 49586
rect 14590 49534 14642 49586
rect 14814 49534 14866 49586
rect 15486 49534 15538 49586
rect 15822 49534 15874 49586
rect 20750 49534 20802 49586
rect 21198 49534 21250 49586
rect 21310 49534 21362 49586
rect 21870 49534 21922 49586
rect 30942 49534 30994 49586
rect 35758 49534 35810 49586
rect 38670 49534 38722 49586
rect 39678 49534 39730 49586
rect 41806 49534 41858 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 4174 49198 4226 49250
rect 4958 49198 5010 49250
rect 6862 49198 6914 49250
rect 7086 49198 7138 49250
rect 21870 49198 21922 49250
rect 22654 49198 22706 49250
rect 36094 49198 36146 49250
rect 39006 49198 39058 49250
rect 43038 49198 43090 49250
rect 49086 49198 49138 49250
rect 50542 49198 50594 49250
rect 7758 49086 7810 49138
rect 16718 49086 16770 49138
rect 19966 49086 20018 49138
rect 23998 49086 24050 49138
rect 28142 49086 28194 49138
rect 29598 49086 29650 49138
rect 34078 49086 34130 49138
rect 37550 49086 37602 49138
rect 40238 49086 40290 49138
rect 44830 49086 44882 49138
rect 4062 48974 4114 49026
rect 4510 48974 4562 49026
rect 4734 48974 4786 49026
rect 5854 48974 5906 49026
rect 6078 48974 6130 49026
rect 7198 48974 7250 49026
rect 9774 48974 9826 49026
rect 9998 48974 10050 49026
rect 10222 48974 10274 49026
rect 13470 48974 13522 49026
rect 16606 48974 16658 49026
rect 17166 48974 17218 49026
rect 21310 48974 21362 49026
rect 21534 48974 21586 49026
rect 22990 48974 23042 49026
rect 24110 48974 24162 49026
rect 27806 48974 27858 49026
rect 28590 48974 28642 49026
rect 29150 48974 29202 49026
rect 29486 48974 29538 49026
rect 30718 48974 30770 49026
rect 31278 48974 31330 49026
rect 34302 48974 34354 49026
rect 36206 48974 36258 49026
rect 37102 48974 37154 49026
rect 37438 48974 37490 49026
rect 38334 48974 38386 49026
rect 39118 48974 39170 49026
rect 39790 48974 39842 49026
rect 40686 48974 40738 49026
rect 41358 48974 41410 49026
rect 41694 48974 41746 49026
rect 42030 48974 42082 49026
rect 42366 48974 42418 49026
rect 43374 48974 43426 49026
rect 44046 48974 44098 49026
rect 47630 48974 47682 49026
rect 49982 48974 50034 49026
rect 50654 48974 50706 49026
rect 50878 48974 50930 49026
rect 3950 48862 4002 48914
rect 6750 48862 6802 48914
rect 7646 48862 7698 48914
rect 9662 48862 9714 48914
rect 14142 48862 14194 48914
rect 15150 48862 15202 48914
rect 17838 48862 17890 48914
rect 20302 48862 20354 48914
rect 20638 48862 20690 48914
rect 23214 48862 23266 48914
rect 23662 48862 23714 48914
rect 23886 48862 23938 48914
rect 27470 48862 27522 48914
rect 27582 48862 27634 48914
rect 30382 48862 30434 48914
rect 31950 48862 32002 48914
rect 34750 48862 34802 48914
rect 34974 48862 35026 48914
rect 37662 48862 37714 48914
rect 39454 48862 39506 48914
rect 41582 48862 41634 48914
rect 42142 48862 42194 48914
rect 44158 48862 44210 48914
rect 46958 48862 47010 48914
rect 49310 48862 49362 48914
rect 49758 48862 49810 48914
rect 50990 48862 51042 48914
rect 4622 48750 4674 48802
rect 6414 48750 6466 48802
rect 7870 48750 7922 48802
rect 8430 48750 8482 48802
rect 11006 48750 11058 48802
rect 11342 48750 11394 48802
rect 22766 48750 22818 48802
rect 25342 48750 25394 48802
rect 25678 48750 25730 48802
rect 26798 48750 26850 48802
rect 27246 48750 27298 48802
rect 28030 48750 28082 48802
rect 28254 48750 28306 48802
rect 29710 48750 29762 48802
rect 34638 48750 34690 48802
rect 35422 48750 35474 48802
rect 36094 48750 36146 48802
rect 37998 48750 38050 48802
rect 48750 48750 48802 48802
rect 51438 48750 51490 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 4286 48414 4338 48466
rect 10334 48414 10386 48466
rect 17502 48414 17554 48466
rect 18398 48414 18450 48466
rect 19406 48414 19458 48466
rect 19854 48414 19906 48466
rect 20078 48414 20130 48466
rect 20526 48414 20578 48466
rect 20974 48414 21026 48466
rect 23326 48414 23378 48466
rect 23998 48414 24050 48466
rect 27582 48414 27634 48466
rect 27694 48414 27746 48466
rect 28814 48414 28866 48466
rect 6750 48302 6802 48354
rect 7870 48302 7922 48354
rect 12126 48302 12178 48354
rect 14142 48302 14194 48354
rect 15598 48302 15650 48354
rect 17726 48302 17778 48354
rect 18622 48302 18674 48354
rect 20414 48302 20466 48354
rect 23774 48302 23826 48354
rect 24670 48302 24722 48354
rect 26686 48302 26738 48354
rect 30718 48302 30770 48354
rect 43262 48302 43314 48354
rect 44046 48302 44098 48354
rect 44494 48302 44546 48354
rect 46958 48302 47010 48354
rect 50094 48302 50146 48354
rect 51214 48302 51266 48354
rect 2830 48190 2882 48242
rect 3054 48190 3106 48242
rect 4062 48190 4114 48242
rect 7534 48190 7586 48242
rect 8094 48190 8146 48242
rect 8654 48190 8706 48242
rect 9774 48190 9826 48242
rect 11342 48190 11394 48242
rect 14702 48190 14754 48242
rect 16830 48190 16882 48242
rect 17278 48190 17330 48242
rect 17950 48190 18002 48242
rect 19182 48190 19234 48242
rect 19742 48190 19794 48242
rect 23662 48190 23714 48242
rect 24334 48190 24386 48242
rect 25790 48190 25842 48242
rect 26014 48190 26066 48242
rect 26462 48190 26514 48242
rect 27358 48190 27410 48242
rect 27806 48190 27858 48242
rect 27918 48190 27970 48242
rect 28702 48190 28754 48242
rect 28926 48190 28978 48242
rect 29374 48190 29426 48242
rect 32510 48190 32562 48242
rect 33294 48190 33346 48242
rect 36206 48190 36258 48242
rect 43374 48190 43426 48242
rect 43822 48190 43874 48242
rect 44606 48190 44658 48242
rect 45390 48190 45442 48242
rect 48638 48190 48690 48242
rect 48974 48190 49026 48242
rect 49198 48190 49250 48242
rect 49758 48190 49810 48242
rect 50542 48190 50594 48242
rect 4622 48078 4674 48130
rect 8766 48078 8818 48130
rect 11678 48078 11730 48130
rect 14814 48078 14866 48130
rect 18398 48078 18450 48130
rect 21422 48078 21474 48130
rect 22766 48078 22818 48130
rect 29150 48078 29202 48130
rect 34302 48078 34354 48130
rect 48190 48078 48242 48130
rect 48862 48078 48914 48130
rect 53342 48078 53394 48130
rect 2718 47966 2770 48018
rect 8990 47966 9042 48018
rect 9998 47966 10050 48018
rect 12350 47966 12402 48018
rect 12686 47966 12738 48018
rect 22990 47966 23042 48018
rect 24334 47966 24386 48018
rect 25454 47966 25506 48018
rect 29598 47966 29650 48018
rect 43262 47966 43314 48018
rect 44718 47966 44770 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 13582 47630 13634 47682
rect 25678 47630 25730 47682
rect 33070 47630 33122 47682
rect 45166 47630 45218 47682
rect 46398 47630 46450 47682
rect 50206 47630 50258 47682
rect 2494 47518 2546 47570
rect 4622 47518 4674 47570
rect 8878 47518 8930 47570
rect 11006 47518 11058 47570
rect 12910 47518 12962 47570
rect 18958 47518 19010 47570
rect 25118 47518 25170 47570
rect 27246 47518 27298 47570
rect 29374 47518 29426 47570
rect 29710 47518 29762 47570
rect 31054 47518 31106 47570
rect 31838 47518 31890 47570
rect 36430 47518 36482 47570
rect 44270 47518 44322 47570
rect 47966 47518 48018 47570
rect 49646 47518 49698 47570
rect 51326 47518 51378 47570
rect 1822 47406 1874 47458
rect 5966 47406 6018 47458
rect 7086 47406 7138 47458
rect 8094 47406 8146 47458
rect 13470 47406 13522 47458
rect 14030 47406 14082 47458
rect 17838 47406 17890 47458
rect 18510 47406 18562 47458
rect 19630 47406 19682 47458
rect 20526 47406 20578 47458
rect 21310 47406 21362 47458
rect 22766 47406 22818 47458
rect 23102 47406 23154 47458
rect 25678 47406 25730 47458
rect 27694 47406 27746 47458
rect 27918 47406 27970 47458
rect 28478 47406 28530 47458
rect 29038 47406 29090 47458
rect 29822 47406 29874 47458
rect 30830 47406 30882 47458
rect 31166 47406 31218 47458
rect 32174 47406 32226 47458
rect 32734 47406 32786 47458
rect 33182 47406 33234 47458
rect 33518 47406 33570 47458
rect 41470 47406 41522 47458
rect 44942 47406 44994 47458
rect 45390 47406 45442 47458
rect 45838 47406 45890 47458
rect 46062 47406 46114 47458
rect 46510 47406 46562 47458
rect 47294 47406 47346 47458
rect 47630 47406 47682 47458
rect 48302 47406 48354 47458
rect 48526 47406 48578 47458
rect 48750 47406 48802 47458
rect 49870 47406 49922 47458
rect 50654 47406 50706 47458
rect 51214 47406 51266 47458
rect 51550 47406 51602 47458
rect 6078 47294 6130 47346
rect 7534 47294 7586 47346
rect 14142 47294 14194 47346
rect 17166 47294 17218 47346
rect 19406 47294 19458 47346
rect 22542 47294 22594 47346
rect 25342 47294 25394 47346
rect 27582 47294 27634 47346
rect 28366 47294 28418 47346
rect 31390 47294 31442 47346
rect 34302 47294 34354 47346
rect 42142 47294 42194 47346
rect 44830 47294 44882 47346
rect 49086 47294 49138 47346
rect 5070 47182 5122 47234
rect 6974 47182 7026 47234
rect 12798 47182 12850 47234
rect 13582 47182 13634 47234
rect 15598 47182 15650 47234
rect 20750 47182 20802 47234
rect 21422 47182 21474 47234
rect 21646 47182 21698 47234
rect 22766 47182 22818 47234
rect 24110 47182 24162 47234
rect 24558 47182 24610 47234
rect 26238 47182 26290 47234
rect 26574 47182 26626 47234
rect 28142 47182 28194 47234
rect 37102 47182 37154 47234
rect 46622 47182 46674 47234
rect 48638 47182 48690 47234
rect 50878 47182 50930 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 15710 46846 15762 46898
rect 16382 46846 16434 46898
rect 19294 46846 19346 46898
rect 19742 46846 19794 46898
rect 20750 46846 20802 46898
rect 24110 46846 24162 46898
rect 27358 46846 27410 46898
rect 28814 46846 28866 46898
rect 28926 46846 28978 46898
rect 29710 46846 29762 46898
rect 30158 46846 30210 46898
rect 33070 46846 33122 46898
rect 35758 46846 35810 46898
rect 51102 46846 51154 46898
rect 2494 46734 2546 46786
rect 3950 46734 4002 46786
rect 6414 46734 6466 46786
rect 12126 46734 12178 46786
rect 13358 46734 13410 46786
rect 13918 46734 13970 46786
rect 15486 46734 15538 46786
rect 16270 46734 16322 46786
rect 22878 46734 22930 46786
rect 23102 46734 23154 46786
rect 26686 46734 26738 46786
rect 28142 46734 28194 46786
rect 28478 46734 28530 46786
rect 28590 46734 28642 46786
rect 29150 46734 29202 46786
rect 29262 46734 29314 46786
rect 29822 46734 29874 46786
rect 30494 46734 30546 46786
rect 30942 46734 30994 46786
rect 31166 46734 31218 46786
rect 32062 46734 32114 46786
rect 32398 46734 32450 46786
rect 34414 46734 34466 46786
rect 34638 46734 34690 46786
rect 47182 46734 47234 46786
rect 3166 46622 3218 46674
rect 3390 46622 3442 46674
rect 3726 46622 3778 46674
rect 4062 46622 4114 46674
rect 11006 46622 11058 46674
rect 11230 46622 11282 46674
rect 11566 46622 11618 46674
rect 12014 46622 12066 46674
rect 12798 46622 12850 46674
rect 13134 46622 13186 46674
rect 13694 46622 13746 46674
rect 14366 46622 14418 46674
rect 15150 46622 15202 46674
rect 16046 46622 16098 46674
rect 17726 46622 17778 46674
rect 17950 46622 18002 46674
rect 18622 46622 18674 46674
rect 19518 46622 19570 46674
rect 20414 46622 20466 46674
rect 21310 46622 21362 46674
rect 21758 46622 21810 46674
rect 22094 46622 22146 46674
rect 22318 46622 22370 46674
rect 23438 46622 23490 46674
rect 25342 46622 25394 46674
rect 25678 46622 25730 46674
rect 27134 46622 27186 46674
rect 28030 46622 28082 46674
rect 30830 46622 30882 46674
rect 31278 46622 31330 46674
rect 31726 46622 31778 46674
rect 33294 46622 33346 46674
rect 33966 46622 34018 46674
rect 36318 46622 36370 46674
rect 39678 46622 39730 46674
rect 40014 46622 40066 46674
rect 41022 46622 41074 46674
rect 44494 46622 44546 46674
rect 44718 46622 44770 46674
rect 45838 46622 45890 46674
rect 46062 46622 46114 46674
rect 47070 46622 47122 46674
rect 47406 46622 47458 46674
rect 49310 46622 49362 46674
rect 49758 46622 49810 46674
rect 50094 46622 50146 46674
rect 50318 46622 50370 46674
rect 50542 46622 50594 46674
rect 7758 46510 7810 46562
rect 10558 46510 10610 46562
rect 18734 46510 18786 46562
rect 19406 46510 19458 46562
rect 20190 46510 20242 46562
rect 24670 46510 24722 46562
rect 26238 46510 26290 46562
rect 34302 46510 34354 46562
rect 35422 46510 35474 46562
rect 37102 46510 37154 46562
rect 39230 46510 39282 46562
rect 40238 46510 40290 46562
rect 41694 46510 41746 46562
rect 43822 46510 43874 46562
rect 46174 46510 46226 46562
rect 46622 46510 46674 46562
rect 48862 46510 48914 46562
rect 6302 46398 6354 46450
rect 6638 46398 6690 46450
rect 10670 46398 10722 46450
rect 11454 46398 11506 46450
rect 14030 46398 14082 46450
rect 15822 46398 15874 46450
rect 16382 46398 16434 46450
rect 17390 46398 17442 46450
rect 26798 46398 26850 46450
rect 27470 46398 27522 46450
rect 29710 46398 29762 46450
rect 32510 46398 32562 46450
rect 35422 46398 35474 46450
rect 35982 46398 36034 46450
rect 40350 46398 40402 46450
rect 45054 46398 45106 46450
rect 45726 46398 45778 46450
rect 50654 46398 50706 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 6414 46062 6466 46114
rect 14926 46062 14978 46114
rect 17166 46062 17218 46114
rect 23438 46062 23490 46114
rect 23662 46062 23714 46114
rect 31390 46062 31442 46114
rect 43822 46062 43874 46114
rect 44382 46062 44434 46114
rect 51550 46062 51602 46114
rect 4622 45950 4674 46002
rect 10894 45950 10946 46002
rect 11790 45950 11842 46002
rect 13694 45950 13746 46002
rect 14590 45950 14642 46002
rect 15038 45950 15090 46002
rect 19854 45950 19906 46002
rect 21758 45950 21810 46002
rect 24222 45950 24274 46002
rect 29486 45950 29538 46002
rect 31838 45950 31890 46002
rect 32958 45950 33010 46002
rect 39566 45950 39618 46002
rect 40238 45950 40290 46002
rect 47294 45950 47346 46002
rect 49422 45950 49474 46002
rect 1822 45838 1874 45890
rect 5630 45838 5682 45890
rect 6190 45838 6242 45890
rect 7086 45838 7138 45890
rect 7982 45838 8034 45890
rect 12574 45838 12626 45890
rect 14142 45838 14194 45890
rect 17726 45838 17778 45890
rect 18846 45838 18898 45890
rect 20638 45838 20690 45890
rect 21310 45838 21362 45890
rect 21534 45838 21586 45890
rect 22542 45838 22594 45890
rect 22990 45838 23042 45890
rect 23886 45838 23938 45890
rect 25006 45838 25058 45890
rect 25342 45838 25394 45890
rect 26798 45838 26850 45890
rect 27582 45838 27634 45890
rect 28030 45838 28082 45890
rect 29374 45838 29426 45890
rect 29598 45838 29650 45890
rect 30046 45838 30098 45890
rect 31054 45838 31106 45890
rect 32062 45838 32114 45890
rect 32510 45838 32562 45890
rect 39230 45838 39282 45890
rect 39902 45838 39954 45890
rect 40462 45838 40514 45890
rect 40910 45838 40962 45890
rect 44046 45838 44098 45890
rect 44942 45838 44994 45890
rect 45838 45838 45890 45890
rect 46622 45838 46674 45890
rect 2494 45726 2546 45778
rect 5854 45726 5906 45778
rect 8766 45726 8818 45778
rect 12910 45726 12962 45778
rect 15710 45726 15762 45778
rect 15822 45726 15874 45778
rect 17054 45726 17106 45778
rect 18286 45726 18338 45778
rect 20302 45726 20354 45778
rect 25902 45726 25954 45778
rect 28254 45726 28306 45778
rect 29150 45726 29202 45778
rect 30158 45726 30210 45778
rect 30718 45726 30770 45778
rect 31726 45726 31778 45778
rect 45614 45726 45666 45778
rect 51662 45726 51714 45778
rect 5070 45614 5122 45666
rect 7646 45614 7698 45666
rect 16046 45614 16098 45666
rect 17166 45614 17218 45666
rect 17950 45614 18002 45666
rect 19406 45614 19458 45666
rect 22206 45614 22258 45666
rect 24110 45614 24162 45666
rect 24334 45614 24386 45666
rect 25566 45614 25618 45666
rect 25678 45614 25730 45666
rect 26014 45614 26066 45666
rect 26238 45614 26290 45666
rect 26910 45614 26962 45666
rect 27022 45614 27074 45666
rect 27246 45614 27298 45666
rect 27806 45614 27858 45666
rect 31278 45614 31330 45666
rect 49870 45614 49922 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 2606 45278 2658 45330
rect 5630 45278 5682 45330
rect 9998 45278 10050 45330
rect 12350 45278 12402 45330
rect 14478 45278 14530 45330
rect 14702 45278 14754 45330
rect 15150 45278 15202 45330
rect 16830 45278 16882 45330
rect 25678 45278 25730 45330
rect 39678 45278 39730 45330
rect 44494 45278 44546 45330
rect 2494 45166 2546 45218
rect 4510 45166 4562 45218
rect 5966 45166 6018 45218
rect 8654 45166 8706 45218
rect 8990 45166 9042 45218
rect 15374 45166 15426 45218
rect 17726 45166 17778 45218
rect 18398 45166 18450 45218
rect 25902 45166 25954 45218
rect 27918 45166 27970 45218
rect 31390 45166 31442 45218
rect 32286 45166 32338 45218
rect 32510 45166 32562 45218
rect 38558 45166 38610 45218
rect 39566 45166 39618 45218
rect 40238 45166 40290 45218
rect 40350 45166 40402 45218
rect 41470 45166 41522 45218
rect 42366 45166 42418 45218
rect 50206 45166 50258 45218
rect 2718 45054 2770 45106
rect 3166 45054 3218 45106
rect 4958 45054 5010 45106
rect 5406 45054 5458 45106
rect 10670 45054 10722 45106
rect 11006 45054 11058 45106
rect 12014 45054 12066 45106
rect 14366 45054 14418 45106
rect 15486 45054 15538 45106
rect 18062 45054 18114 45106
rect 18622 45054 18674 45106
rect 18958 45054 19010 45106
rect 20638 45054 20690 45106
rect 21534 45054 21586 45106
rect 23214 45054 23266 45106
rect 23886 45054 23938 45106
rect 26686 45054 26738 45106
rect 27246 45054 27298 45106
rect 27470 45054 27522 45106
rect 28926 45054 28978 45106
rect 30046 45054 30098 45106
rect 30718 45054 30770 45106
rect 31278 45054 31330 45106
rect 33742 45054 33794 45106
rect 33966 45054 34018 45106
rect 34414 45054 34466 45106
rect 34750 45054 34802 45106
rect 38334 45054 38386 45106
rect 41022 45054 41074 45106
rect 41582 45054 41634 45106
rect 41694 45054 41746 45106
rect 41918 45054 41970 45106
rect 42478 45054 42530 45106
rect 49422 45054 49474 45106
rect 10558 44942 10610 44994
rect 11790 44942 11842 44994
rect 15934 44942 15986 44994
rect 16718 44942 16770 44994
rect 20302 44942 20354 44994
rect 23550 44942 23602 44994
rect 26350 44942 26402 44994
rect 28702 44942 28754 44994
rect 29262 44942 29314 44994
rect 29598 44942 29650 44994
rect 31390 44942 31442 44994
rect 33406 44942 33458 44994
rect 34190 44942 34242 44994
rect 35422 44942 35474 44994
rect 37550 44942 37602 44994
rect 40798 44942 40850 44994
rect 41022 44942 41074 44994
rect 42142 44942 42194 44994
rect 49086 44942 49138 44994
rect 52334 44942 52386 44994
rect 17950 44830 18002 44882
rect 18286 44830 18338 44882
rect 32174 44830 32226 44882
rect 39678 44830 39730 44882
rect 40238 44830 40290 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 3614 44494 3666 44546
rect 4174 44494 4226 44546
rect 10110 44494 10162 44546
rect 10446 44494 10498 44546
rect 15486 44494 15538 44546
rect 16494 44494 16546 44546
rect 17502 44494 17554 44546
rect 29150 44494 29202 44546
rect 29374 44494 29426 44546
rect 32510 44494 32562 44546
rect 34638 44494 34690 44546
rect 2494 44382 2546 44434
rect 8542 44382 8594 44434
rect 10222 44382 10274 44434
rect 11790 44382 11842 44434
rect 16606 44382 16658 44434
rect 17054 44382 17106 44434
rect 25006 44382 25058 44434
rect 25790 44382 25842 44434
rect 30942 44382 30994 44434
rect 32846 44382 32898 44434
rect 34078 44382 34130 44434
rect 37774 44382 37826 44434
rect 39342 44382 39394 44434
rect 40126 44382 40178 44434
rect 40798 44382 40850 44434
rect 41918 44382 41970 44434
rect 44830 44382 44882 44434
rect 2270 44270 2322 44322
rect 2718 44270 2770 44322
rect 2830 44270 2882 44322
rect 3390 44270 3442 44322
rect 3726 44270 3778 44322
rect 4510 44270 4562 44322
rect 4958 44270 5010 44322
rect 5630 44270 5682 44322
rect 10670 44270 10722 44322
rect 11118 44270 11170 44322
rect 11454 44270 11506 44322
rect 12574 44270 12626 44322
rect 13582 44270 13634 44322
rect 13694 44270 13746 44322
rect 14030 44270 14082 44322
rect 14254 44270 14306 44322
rect 14478 44270 14530 44322
rect 15038 44270 15090 44322
rect 17278 44270 17330 44322
rect 17950 44270 18002 44322
rect 18286 44270 18338 44322
rect 18622 44270 18674 44322
rect 19406 44270 19458 44322
rect 19854 44270 19906 44322
rect 22318 44270 22370 44322
rect 23326 44270 23378 44322
rect 25678 44270 25730 44322
rect 26462 44270 26514 44322
rect 27358 44270 27410 44322
rect 28254 44270 28306 44322
rect 28590 44270 28642 44322
rect 29598 44270 29650 44322
rect 29822 44270 29874 44322
rect 30046 44270 30098 44322
rect 30382 44270 30434 44322
rect 31278 44270 31330 44322
rect 31614 44270 31666 44322
rect 31950 44270 32002 44322
rect 33518 44270 33570 44322
rect 33742 44270 33794 44322
rect 38782 44270 38834 44322
rect 39790 44270 39842 44322
rect 41246 44270 41298 44322
rect 47742 44270 47794 44322
rect 3278 44158 3330 44210
rect 6414 44158 6466 44210
rect 11230 44158 11282 44210
rect 12238 44158 12290 44210
rect 14926 44158 14978 44210
rect 15486 44158 15538 44210
rect 15934 44158 15986 44210
rect 17726 44158 17778 44210
rect 19294 44158 19346 44210
rect 22206 44158 22258 44210
rect 23214 44158 23266 44210
rect 26014 44158 26066 44210
rect 26686 44158 26738 44210
rect 28478 44158 28530 44210
rect 33966 44158 34018 44210
rect 34526 44158 34578 44210
rect 38446 44158 38498 44210
rect 46958 44158 47010 44210
rect 4286 44046 4338 44098
rect 5070 44046 5122 44098
rect 9102 44046 9154 44098
rect 9550 44046 9602 44098
rect 12350 44046 12402 44098
rect 13806 44046 13858 44098
rect 14702 44046 14754 44098
rect 16494 44046 16546 44098
rect 20190 44046 20242 44098
rect 29934 44046 29986 44098
rect 30830 44046 30882 44098
rect 31054 44046 31106 44098
rect 31614 44046 31666 44098
rect 32734 44046 32786 44098
rect 34078 44046 34130 44098
rect 34638 44046 34690 44098
rect 44158 44046 44210 44098
rect 48190 44046 48242 44098
rect 50878 44046 50930 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 5070 43710 5122 43762
rect 5854 43710 5906 43762
rect 12910 43710 12962 43762
rect 19294 43710 19346 43762
rect 22430 43710 22482 43762
rect 23662 43710 23714 43762
rect 26798 43710 26850 43762
rect 39790 43710 39842 43762
rect 41358 43710 41410 43762
rect 46174 43710 46226 43762
rect 2494 43598 2546 43650
rect 4958 43598 5010 43650
rect 10222 43598 10274 43650
rect 10334 43598 10386 43650
rect 10894 43598 10946 43650
rect 11118 43598 11170 43650
rect 11230 43598 11282 43650
rect 12798 43598 12850 43650
rect 13806 43598 13858 43650
rect 15374 43598 15426 43650
rect 16382 43598 16434 43650
rect 17726 43598 17778 43650
rect 18846 43598 18898 43650
rect 20638 43598 20690 43650
rect 24222 43598 24274 43650
rect 24670 43598 24722 43650
rect 25342 43598 25394 43650
rect 27022 43598 27074 43650
rect 29598 43598 29650 43650
rect 33406 43598 33458 43650
rect 34414 43598 34466 43650
rect 34638 43598 34690 43650
rect 38558 43598 38610 43650
rect 39118 43598 39170 43650
rect 39230 43598 39282 43650
rect 39566 43598 39618 43650
rect 40350 43598 40402 43650
rect 41918 43598 41970 43650
rect 42366 43598 42418 43650
rect 46846 43598 46898 43650
rect 50094 43598 50146 43650
rect 50430 43598 50482 43650
rect 1822 43486 1874 43538
rect 5518 43486 5570 43538
rect 5742 43486 5794 43538
rect 6638 43486 6690 43538
rect 11454 43486 11506 43538
rect 11790 43486 11842 43538
rect 12014 43486 12066 43538
rect 12238 43486 12290 43538
rect 12686 43486 12738 43538
rect 13134 43486 13186 43538
rect 13358 43486 13410 43538
rect 13694 43486 13746 43538
rect 13918 43486 13970 43538
rect 14366 43486 14418 43538
rect 15150 43486 15202 43538
rect 16270 43486 16322 43538
rect 16606 43486 16658 43538
rect 16942 43486 16994 43538
rect 18174 43486 18226 43538
rect 18398 43486 18450 43538
rect 19518 43486 19570 43538
rect 21534 43486 21586 43538
rect 21870 43486 21922 43538
rect 23214 43486 23266 43538
rect 23550 43486 23602 43538
rect 23774 43486 23826 43538
rect 24446 43486 24498 43538
rect 25678 43486 25730 43538
rect 26126 43486 26178 43538
rect 26462 43486 26514 43538
rect 27358 43486 27410 43538
rect 27806 43486 27858 43538
rect 28254 43486 28306 43538
rect 28478 43486 28530 43538
rect 28702 43486 28754 43538
rect 28926 43486 28978 43538
rect 29710 43486 29762 43538
rect 30382 43486 30434 43538
rect 31054 43486 31106 43538
rect 31166 43486 31218 43538
rect 33070 43486 33122 43538
rect 35086 43486 35138 43538
rect 38446 43486 38498 43538
rect 38782 43486 38834 43538
rect 38894 43486 38946 43538
rect 40798 43486 40850 43538
rect 41246 43486 41298 43538
rect 41470 43486 41522 43538
rect 42142 43486 42194 43538
rect 44830 43486 44882 43538
rect 45278 43486 45330 43538
rect 49086 43486 49138 43538
rect 49646 43486 49698 43538
rect 4622 43374 4674 43426
rect 7422 43374 7474 43426
rect 9886 43374 9938 43426
rect 14814 43374 14866 43426
rect 16158 43374 16210 43426
rect 17502 43374 17554 43426
rect 24558 43374 24610 43426
rect 27134 43374 27186 43426
rect 30494 43374 30546 43426
rect 34750 43374 34802 43426
rect 35870 43374 35922 43426
rect 37998 43374 38050 43426
rect 39902 43374 39954 43426
rect 42254 43374 42306 43426
rect 45390 43374 45442 43426
rect 46174 43374 46226 43426
rect 47294 43374 47346 43426
rect 49758 43374 49810 43426
rect 51102 43374 51154 43426
rect 5854 43262 5906 43314
rect 10222 43262 10274 43314
rect 11678 43262 11730 43314
rect 18622 43262 18674 43314
rect 19182 43262 19234 43314
rect 28814 43262 28866 43314
rect 45838 43262 45890 43314
rect 46062 43262 46114 43314
rect 51326 43262 51378 43314
rect 51662 43262 51714 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 3390 42926 3442 42978
rect 3726 42926 3778 42978
rect 7198 42926 7250 42978
rect 7534 42926 7586 42978
rect 11678 42926 11730 42978
rect 12910 42926 12962 42978
rect 16046 42926 16098 42978
rect 18846 42926 18898 42978
rect 22654 42926 22706 42978
rect 30046 42926 30098 42978
rect 34526 42926 34578 42978
rect 45278 42926 45330 42978
rect 45838 42926 45890 42978
rect 3950 42814 4002 42866
rect 4734 42814 4786 42866
rect 6526 42814 6578 42866
rect 8654 42814 8706 42866
rect 10782 42814 10834 42866
rect 11454 42814 11506 42866
rect 14702 42814 14754 42866
rect 15822 42814 15874 42866
rect 17054 42814 17106 42866
rect 20526 42814 20578 42866
rect 23550 42814 23602 42866
rect 25566 42814 25618 42866
rect 26350 42814 26402 42866
rect 27582 42814 27634 42866
rect 29150 42814 29202 42866
rect 29486 42814 29538 42866
rect 30942 42814 30994 42866
rect 36094 42814 36146 42866
rect 39902 42814 39954 42866
rect 42142 42814 42194 42866
rect 45838 42814 45890 42866
rect 50206 42814 50258 42866
rect 5854 42702 5906 42754
rect 6638 42702 6690 42754
rect 6974 42702 7026 42754
rect 7870 42702 7922 42754
rect 12798 42702 12850 42754
rect 13358 42702 13410 42754
rect 13694 42702 13746 42754
rect 13918 42702 13970 42754
rect 14142 42702 14194 42754
rect 15598 42702 15650 42754
rect 16270 42702 16322 42754
rect 16942 42702 16994 42754
rect 17726 42702 17778 42754
rect 19406 42702 19458 42754
rect 19854 42702 19906 42754
rect 22318 42702 22370 42754
rect 22990 42702 23042 42754
rect 24894 42702 24946 42754
rect 25454 42702 25506 42754
rect 26462 42702 26514 42754
rect 26798 42702 26850 42754
rect 28254 42702 28306 42754
rect 28590 42702 28642 42754
rect 29934 42702 29986 42754
rect 30606 42702 30658 42754
rect 30830 42702 30882 42754
rect 34750 42702 34802 42754
rect 36990 42702 37042 42754
rect 40350 42702 40402 42754
rect 41134 42702 41186 42754
rect 41694 42702 41746 42754
rect 42366 42702 42418 42754
rect 46286 42702 46338 42754
rect 46846 42702 46898 42754
rect 47406 42702 47458 42754
rect 50542 42702 50594 42754
rect 50766 42702 50818 42754
rect 5630 42590 5682 42642
rect 6302 42590 6354 42642
rect 14366 42590 14418 42642
rect 14814 42590 14866 42642
rect 15486 42590 15538 42642
rect 17166 42590 17218 42642
rect 17950 42590 18002 42642
rect 18062 42590 18114 42642
rect 18510 42590 18562 42642
rect 18734 42590 18786 42642
rect 22094 42590 22146 42642
rect 23214 42590 23266 42642
rect 26238 42590 26290 42642
rect 27134 42590 27186 42642
rect 28478 42590 28530 42642
rect 37774 42590 37826 42642
rect 41806 42590 41858 42642
rect 46622 42590 46674 42642
rect 48078 42590 48130 42642
rect 51102 42590 51154 42642
rect 51438 42590 51490 42642
rect 51662 42590 51714 42642
rect 51998 42590 52050 42642
rect 5070 42478 5122 42530
rect 12014 42478 12066 42530
rect 12686 42478 12738 42530
rect 13806 42478 13858 42530
rect 17390 42478 17442 42530
rect 19966 42478 20018 42530
rect 26014 42478 26066 42530
rect 28030 42478 28082 42530
rect 29374 42478 29426 42530
rect 30382 42478 30434 42530
rect 31390 42478 31442 42530
rect 32622 42478 32674 42530
rect 34190 42478 34242 42530
rect 34974 42478 35026 42530
rect 35086 42478 35138 42530
rect 35198 42478 35250 42530
rect 35646 42478 35698 42530
rect 42702 42478 42754 42530
rect 45390 42478 45442 42530
rect 51774 42478 51826 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 4398 42142 4450 42194
rect 11118 42142 11170 42194
rect 14366 42142 14418 42194
rect 14478 42030 14530 42082
rect 14926 42030 14978 42082
rect 17838 42030 17890 42082
rect 18510 42030 18562 42082
rect 18622 42086 18674 42138
rect 27470 42142 27522 42194
rect 28366 42142 28418 42194
rect 28590 42142 28642 42194
rect 29710 42142 29762 42194
rect 31278 42142 31330 42194
rect 32286 42142 32338 42194
rect 36654 42142 36706 42194
rect 37102 42142 37154 42194
rect 19294 42030 19346 42082
rect 19742 42030 19794 42082
rect 19966 42030 20018 42082
rect 22878 42030 22930 42082
rect 27134 42030 27186 42082
rect 27246 42030 27298 42082
rect 30382 42030 30434 42082
rect 32062 42030 32114 42082
rect 33294 42030 33346 42082
rect 35534 42030 35586 42082
rect 36094 42030 36146 42082
rect 53006 42030 53058 42082
rect 53790 42030 53842 42082
rect 2830 41918 2882 41970
rect 3390 41918 3442 41970
rect 3838 41918 3890 41970
rect 4062 41918 4114 41970
rect 4734 41918 4786 41970
rect 4958 41918 5010 41970
rect 5294 41918 5346 41970
rect 8766 41918 8818 41970
rect 11342 41918 11394 41970
rect 12238 41918 12290 41970
rect 15486 41918 15538 41970
rect 16046 41918 16098 41970
rect 16270 41918 16322 41970
rect 16494 41918 16546 41970
rect 16942 41918 16994 41970
rect 17390 41918 17442 41970
rect 17950 41918 18002 41970
rect 18174 41918 18226 41970
rect 20302 41918 20354 41970
rect 20750 41918 20802 41970
rect 21534 41918 21586 41970
rect 21982 41918 22034 41970
rect 22990 41918 23042 41970
rect 23102 41918 23154 41970
rect 25342 41918 25394 41970
rect 26014 41918 26066 41970
rect 26462 41918 26514 41970
rect 27806 41918 27858 41970
rect 28142 41918 28194 41970
rect 28814 41918 28866 41970
rect 29038 41918 29090 41970
rect 29486 41918 29538 41970
rect 30046 41918 30098 41970
rect 30942 41918 30994 41970
rect 31614 41918 31666 41970
rect 34974 41918 35026 41970
rect 35310 41918 35362 41970
rect 35870 41918 35922 41970
rect 38670 41918 38722 41970
rect 38894 41918 38946 41970
rect 39790 41918 39842 41970
rect 40126 41918 40178 41970
rect 42254 41918 42306 41970
rect 43262 41918 43314 41970
rect 44046 41918 44098 41970
rect 45390 41918 45442 41970
rect 49422 41918 49474 41970
rect 49758 41918 49810 41970
rect 51774 41918 51826 41970
rect 52782 41918 52834 41970
rect 53678 41918 53730 41970
rect 3166 41806 3218 41858
rect 3950 41806 4002 41858
rect 5854 41806 5906 41858
rect 7646 41806 7698 41858
rect 9662 41806 9714 41858
rect 13918 41806 13970 41858
rect 16382 41806 16434 41858
rect 19406 41806 19458 41858
rect 19966 41806 20018 41858
rect 27694 41806 27746 41858
rect 29598 41806 29650 41858
rect 31838 41806 31890 41858
rect 32174 41806 32226 41858
rect 33182 41806 33234 41858
rect 35422 41806 35474 41858
rect 36206 41806 36258 41858
rect 38334 41806 38386 41858
rect 45614 41806 45666 41858
rect 48862 41806 48914 41858
rect 50766 41806 50818 41858
rect 51662 41806 51714 41858
rect 53566 41806 53618 41858
rect 2830 41694 2882 41746
rect 5630 41694 5682 41746
rect 14366 41694 14418 41746
rect 14814 41694 14866 41746
rect 18622 41694 18674 41746
rect 19070 41694 19122 41746
rect 20750 41694 20802 41746
rect 21086 41694 21138 41746
rect 23550 41694 23602 41746
rect 26238 41694 26290 41746
rect 28702 41694 28754 41746
rect 33070 41694 33122 41746
rect 39118 41694 39170 41746
rect 39342 41694 39394 41746
rect 39454 41694 39506 41746
rect 39790 41694 39842 41746
rect 46062 41694 46114 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 6414 41358 6466 41410
rect 6862 41358 6914 41410
rect 13470 41358 13522 41410
rect 13582 41358 13634 41410
rect 15262 41358 15314 41410
rect 18286 41358 18338 41410
rect 18622 41358 18674 41410
rect 19966 41358 20018 41410
rect 20302 41358 20354 41410
rect 22542 41358 22594 41410
rect 25342 41358 25394 41410
rect 27582 41358 27634 41410
rect 49982 41358 50034 41410
rect 51774 41358 51826 41410
rect 2494 41246 2546 41298
rect 4622 41246 4674 41298
rect 5070 41246 5122 41298
rect 7758 41246 7810 41298
rect 8878 41246 8930 41298
rect 11006 41246 11058 41298
rect 11902 41246 11954 41298
rect 14254 41246 14306 41298
rect 14478 41246 14530 41298
rect 14814 41246 14866 41298
rect 16158 41246 16210 41298
rect 16606 41246 16658 41298
rect 19630 41246 19682 41298
rect 23326 41246 23378 41298
rect 32734 41246 32786 41298
rect 34862 41246 34914 41298
rect 36206 41246 36258 41298
rect 43038 41246 43090 41298
rect 44830 41246 44882 41298
rect 48862 41246 48914 41298
rect 1822 41134 1874 41186
rect 5966 41134 6018 41186
rect 6190 41134 6242 41186
rect 6974 41134 7026 41186
rect 8094 41134 8146 41186
rect 12238 41134 12290 41186
rect 13694 41134 13746 41186
rect 14030 41134 14082 41186
rect 15038 41134 15090 41186
rect 17390 41134 17442 41186
rect 17726 41134 17778 41186
rect 17950 41134 18002 41186
rect 18286 41134 18338 41186
rect 19742 41134 19794 41186
rect 20190 41134 20242 41186
rect 21422 41134 21474 41186
rect 21982 41134 22034 41186
rect 22206 41134 22258 41186
rect 22654 41134 22706 41186
rect 25454 41134 25506 41186
rect 25790 41134 25842 41186
rect 26238 41134 26290 41186
rect 26798 41134 26850 41186
rect 27134 41134 27186 41186
rect 27694 41134 27746 41186
rect 29934 41134 29986 41186
rect 32062 41134 32114 41186
rect 35310 41134 35362 41186
rect 35758 41134 35810 41186
rect 36990 41134 37042 41186
rect 37550 41134 37602 41186
rect 39566 41134 39618 41186
rect 42030 41134 42082 41186
rect 42814 41134 42866 41186
rect 43822 41134 43874 41186
rect 47742 41134 47794 41186
rect 50990 41134 51042 41186
rect 51214 41134 51266 41186
rect 51326 41134 51378 41186
rect 6526 41022 6578 41074
rect 7086 41022 7138 41074
rect 19182 41022 19234 41074
rect 19294 41022 19346 41074
rect 22430 41022 22482 41074
rect 22990 41022 23042 41074
rect 23438 41022 23490 41074
rect 29486 41022 29538 41074
rect 30606 41022 30658 41074
rect 35422 41022 35474 41074
rect 37214 41022 37266 41074
rect 39678 41022 39730 41074
rect 41582 41022 41634 41074
rect 42478 41022 42530 41074
rect 44270 41022 44322 41074
rect 46958 41022 47010 41074
rect 49982 41022 50034 41074
rect 50094 41022 50146 41074
rect 50430 41022 50482 41074
rect 50542 41022 50594 41074
rect 12574 40910 12626 40962
rect 15598 40910 15650 40962
rect 16046 40910 16098 40962
rect 17054 40910 17106 40962
rect 17614 40910 17666 40962
rect 19070 40910 19122 40962
rect 21646 40910 21698 40962
rect 22878 40910 22930 40962
rect 25342 40910 25394 40962
rect 29150 40910 29202 40962
rect 29262 40910 29314 40962
rect 29374 40910 29426 40962
rect 30270 40910 30322 40962
rect 35646 40910 35698 40962
rect 37102 40910 37154 40962
rect 38110 40910 38162 40962
rect 38894 40910 38946 40962
rect 39230 40910 39282 40962
rect 39902 40910 39954 40962
rect 41470 40910 41522 40962
rect 41694 40910 41746 40962
rect 43710 40910 43762 40962
rect 44158 40910 44210 40962
rect 48190 40910 48242 40962
rect 49422 40910 49474 40962
rect 50766 40910 50818 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 4510 40574 4562 40626
rect 8990 40574 9042 40626
rect 13918 40574 13970 40626
rect 14478 40574 14530 40626
rect 14590 40574 14642 40626
rect 15710 40574 15762 40626
rect 16382 40574 16434 40626
rect 22094 40574 22146 40626
rect 24670 40574 24722 40626
rect 28702 40574 28754 40626
rect 29710 40574 29762 40626
rect 32286 40574 32338 40626
rect 38446 40574 38498 40626
rect 44382 40574 44434 40626
rect 45278 40574 45330 40626
rect 45950 40574 46002 40626
rect 46846 40574 46898 40626
rect 47182 40574 47234 40626
rect 48974 40574 49026 40626
rect 49198 40574 49250 40626
rect 51438 40574 51490 40626
rect 51662 40574 51714 40626
rect 51998 40574 52050 40626
rect 52222 40574 52274 40626
rect 52558 40574 52610 40626
rect 7758 40462 7810 40514
rect 10334 40462 10386 40514
rect 13134 40462 13186 40514
rect 16046 40462 16098 40514
rect 16158 40462 16210 40514
rect 16718 40462 16770 40514
rect 16830 40462 16882 40514
rect 22318 40462 22370 40514
rect 22430 40462 22482 40514
rect 24558 40462 24610 40514
rect 26238 40462 26290 40514
rect 26798 40462 26850 40514
rect 26910 40462 26962 40514
rect 27358 40462 27410 40514
rect 27470 40462 27522 40514
rect 28366 40462 28418 40514
rect 29038 40462 29090 40514
rect 30942 40462 30994 40514
rect 32510 40462 32562 40514
rect 35758 40462 35810 40514
rect 38222 40462 38274 40514
rect 39790 40462 39842 40514
rect 45614 40462 45666 40514
rect 46286 40462 46338 40514
rect 50990 40462 51042 40514
rect 51326 40462 51378 40514
rect 51886 40462 51938 40514
rect 8430 40350 8482 40402
rect 9550 40350 9602 40402
rect 12798 40350 12850 40402
rect 13918 40350 13970 40402
rect 14702 40350 14754 40402
rect 15038 40350 15090 40402
rect 15486 40350 15538 40402
rect 16494 40350 16546 40402
rect 17502 40350 17554 40402
rect 18734 40350 18786 40402
rect 19630 40350 19682 40402
rect 19966 40350 20018 40402
rect 20414 40350 20466 40402
rect 21198 40350 21250 40402
rect 21646 40350 21698 40402
rect 21870 40350 21922 40402
rect 25230 40350 25282 40402
rect 26014 40350 26066 40402
rect 28142 40350 28194 40402
rect 29374 40350 29426 40402
rect 29934 40350 29986 40402
rect 30830 40350 30882 40402
rect 31950 40350 32002 40402
rect 35086 40350 35138 40402
rect 39006 40350 39058 40402
rect 40014 40350 40066 40402
rect 41358 40350 41410 40402
rect 41918 40350 41970 40402
rect 42254 40350 42306 40402
rect 42590 40350 42642 40402
rect 42926 40350 42978 40402
rect 43262 40350 43314 40402
rect 43598 40350 43650 40402
rect 43822 40350 43874 40402
rect 44942 40350 44994 40402
rect 48190 40350 48242 40402
rect 48750 40350 48802 40402
rect 49534 40350 49586 40402
rect 49758 40350 49810 40402
rect 50094 40350 50146 40402
rect 50318 40350 50370 40402
rect 50766 40350 50818 40402
rect 4622 40238 4674 40290
rect 4846 40238 4898 40290
rect 5630 40238 5682 40290
rect 12462 40238 12514 40290
rect 18062 40238 18114 40290
rect 18510 40238 18562 40290
rect 21758 40238 21810 40290
rect 25678 40238 25730 40290
rect 29822 40238 29874 40290
rect 37886 40238 37938 40290
rect 38334 40238 38386 40290
rect 42030 40238 42082 40290
rect 42478 40238 42530 40290
rect 47742 40238 47794 40290
rect 49198 40238 49250 40290
rect 49646 40238 49698 40290
rect 50878 40238 50930 40290
rect 4510 40126 4562 40178
rect 18286 40126 18338 40178
rect 19182 40126 19234 40178
rect 26910 40126 26962 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 6190 39790 6242 39842
rect 15374 39790 15426 39842
rect 15822 39790 15874 39842
rect 26686 39790 26738 39842
rect 27246 39790 27298 39842
rect 28590 39790 28642 39842
rect 29934 39790 29986 39842
rect 5070 39678 5122 39730
rect 8766 39678 8818 39730
rect 11454 39678 11506 39730
rect 12686 39678 12738 39730
rect 16158 39678 16210 39730
rect 18062 39678 18114 39730
rect 20750 39678 20802 39730
rect 23550 39678 23602 39730
rect 25118 39678 25170 39730
rect 30046 39678 30098 39730
rect 36430 39678 36482 39730
rect 37774 39678 37826 39730
rect 39902 39678 39954 39730
rect 41918 39678 41970 39730
rect 42478 39678 42530 39730
rect 48862 39678 48914 39730
rect 4734 39566 4786 39618
rect 5518 39566 5570 39618
rect 12238 39566 12290 39618
rect 12574 39566 12626 39618
rect 15486 39566 15538 39618
rect 17838 39566 17890 39618
rect 19630 39566 19682 39618
rect 21310 39566 21362 39618
rect 21870 39566 21922 39618
rect 22430 39566 22482 39618
rect 25006 39566 25058 39618
rect 25342 39566 25394 39618
rect 25678 39566 25730 39618
rect 26574 39566 26626 39618
rect 27694 39566 27746 39618
rect 27918 39566 27970 39618
rect 28590 39566 28642 39618
rect 29038 39566 29090 39618
rect 32510 39566 32562 39618
rect 33406 39566 33458 39618
rect 37102 39566 37154 39618
rect 41246 39566 41298 39618
rect 41694 39566 41746 39618
rect 42702 39566 42754 39618
rect 44830 39566 44882 39618
rect 45390 39566 45442 39618
rect 46286 39566 46338 39618
rect 47182 39566 47234 39618
rect 47518 39566 47570 39618
rect 47966 39566 48018 39618
rect 48414 39566 48466 39618
rect 48638 39566 48690 39618
rect 49310 39566 49362 39618
rect 49758 39566 49810 39618
rect 49870 39566 49922 39618
rect 50318 39566 50370 39618
rect 50654 39566 50706 39618
rect 13022 39454 13074 39506
rect 14590 39454 14642 39506
rect 14926 39454 14978 39506
rect 17054 39454 17106 39506
rect 18286 39454 18338 39506
rect 26014 39454 26066 39506
rect 28254 39454 28306 39506
rect 29598 39454 29650 39506
rect 32286 39454 32338 39506
rect 32846 39454 32898 39506
rect 33070 39454 33122 39506
rect 44270 39454 44322 39506
rect 45838 39454 45890 39506
rect 46174 39454 46226 39506
rect 46846 39454 46898 39506
rect 46958 39454 47010 39506
rect 49086 39454 49138 39506
rect 49646 39454 49698 39506
rect 51214 39454 51266 39506
rect 51662 39454 51714 39506
rect 4062 39342 4114 39394
rect 4174 39342 4226 39394
rect 4286 39342 4338 39394
rect 5854 39342 5906 39394
rect 6078 39342 6130 39394
rect 6414 39342 6466 39394
rect 6750 39342 6802 39394
rect 15374 39342 15426 39394
rect 16046 39342 16098 39394
rect 20190 39342 20242 39394
rect 22542 39342 22594 39394
rect 22766 39342 22818 39394
rect 23102 39342 23154 39394
rect 23998 39342 24050 39394
rect 26686 39342 26738 39394
rect 29374 39342 29426 39394
rect 29710 39342 29762 39394
rect 30158 39342 30210 39394
rect 31950 39342 32002 39394
rect 32622 39342 32674 39394
rect 33294 39342 33346 39394
rect 43710 39342 43762 39394
rect 45278 39342 45330 39394
rect 45502 39342 45554 39394
rect 46062 39342 46114 39394
rect 50990 39342 51042 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 6190 39006 6242 39058
rect 7646 39006 7698 39058
rect 15150 39006 15202 39058
rect 16270 39006 16322 39058
rect 18846 39006 18898 39058
rect 25230 39006 25282 39058
rect 29038 39006 29090 39058
rect 29262 39006 29314 39058
rect 33742 39006 33794 39058
rect 34190 39006 34242 39058
rect 37662 39006 37714 39058
rect 41582 39006 41634 39058
rect 46958 39006 47010 39058
rect 2494 38894 2546 38946
rect 5182 38894 5234 38946
rect 5294 38894 5346 38946
rect 5854 38894 5906 38946
rect 13806 38894 13858 38946
rect 14478 38894 14530 38946
rect 15374 38894 15426 38946
rect 16158 38894 16210 38946
rect 18398 38894 18450 38946
rect 19742 38894 19794 38946
rect 22542 38894 22594 38946
rect 28926 38894 28978 38946
rect 37438 38894 37490 38946
rect 37998 38894 38050 38946
rect 38558 38894 38610 38946
rect 41918 38894 41970 38946
rect 45502 38894 45554 38946
rect 45950 38894 46002 38946
rect 47742 38894 47794 38946
rect 47854 38894 47906 38946
rect 47966 38894 48018 38946
rect 49758 38894 49810 38946
rect 51214 38894 51266 38946
rect 1822 38782 1874 38834
rect 5406 38782 5458 38834
rect 6526 38782 6578 38834
rect 6974 38782 7026 38834
rect 7422 38782 7474 38834
rect 14590 38782 14642 38834
rect 14926 38782 14978 38834
rect 15262 38782 15314 38834
rect 15598 38782 15650 38834
rect 16494 38782 16546 38834
rect 17726 38782 17778 38834
rect 17950 38782 18002 38834
rect 20302 38782 20354 38834
rect 20526 38782 20578 38834
rect 21758 38782 21810 38834
rect 25454 38782 25506 38834
rect 31278 38782 31330 38834
rect 33966 38782 34018 38834
rect 37326 38782 37378 38834
rect 37886 38782 37938 38834
rect 38222 38782 38274 38834
rect 38670 38782 38722 38834
rect 41582 38782 41634 38834
rect 42590 38782 42642 38834
rect 43374 38782 43426 38834
rect 43934 38782 43986 38834
rect 44606 38782 44658 38834
rect 45054 38782 45106 38834
rect 46622 38782 46674 38834
rect 49198 38782 49250 38834
rect 49646 38782 49698 38834
rect 50430 38782 50482 38834
rect 4622 38670 4674 38722
rect 6750 38670 6802 38722
rect 7534 38670 7586 38722
rect 12798 38670 12850 38722
rect 14254 38670 14306 38722
rect 18286 38670 18338 38722
rect 24670 38670 24722 38722
rect 26014 38670 26066 38722
rect 26462 38670 26514 38722
rect 27694 38670 27746 38722
rect 30830 38670 30882 38722
rect 34078 38670 34130 38722
rect 39230 38670 39282 38722
rect 42478 38670 42530 38722
rect 44158 38670 44210 38722
rect 46398 38670 46450 38722
rect 53342 38670 53394 38722
rect 17390 38558 17442 38610
rect 38558 38558 38610 38610
rect 47294 38558 47346 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 27022 38222 27074 38274
rect 45838 38222 45890 38274
rect 4622 38110 4674 38162
rect 8766 38110 8818 38162
rect 9662 38110 9714 38162
rect 17614 38110 17666 38162
rect 19966 38110 20018 38162
rect 21758 38110 21810 38162
rect 22990 38110 23042 38162
rect 27358 38110 27410 38162
rect 27918 38110 27970 38162
rect 32510 38110 32562 38162
rect 34638 38110 34690 38162
rect 55022 38110 55074 38162
rect 1822 37998 1874 38050
rect 5966 37998 6018 38050
rect 12574 37998 12626 38050
rect 14702 37998 14754 38050
rect 15038 37998 15090 38050
rect 15822 37998 15874 38050
rect 18174 37998 18226 38050
rect 24782 37998 24834 38050
rect 25230 37998 25282 38050
rect 28590 37998 28642 38050
rect 29486 37998 29538 38050
rect 30270 37998 30322 38050
rect 31726 37998 31778 38050
rect 37214 37998 37266 38050
rect 37998 37998 38050 38050
rect 38110 37998 38162 38050
rect 38222 37998 38274 38050
rect 38446 37998 38498 38050
rect 39678 37998 39730 38050
rect 43710 37998 43762 38050
rect 44718 37998 44770 38050
rect 45726 37998 45778 38050
rect 47070 37998 47122 38050
rect 48302 37998 48354 38050
rect 48974 37998 49026 38050
rect 49646 37998 49698 38050
rect 51326 37998 51378 38050
rect 51774 37998 51826 38050
rect 52894 37998 52946 38050
rect 54574 37998 54626 38050
rect 2494 37886 2546 37938
rect 6638 37886 6690 37938
rect 11790 37886 11842 37938
rect 14366 37886 14418 37938
rect 14814 37886 14866 37938
rect 18734 37886 18786 37938
rect 21422 37886 21474 37938
rect 23998 37886 24050 37938
rect 24334 37886 24386 37938
rect 26574 37886 26626 37938
rect 29822 37886 29874 37938
rect 30718 37886 30770 37938
rect 31054 37886 31106 37938
rect 37326 37886 37378 37938
rect 38782 37886 38834 37938
rect 39342 37886 39394 37938
rect 42478 37886 42530 37938
rect 42814 37886 42866 37938
rect 44942 37886 44994 37938
rect 45166 37886 45218 37938
rect 45390 37886 45442 37938
rect 45838 37886 45890 37938
rect 46398 37886 46450 37938
rect 48862 37886 48914 37938
rect 52782 37886 52834 37938
rect 53342 37886 53394 37938
rect 5070 37774 5122 37826
rect 9214 37774 9266 37826
rect 13694 37774 13746 37826
rect 14030 37774 14082 37826
rect 19630 37774 19682 37826
rect 21310 37774 21362 37826
rect 21870 37774 21922 37826
rect 22542 37774 22594 37826
rect 26014 37774 26066 37826
rect 26238 37774 26290 37826
rect 27246 37774 27298 37826
rect 28254 37774 28306 37826
rect 35086 37774 35138 37826
rect 36206 37774 36258 37826
rect 37102 37774 37154 37826
rect 37774 37774 37826 37826
rect 38670 37774 38722 37826
rect 39454 37774 39506 37826
rect 43486 37774 43538 37826
rect 43822 37774 43874 37826
rect 44382 37774 44434 37826
rect 51102 37774 51154 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 3502 37438 3554 37490
rect 4398 37438 4450 37490
rect 5182 37438 5234 37490
rect 6526 37438 6578 37490
rect 6638 37438 6690 37490
rect 14142 37438 14194 37490
rect 17502 37438 17554 37490
rect 18174 37438 18226 37490
rect 22990 37438 23042 37490
rect 31502 37438 31554 37490
rect 36430 37438 36482 37490
rect 40238 37438 40290 37490
rect 50206 37438 50258 37490
rect 50990 37438 51042 37490
rect 3726 37326 3778 37378
rect 3950 37326 4002 37378
rect 4622 37326 4674 37378
rect 4846 37326 4898 37378
rect 5518 37326 5570 37378
rect 6750 37326 6802 37378
rect 11790 37326 11842 37378
rect 15374 37326 15426 37378
rect 16382 37326 16434 37378
rect 17390 37326 17442 37378
rect 17838 37326 17890 37378
rect 20862 37326 20914 37378
rect 22094 37326 22146 37378
rect 24334 37326 24386 37378
rect 27918 37326 27970 37378
rect 36206 37326 36258 37378
rect 37102 37326 37154 37378
rect 37214 37326 37266 37378
rect 37662 37326 37714 37378
rect 37998 37326 38050 37378
rect 44158 37326 44210 37378
rect 45726 37326 45778 37378
rect 56142 37326 56194 37378
rect 3390 37214 3442 37266
rect 4286 37214 4338 37266
rect 11118 37214 11170 37266
rect 14366 37214 14418 37266
rect 15598 37214 15650 37266
rect 16046 37214 16098 37266
rect 18622 37214 18674 37266
rect 19070 37214 19122 37266
rect 19630 37214 19682 37266
rect 20078 37214 20130 37266
rect 20302 37214 20354 37266
rect 21198 37214 21250 37266
rect 21646 37214 21698 37266
rect 22430 37214 22482 37266
rect 23326 37214 23378 37266
rect 23886 37214 23938 37266
rect 24670 37214 24722 37266
rect 25230 37214 25282 37266
rect 25902 37214 25954 37266
rect 27246 37214 27298 37266
rect 30494 37214 30546 37266
rect 31166 37214 31218 37266
rect 32398 37214 32450 37266
rect 33070 37214 33122 37266
rect 36542 37214 36594 37266
rect 36990 37214 37042 37266
rect 38222 37214 38274 37266
rect 39790 37214 39842 37266
rect 43822 37214 43874 37266
rect 44830 37214 44882 37266
rect 45838 37214 45890 37266
rect 48750 37214 48802 37266
rect 48974 37214 49026 37266
rect 49422 37214 49474 37266
rect 54126 37214 54178 37266
rect 55022 37214 55074 37266
rect 13918 37102 13970 37154
rect 19854 37102 19906 37154
rect 24446 37102 24498 37154
rect 26126 37102 26178 37154
rect 26686 37102 26738 37154
rect 30046 37102 30098 37154
rect 30942 37102 30994 37154
rect 32062 37102 32114 37154
rect 33854 37102 33906 37154
rect 35982 37102 36034 37154
rect 40910 37102 40962 37154
rect 43038 37102 43090 37154
rect 45278 37102 45330 37154
rect 48190 37102 48242 37154
rect 49198 37102 49250 37154
rect 50430 37102 50482 37154
rect 51326 37102 51378 37154
rect 53454 37102 53506 37154
rect 54574 37102 54626 37154
rect 56702 37102 56754 37154
rect 57262 37102 57314 37154
rect 18622 36990 18674 37042
rect 22654 36990 22706 37042
rect 22990 36990 23042 37042
rect 54798 36990 54850 37042
rect 55470 36990 55522 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 14590 36654 14642 36706
rect 15598 36654 15650 36706
rect 33742 36654 33794 36706
rect 37214 36654 37266 36706
rect 37550 36654 37602 36706
rect 48862 36654 48914 36706
rect 16158 36542 16210 36594
rect 22094 36542 22146 36594
rect 22542 36542 22594 36594
rect 28142 36542 28194 36594
rect 28590 36542 28642 36594
rect 30046 36542 30098 36594
rect 33854 36542 33906 36594
rect 38558 36542 38610 36594
rect 39006 36542 39058 36594
rect 40350 36542 40402 36594
rect 42478 36542 42530 36594
rect 46846 36542 46898 36594
rect 47630 36542 47682 36594
rect 51662 36542 51714 36594
rect 54686 36542 54738 36594
rect 55582 36542 55634 36594
rect 13694 36430 13746 36482
rect 14030 36430 14082 36482
rect 14254 36430 14306 36482
rect 14478 36430 14530 36482
rect 15262 36430 15314 36482
rect 15934 36430 15986 36482
rect 17278 36430 17330 36482
rect 18958 36430 19010 36482
rect 19406 36430 19458 36482
rect 19742 36430 19794 36482
rect 20078 36430 20130 36482
rect 20526 36430 20578 36482
rect 21982 36430 22034 36482
rect 22430 36430 22482 36482
rect 23326 36430 23378 36482
rect 23998 36430 24050 36482
rect 27358 36430 27410 36482
rect 29486 36430 29538 36482
rect 31166 36430 31218 36482
rect 31502 36430 31554 36482
rect 36094 36430 36146 36482
rect 36990 36430 37042 36482
rect 38334 36430 38386 36482
rect 39566 36430 39618 36482
rect 43934 36430 43986 36482
rect 44830 36430 44882 36482
rect 45166 36430 45218 36482
rect 45278 36430 45330 36482
rect 45502 36430 45554 36482
rect 45726 36430 45778 36482
rect 46062 36430 46114 36482
rect 47742 36430 47794 36482
rect 48190 36430 48242 36482
rect 49870 36430 49922 36482
rect 50206 36430 50258 36482
rect 52670 36430 52722 36482
rect 54126 36430 54178 36482
rect 54798 36430 54850 36482
rect 55470 36430 55522 36482
rect 56030 36430 56082 36482
rect 56366 36430 56418 36482
rect 13806 36318 13858 36370
rect 18062 36318 18114 36370
rect 20750 36318 20802 36370
rect 25230 36318 25282 36370
rect 27694 36318 27746 36370
rect 32510 36318 32562 36370
rect 33966 36318 34018 36370
rect 35870 36318 35922 36370
rect 46398 36318 46450 36370
rect 47518 36318 47570 36370
rect 50878 36318 50930 36370
rect 52894 36318 52946 36370
rect 56702 36318 56754 36370
rect 57038 36318 57090 36370
rect 12910 36206 12962 36258
rect 14926 36206 14978 36258
rect 17166 36206 17218 36258
rect 19518 36206 19570 36258
rect 20302 36206 20354 36258
rect 23102 36206 23154 36258
rect 23774 36206 23826 36258
rect 23886 36206 23938 36258
rect 24558 36206 24610 36258
rect 24894 36206 24946 36258
rect 25566 36206 25618 36258
rect 30830 36206 30882 36258
rect 31838 36206 31890 36258
rect 32174 36206 32226 36258
rect 42926 36206 42978 36258
rect 43598 36206 43650 36258
rect 44270 36206 44322 36258
rect 45166 36206 45218 36258
rect 48638 36206 48690 36258
rect 48750 36206 48802 36258
rect 52110 36206 52162 36258
rect 53118 36206 53170 36258
rect 54014 36206 54066 36258
rect 56254 36206 56306 36258
rect 57150 36206 57202 36258
rect 57262 36206 57314 36258
rect 57822 36206 57874 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 14926 35870 14978 35922
rect 17390 35870 17442 35922
rect 18398 35870 18450 35922
rect 18622 35870 18674 35922
rect 18958 35870 19010 35922
rect 25230 35870 25282 35922
rect 25566 35870 25618 35922
rect 28030 35870 28082 35922
rect 29262 35870 29314 35922
rect 29374 35870 29426 35922
rect 29710 35870 29762 35922
rect 30270 35870 30322 35922
rect 30718 35870 30770 35922
rect 43486 35870 43538 35922
rect 43822 35870 43874 35922
rect 45502 35870 45554 35922
rect 45950 35870 46002 35922
rect 54574 35870 54626 35922
rect 57934 35870 57986 35922
rect 15822 35758 15874 35810
rect 16830 35758 16882 35810
rect 19070 35758 19122 35810
rect 21534 35758 21586 35810
rect 28590 35758 28642 35810
rect 30494 35758 30546 35810
rect 33742 35758 33794 35810
rect 36654 35758 36706 35810
rect 47070 35758 47122 35810
rect 54462 35758 54514 35810
rect 56030 35758 56082 35810
rect 12014 35646 12066 35698
rect 16046 35646 16098 35698
rect 17726 35646 17778 35698
rect 17950 35646 18002 35698
rect 22318 35646 22370 35698
rect 23214 35646 23266 35698
rect 23886 35646 23938 35698
rect 26126 35646 26178 35698
rect 28254 35646 28306 35698
rect 28814 35646 28866 35698
rect 29486 35646 29538 35698
rect 34078 35646 34130 35698
rect 37326 35646 37378 35698
rect 37550 35646 37602 35698
rect 38222 35646 38274 35698
rect 39118 35646 39170 35698
rect 39454 35646 39506 35698
rect 39790 35646 39842 35698
rect 40238 35646 40290 35698
rect 44718 35646 44770 35698
rect 44942 35646 44994 35698
rect 45166 35646 45218 35698
rect 45726 35646 45778 35698
rect 47630 35646 47682 35698
rect 47966 35646 48018 35698
rect 48750 35646 48802 35698
rect 49646 35646 49698 35698
rect 50766 35646 50818 35698
rect 51438 35646 51490 35698
rect 52558 35646 52610 35698
rect 54798 35646 54850 35698
rect 55358 35646 55410 35698
rect 56590 35646 56642 35698
rect 56926 35646 56978 35698
rect 57150 35646 57202 35698
rect 12686 35534 12738 35586
rect 15598 35534 15650 35586
rect 18510 35534 18562 35586
rect 19406 35534 19458 35586
rect 23438 35534 23490 35586
rect 27918 35534 27970 35586
rect 30382 35534 30434 35586
rect 38334 35534 38386 35586
rect 44382 35534 44434 35586
rect 45614 35534 45666 35586
rect 46622 35534 46674 35586
rect 50430 35534 50482 35586
rect 53342 35534 53394 35586
rect 55134 35534 55186 35586
rect 56702 35534 56754 35586
rect 57822 35534 57874 35586
rect 16382 35422 16434 35474
rect 16718 35422 16770 35474
rect 23326 35422 23378 35474
rect 39790 35422 39842 35474
rect 44606 35422 44658 35474
rect 48750 35422 48802 35474
rect 49086 35422 49138 35474
rect 57150 35422 57202 35474
rect 57710 35422 57762 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 13806 35086 13858 35138
rect 18958 35086 19010 35138
rect 29486 35086 29538 35138
rect 30606 35086 30658 35138
rect 34638 35086 34690 35138
rect 35086 35086 35138 35138
rect 43822 35086 43874 35138
rect 45278 35086 45330 35138
rect 51550 35086 51602 35138
rect 52894 35086 52946 35138
rect 57150 35086 57202 35138
rect 13582 34974 13634 35026
rect 15038 34974 15090 35026
rect 18174 34974 18226 35026
rect 18734 34974 18786 35026
rect 20526 34974 20578 35026
rect 22430 34974 22482 35026
rect 23886 34974 23938 35026
rect 26014 34974 26066 35026
rect 34414 34974 34466 35026
rect 34862 34974 34914 35026
rect 38110 34974 38162 35026
rect 40014 34974 40066 35026
rect 42142 34974 42194 35026
rect 47182 34974 47234 35026
rect 51102 34974 51154 35026
rect 53342 34974 53394 35026
rect 54126 34974 54178 35026
rect 15374 34862 15426 34914
rect 19294 34862 19346 34914
rect 19630 34862 19682 34914
rect 20638 34862 20690 34914
rect 21310 34862 21362 34914
rect 21422 34862 21474 34914
rect 23214 34862 23266 34914
rect 26462 34862 26514 34914
rect 27022 34862 27074 34914
rect 29150 34862 29202 34914
rect 30270 34862 30322 34914
rect 33406 34862 33458 34914
rect 39342 34862 39394 34914
rect 44158 34862 44210 34914
rect 44718 34862 44770 34914
rect 45166 34862 45218 34914
rect 45502 34862 45554 34914
rect 46286 34862 46338 34914
rect 47070 34862 47122 34914
rect 47294 34862 47346 34914
rect 48526 34862 48578 34914
rect 49310 34862 49362 34914
rect 49534 34862 49586 34914
rect 50990 34862 51042 34914
rect 52670 34862 52722 34914
rect 56814 34862 56866 34914
rect 57150 34862 57202 34914
rect 13582 34750 13634 34802
rect 16046 34750 16098 34802
rect 20750 34750 20802 34802
rect 21982 34750 22034 34802
rect 33182 34750 33234 34802
rect 37886 34750 37938 34802
rect 45726 34750 45778 34802
rect 46398 34750 46450 34802
rect 53230 34750 53282 34802
rect 53454 34750 53506 34802
rect 54350 34750 54402 34802
rect 56030 34750 56082 34802
rect 56590 34750 56642 34802
rect 57822 34750 57874 34802
rect 19070 34638 19122 34690
rect 29374 34638 29426 34690
rect 30494 34638 30546 34690
rect 33854 34638 33906 34690
rect 33966 34638 34018 34690
rect 34078 34638 34130 34690
rect 35534 34638 35586 34690
rect 36318 34638 36370 34690
rect 37102 34638 37154 34690
rect 42590 34638 42642 34690
rect 43486 34638 43538 34690
rect 43934 34638 43986 34690
rect 45166 34638 45218 34690
rect 46846 34638 46898 34690
rect 55918 34638 55970 34690
rect 57038 34638 57090 34690
rect 57710 34638 57762 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 15598 34302 15650 34354
rect 16382 34302 16434 34354
rect 21870 34302 21922 34354
rect 22766 34302 22818 34354
rect 25454 34302 25506 34354
rect 36430 34302 36482 34354
rect 46398 34302 46450 34354
rect 48974 34302 49026 34354
rect 49982 34302 50034 34354
rect 16606 34190 16658 34242
rect 16830 34190 16882 34242
rect 25902 34190 25954 34242
rect 27134 34190 27186 34242
rect 30382 34190 30434 34242
rect 36542 34190 36594 34242
rect 41022 34190 41074 34242
rect 42590 34190 42642 34242
rect 43822 34190 43874 34242
rect 48190 34190 48242 34242
rect 50206 34190 50258 34242
rect 50654 34190 50706 34242
rect 56030 34190 56082 34242
rect 14478 34078 14530 34130
rect 16270 34078 16322 34130
rect 17950 34078 18002 34130
rect 20862 34078 20914 34130
rect 24670 34078 24722 34130
rect 26462 34078 26514 34130
rect 29598 34078 29650 34130
rect 33182 34078 33234 34130
rect 37102 34078 37154 34130
rect 38782 34078 38834 34130
rect 40910 34078 40962 34130
rect 42030 34078 42082 34130
rect 43150 34078 43202 34130
rect 47630 34078 47682 34130
rect 48078 34078 48130 34130
rect 48750 34078 48802 34130
rect 49198 34078 49250 34130
rect 49422 34078 49474 34130
rect 51774 34078 51826 34130
rect 53118 34078 53170 34130
rect 53566 34078 53618 34130
rect 53902 34078 53954 34130
rect 56478 34078 56530 34130
rect 56814 34078 56866 34130
rect 57262 34078 57314 34130
rect 19742 33966 19794 34018
rect 20302 33966 20354 34018
rect 21310 33966 21362 34018
rect 23214 33966 23266 34018
rect 24446 33966 24498 34018
rect 29262 33966 29314 34018
rect 32510 33966 32562 34018
rect 33854 33966 33906 34018
rect 35982 33966 36034 34018
rect 37214 33966 37266 34018
rect 41694 33966 41746 34018
rect 45950 33966 46002 34018
rect 49086 33966 49138 34018
rect 49870 33966 49922 34018
rect 55582 33966 55634 34018
rect 57374 33966 57426 34018
rect 14478 33854 14530 33906
rect 14814 33854 14866 33906
rect 24334 33854 24386 33906
rect 26014 33854 26066 33906
rect 36430 33854 36482 33906
rect 38222 33854 38274 33906
rect 51214 33854 51266 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 44046 33518 44098 33570
rect 47182 33518 47234 33570
rect 50094 33518 50146 33570
rect 14254 33406 14306 33458
rect 16382 33406 16434 33458
rect 17278 33406 17330 33458
rect 19406 33406 19458 33458
rect 20078 33406 20130 33458
rect 24446 33406 24498 33458
rect 29934 33406 29986 33458
rect 30382 33406 30434 33458
rect 32734 33406 32786 33458
rect 33518 33406 33570 33458
rect 39902 33406 39954 33458
rect 42254 33406 42306 33458
rect 51214 33406 51266 33458
rect 51662 33406 51714 33458
rect 55806 33406 55858 33458
rect 57934 33406 57986 33458
rect 13582 33294 13634 33346
rect 18062 33294 18114 33346
rect 18846 33294 18898 33346
rect 22542 33294 22594 33346
rect 23662 33294 23714 33346
rect 29486 33294 29538 33346
rect 35086 33294 35138 33346
rect 35758 33294 35810 33346
rect 36318 33294 36370 33346
rect 37102 33294 37154 33346
rect 43934 33294 43986 33346
rect 47070 33294 47122 33346
rect 49982 33294 50034 33346
rect 50878 33294 50930 33346
rect 51102 33294 51154 33346
rect 53566 33294 53618 33346
rect 54014 33294 54066 33346
rect 55022 33294 55074 33346
rect 16830 33182 16882 33234
rect 18734 33182 18786 33234
rect 22206 33182 22258 33234
rect 29150 33182 29202 33234
rect 33070 33182 33122 33234
rect 34750 33182 34802 33234
rect 35422 33182 35474 33234
rect 36206 33182 36258 33234
rect 37774 33182 37826 33234
rect 46510 33182 46562 33234
rect 46734 33182 46786 33234
rect 52110 33182 52162 33234
rect 53006 33182 53058 33234
rect 54686 33182 54738 33234
rect 17950 33070 18002 33122
rect 20526 33070 20578 33122
rect 21422 33070 21474 33122
rect 21870 33070 21922 33122
rect 22318 33070 22370 33122
rect 23326 33070 23378 33122
rect 26686 33070 26738 33122
rect 29262 33070 29314 33122
rect 36430 33070 36482 33122
rect 40350 33070 40402 33122
rect 42814 33070 42866 33122
rect 43262 33070 43314 33122
rect 43822 33070 43874 33122
rect 46622 33070 46674 33122
rect 47182 33070 47234 33122
rect 54126 33070 54178 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 16382 32734 16434 32786
rect 31950 32734 32002 32786
rect 34078 32734 34130 32786
rect 35646 32734 35698 32786
rect 37326 32734 37378 32786
rect 42142 32734 42194 32786
rect 43374 32734 43426 32786
rect 46398 32734 46450 32786
rect 46846 32734 46898 32786
rect 47182 32734 47234 32786
rect 52222 32734 52274 32786
rect 56702 32734 56754 32786
rect 29374 32622 29426 32674
rect 33742 32622 33794 32674
rect 34302 32622 34354 32674
rect 36878 32622 36930 32674
rect 46958 32622 47010 32674
rect 50094 32622 50146 32674
rect 50206 32622 50258 32674
rect 51662 32622 51714 32674
rect 52782 32622 52834 32674
rect 54798 32622 54850 32674
rect 12462 32510 12514 32562
rect 18286 32510 18338 32562
rect 23662 32510 23714 32562
rect 24446 32510 24498 32562
rect 30158 32510 30210 32562
rect 30830 32510 30882 32562
rect 31278 32510 31330 32562
rect 33966 32510 34018 32562
rect 37102 32510 37154 32562
rect 37438 32510 37490 32562
rect 41806 32510 41858 32562
rect 43710 32510 43762 32562
rect 43934 32510 43986 32562
rect 44382 32510 44434 32562
rect 45838 32510 45890 32562
rect 46062 32510 46114 32562
rect 47518 32510 47570 32562
rect 49310 32510 49362 32562
rect 49758 32510 49810 32562
rect 50766 32510 50818 32562
rect 51774 32510 51826 32562
rect 52110 32510 52162 32562
rect 54238 32510 54290 32562
rect 13134 32398 13186 32450
rect 15262 32398 15314 32450
rect 15822 32398 15874 32450
rect 18958 32398 19010 32450
rect 21086 32398 21138 32450
rect 21534 32398 21586 32450
rect 27246 32398 27298 32450
rect 32398 32398 32450 32450
rect 33182 32398 33234 32450
rect 41582 32398 41634 32450
rect 42926 32398 42978 32450
rect 43822 32398 43874 32450
rect 48862 32398 48914 32450
rect 51326 32398 51378 32450
rect 15934 32286 15986 32338
rect 46286 32286 46338 32338
rect 46510 32286 46562 32338
rect 50206 32286 50258 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 25342 31950 25394 32002
rect 37550 31950 37602 32002
rect 38110 31950 38162 32002
rect 46958 31950 47010 32002
rect 50990 31950 51042 32002
rect 13918 31838 13970 31890
rect 14478 31838 14530 31890
rect 14814 31838 14866 31890
rect 15598 31838 15650 31890
rect 18958 31838 19010 31890
rect 21870 31838 21922 31890
rect 24894 31838 24946 31890
rect 25678 31838 25730 31890
rect 26462 31838 26514 31890
rect 27358 31838 27410 31890
rect 33630 31838 33682 31890
rect 36206 31838 36258 31890
rect 44270 31838 44322 31890
rect 44942 31838 44994 31890
rect 51998 31838 52050 31890
rect 53118 31838 53170 31890
rect 55246 31838 55298 31890
rect 57374 31838 57426 31890
rect 13806 31726 13858 31778
rect 14142 31726 14194 31778
rect 15710 31726 15762 31778
rect 16494 31726 16546 31778
rect 17502 31726 17554 31778
rect 19070 31726 19122 31778
rect 20078 31726 20130 31778
rect 20526 31726 20578 31778
rect 21310 31726 21362 31778
rect 22654 31726 22706 31778
rect 26686 31726 26738 31778
rect 30382 31726 30434 31778
rect 32174 31726 32226 31778
rect 32734 31726 32786 31778
rect 33854 31726 33906 31778
rect 37326 31726 37378 31778
rect 37550 31726 37602 31778
rect 41470 31726 41522 31778
rect 46734 31726 46786 31778
rect 47182 31726 47234 31778
rect 49086 31726 49138 31778
rect 50990 31726 51042 31778
rect 51326 31726 51378 31778
rect 52670 31726 52722 31778
rect 54014 31726 54066 31778
rect 54798 31726 54850 31778
rect 58046 31726 58098 31778
rect 14590 31614 14642 31666
rect 16158 31614 16210 31666
rect 16606 31614 16658 31666
rect 18734 31614 18786 31666
rect 20414 31614 20466 31666
rect 20750 31614 20802 31666
rect 21534 31614 21586 31666
rect 22542 31614 22594 31666
rect 25006 31614 25058 31666
rect 25566 31614 25618 31666
rect 26014 31614 26066 31666
rect 26238 31614 26290 31666
rect 30046 31614 30098 31666
rect 31614 31614 31666 31666
rect 32510 31614 32562 31666
rect 33182 31614 33234 31666
rect 33406 31614 33458 31666
rect 34078 31614 34130 31666
rect 36990 31614 37042 31666
rect 38222 31614 38274 31666
rect 39678 31614 39730 31666
rect 40014 31614 40066 31666
rect 42142 31614 42194 31666
rect 47966 31614 48018 31666
rect 48190 31614 48242 31666
rect 48414 31614 48466 31666
rect 51550 31614 51602 31666
rect 51886 31614 51938 31666
rect 54238 31614 54290 31666
rect 15598 31502 15650 31554
rect 15934 31502 15986 31554
rect 17614 31502 17666 31554
rect 17726 31502 17778 31554
rect 20302 31502 20354 31554
rect 26462 31502 26514 31554
rect 33966 31502 34018 31554
rect 34526 31502 34578 31554
rect 37102 31502 37154 31554
rect 38670 31502 38722 31554
rect 39342 31502 39394 31554
rect 40350 31502 40402 31554
rect 47630 31502 47682 31554
rect 48302 31502 48354 31554
rect 48750 31502 48802 31554
rect 49758 31502 49810 31554
rect 49982 31502 50034 31554
rect 50094 31502 50146 31554
rect 50206 31502 50258 31554
rect 51438 31502 51490 31554
rect 54574 31502 54626 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 13246 31166 13298 31218
rect 24670 31166 24722 31218
rect 29710 31166 29762 31218
rect 40014 31166 40066 31218
rect 40910 31166 40962 31218
rect 41806 31166 41858 31218
rect 43150 31166 43202 31218
rect 43486 31166 43538 31218
rect 44270 31166 44322 31218
rect 45502 31166 45554 31218
rect 49422 31166 49474 31218
rect 13470 31054 13522 31106
rect 13806 31054 13858 31106
rect 29150 31054 29202 31106
rect 30158 31054 30210 31106
rect 33854 31054 33906 31106
rect 37102 31054 37154 31106
rect 39902 31054 39954 31106
rect 40126 31054 40178 31106
rect 42142 31054 42194 31106
rect 42590 31054 42642 31106
rect 42814 31054 42866 31106
rect 44158 31054 44210 31106
rect 44718 31054 44770 31106
rect 50542 31054 50594 31106
rect 51886 31054 51938 31106
rect 52110 31054 52162 31106
rect 14142 30942 14194 30994
rect 15822 30942 15874 30994
rect 16158 30942 16210 30994
rect 17838 30942 17890 30994
rect 18734 30942 18786 30994
rect 21422 30942 21474 30994
rect 22990 30942 23042 30994
rect 28030 30942 28082 30994
rect 30046 30942 30098 30994
rect 33070 30942 33122 30994
rect 36430 30942 36482 30994
rect 44382 30942 44434 30994
rect 44942 30942 44994 30994
rect 45278 30942 45330 30994
rect 45614 30942 45666 30994
rect 46510 30942 46562 30994
rect 47406 30942 47458 30994
rect 49198 30942 49250 30994
rect 49422 30942 49474 30994
rect 49758 30942 49810 30994
rect 50094 30942 50146 30994
rect 50206 30942 50258 30994
rect 52558 30942 52610 30994
rect 53790 30942 53842 30994
rect 54910 30942 54962 30994
rect 55358 30942 55410 30994
rect 16830 30830 16882 30882
rect 17390 30830 17442 30882
rect 18286 30830 18338 30882
rect 19070 30830 19122 30882
rect 22094 30830 22146 30882
rect 23326 30830 23378 30882
rect 25230 30830 25282 30882
rect 27358 30830 27410 30882
rect 30718 30830 30770 30882
rect 35982 30830 36034 30882
rect 39230 30830 39282 30882
rect 41358 30830 41410 30882
rect 42478 30830 42530 30882
rect 46734 30830 46786 30882
rect 47966 30830 48018 30882
rect 50430 30830 50482 30882
rect 50990 30830 51042 30882
rect 52334 30830 52386 30882
rect 52782 30830 52834 30882
rect 53902 30830 53954 30882
rect 13134 30718 13186 30770
rect 14142 30718 14194 30770
rect 18734 30718 18786 30770
rect 21982 30718 22034 30770
rect 24110 30718 24162 30770
rect 29262 30718 29314 30770
rect 30158 30718 30210 30770
rect 30606 30718 30658 30770
rect 45054 30718 45106 30770
rect 46958 30718 47010 30770
rect 47070 30718 47122 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 18622 30382 18674 30434
rect 21310 30382 21362 30434
rect 22766 30382 22818 30434
rect 26350 30382 26402 30434
rect 39006 30382 39058 30434
rect 11790 30270 11842 30322
rect 47742 30270 47794 30322
rect 53454 30270 53506 30322
rect 53678 30270 53730 30322
rect 54574 30270 54626 30322
rect 8990 30158 9042 30210
rect 12238 30158 12290 30210
rect 16718 30158 16770 30210
rect 17166 30158 17218 30210
rect 17390 30158 17442 30210
rect 18622 30158 18674 30210
rect 19518 30158 19570 30210
rect 21646 30158 21698 30210
rect 21870 30158 21922 30210
rect 22094 30158 22146 30210
rect 22430 30158 22482 30210
rect 25790 30158 25842 30210
rect 26126 30158 26178 30210
rect 26574 30158 26626 30210
rect 27134 30158 27186 30210
rect 28366 30158 28418 30210
rect 28702 30158 28754 30210
rect 29038 30158 29090 30210
rect 29486 30158 29538 30210
rect 29598 30158 29650 30210
rect 31054 30158 31106 30210
rect 35758 30158 35810 30210
rect 35870 30158 35922 30210
rect 37438 30158 37490 30210
rect 38222 30158 38274 30210
rect 38670 30158 38722 30210
rect 39230 30158 39282 30210
rect 39790 30158 39842 30210
rect 40238 30158 40290 30210
rect 41134 30158 41186 30210
rect 41694 30158 41746 30210
rect 42030 30158 42082 30210
rect 42590 30158 42642 30210
rect 43038 30158 43090 30210
rect 46398 30158 46450 30210
rect 47070 30158 47122 30210
rect 47854 30158 47906 30210
rect 49534 30158 49586 30210
rect 51886 30158 51938 30210
rect 56702 30158 56754 30210
rect 57374 30158 57426 30210
rect 9662 30046 9714 30098
rect 15710 30046 15762 30098
rect 16606 30046 16658 30098
rect 20078 30046 20130 30098
rect 21422 30046 21474 30098
rect 22318 30046 22370 30098
rect 22878 30046 22930 30098
rect 26910 30046 26962 30098
rect 28478 30046 28530 30098
rect 34414 30046 34466 30098
rect 37662 30046 37714 30098
rect 46062 30046 46114 30098
rect 47294 30046 47346 30098
rect 48862 30046 48914 30098
rect 49870 30046 49922 30098
rect 52110 30046 52162 30098
rect 53006 30046 53058 30098
rect 15934 29934 15986 29986
rect 16046 29934 16098 29986
rect 16158 29934 16210 29986
rect 16494 29934 16546 29986
rect 26574 29934 26626 29986
rect 29262 29934 29314 29986
rect 40574 29934 40626 29986
rect 43262 29934 43314 29986
rect 45726 29934 45778 29986
rect 46734 29934 46786 29986
rect 47630 29934 47682 29986
rect 48078 29934 48130 29986
rect 48526 29934 48578 29986
rect 49422 29934 49474 29986
rect 49646 29934 49698 29986
rect 51550 29934 51602 29986
rect 52782 29934 52834 29986
rect 52894 29934 52946 29986
rect 54014 29934 54066 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 9774 29598 9826 29650
rect 19406 29598 19458 29650
rect 27694 29598 27746 29650
rect 31950 29598 32002 29650
rect 35198 29598 35250 29650
rect 41022 29598 41074 29650
rect 46958 29598 47010 29650
rect 47406 29598 47458 29650
rect 49310 29598 49362 29650
rect 12910 29486 12962 29538
rect 18062 29486 18114 29538
rect 18846 29486 18898 29538
rect 23662 29486 23714 29538
rect 28814 29486 28866 29538
rect 34526 29486 34578 29538
rect 39902 29486 39954 29538
rect 46062 29486 46114 29538
rect 50430 29486 50482 29538
rect 5742 29374 5794 29426
rect 10110 29374 10162 29426
rect 12238 29374 12290 29426
rect 17390 29374 17442 29426
rect 17950 29374 18002 29426
rect 22094 29374 22146 29426
rect 23998 29374 24050 29426
rect 24670 29374 24722 29426
rect 25902 29374 25954 29426
rect 28030 29374 28082 29426
rect 32286 29374 32338 29426
rect 33070 29374 33122 29426
rect 33742 29374 33794 29426
rect 33966 29374 34018 29426
rect 34750 29374 34802 29426
rect 34974 29374 35026 29426
rect 35310 29374 35362 29426
rect 40126 29374 40178 29426
rect 45166 29374 45218 29426
rect 45390 29374 45442 29426
rect 45838 29374 45890 29426
rect 46398 29374 46450 29426
rect 46622 29374 46674 29426
rect 47070 29374 47122 29426
rect 47182 29374 47234 29426
rect 49086 29374 49138 29426
rect 49198 29374 49250 29426
rect 49534 29374 49586 29426
rect 50094 29374 50146 29426
rect 51662 29374 51714 29426
rect 53230 29374 53282 29426
rect 53902 29374 53954 29426
rect 54798 29374 54850 29426
rect 55358 29374 55410 29426
rect 6414 29262 6466 29314
rect 8542 29262 8594 29314
rect 8990 29262 9042 29314
rect 15038 29262 15090 29314
rect 15486 29262 15538 29314
rect 18398 29262 18450 29314
rect 21982 29262 22034 29314
rect 22766 29262 22818 29314
rect 25230 29262 25282 29314
rect 25566 29262 25618 29314
rect 30942 29262 30994 29314
rect 32510 29262 32562 29314
rect 34414 29262 34466 29314
rect 44494 29262 44546 29314
rect 44830 29262 44882 29314
rect 45614 29262 45666 29314
rect 46174 29262 46226 29314
rect 50878 29262 50930 29314
rect 54350 29262 54402 29314
rect 24334 29150 24386 29202
rect 24670 29150 24722 29202
rect 55134 29150 55186 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 10558 28814 10610 28866
rect 18286 28814 18338 28866
rect 21310 28814 21362 28866
rect 27582 28814 27634 28866
rect 28254 28814 28306 28866
rect 29150 28814 29202 28866
rect 45166 28814 45218 28866
rect 53230 28814 53282 28866
rect 14254 28702 14306 28754
rect 16382 28702 16434 28754
rect 16830 28702 16882 28754
rect 25342 28702 25394 28754
rect 28590 28702 28642 28754
rect 30046 28702 30098 28754
rect 32174 28702 32226 28754
rect 33406 28702 33458 28754
rect 35086 28702 35138 28754
rect 36318 28702 36370 28754
rect 37662 28702 37714 28754
rect 38110 28702 38162 28754
rect 38558 28702 38610 28754
rect 41918 28702 41970 28754
rect 42366 28702 42418 28754
rect 43374 28702 43426 28754
rect 43822 28702 43874 28754
rect 44270 28702 44322 28754
rect 49310 28702 49362 28754
rect 51438 28702 51490 28754
rect 52110 28702 52162 28754
rect 53118 28702 53170 28754
rect 54910 28702 54962 28754
rect 7086 28590 7138 28642
rect 7534 28590 7586 28642
rect 7870 28590 7922 28642
rect 10894 28590 10946 28642
rect 11566 28590 11618 28642
rect 13470 28590 13522 28642
rect 21646 28590 21698 28642
rect 23438 28590 23490 28642
rect 24894 28590 24946 28642
rect 25230 28590 25282 28642
rect 27358 28590 27410 28642
rect 27918 28590 27970 28642
rect 29486 28590 29538 28642
rect 32286 28590 32338 28642
rect 33294 28590 33346 28642
rect 33630 28590 33682 28642
rect 33854 28590 33906 28642
rect 34078 28590 34130 28642
rect 34414 28590 34466 28642
rect 34750 28590 34802 28642
rect 37214 28590 37266 28642
rect 41470 28590 41522 28642
rect 42926 28590 42978 28642
rect 45614 28590 45666 28642
rect 46846 28590 46898 28642
rect 47630 28590 47682 28642
rect 48526 28590 48578 28642
rect 53006 28590 53058 28642
rect 53790 28590 53842 28642
rect 54238 28590 54290 28642
rect 55358 28590 55410 28642
rect 55694 28590 55746 28642
rect 56478 28590 56530 28642
rect 6750 28478 6802 28530
rect 8094 28478 8146 28530
rect 8654 28478 8706 28530
rect 11678 28478 11730 28530
rect 18398 28478 18450 28530
rect 26238 28478 26290 28530
rect 27134 28478 27186 28530
rect 28478 28478 28530 28530
rect 32958 28478 33010 28530
rect 35534 28478 35586 28530
rect 40686 28478 40738 28530
rect 45054 28478 45106 28530
rect 46622 28478 46674 28530
rect 47294 28478 47346 28530
rect 51774 28478 51826 28530
rect 55022 28478 55074 28530
rect 56254 28478 56306 28530
rect 19630 28366 19682 28418
rect 21422 28366 21474 28418
rect 22878 28366 22930 28418
rect 27582 28366 27634 28418
rect 29262 28366 29314 28418
rect 34302 28366 34354 28418
rect 35086 28366 35138 28418
rect 35310 28366 35362 28418
rect 42254 28366 42306 28418
rect 42478 28366 42530 28418
rect 46958 28366 47010 28418
rect 48190 28366 48242 28418
rect 51998 28366 52050 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 12910 28030 12962 28082
rect 17502 28030 17554 28082
rect 19070 28030 19122 28082
rect 31838 28030 31890 28082
rect 32174 28030 32226 28082
rect 32398 28030 32450 28082
rect 41022 28030 41074 28082
rect 47742 28030 47794 28082
rect 48862 28030 48914 28082
rect 49534 28030 49586 28082
rect 8206 27918 8258 27970
rect 8878 27918 8930 27970
rect 14478 27918 14530 27970
rect 20414 27918 20466 27970
rect 27694 27918 27746 27970
rect 36542 27918 36594 27970
rect 38446 27918 38498 27970
rect 39678 27918 39730 27970
rect 42366 27918 42418 27970
rect 49982 27918 50034 27970
rect 51774 27918 51826 27970
rect 53902 27918 53954 27970
rect 54126 27918 54178 27970
rect 56590 27918 56642 27970
rect 4062 27806 4114 27858
rect 7646 27806 7698 27858
rect 8094 27806 8146 27858
rect 9550 27806 9602 27858
rect 13806 27806 13858 27858
rect 19742 27806 19794 27858
rect 23998 27806 24050 27858
rect 24334 27806 24386 27858
rect 28366 27806 28418 27858
rect 28814 27806 28866 27858
rect 32510 27806 32562 27858
rect 33182 27806 33234 27858
rect 36430 27806 36482 27858
rect 38558 27806 38610 27858
rect 41694 27806 41746 27858
rect 44830 27806 44882 27858
rect 47854 27806 47906 27858
rect 48974 27806 49026 27858
rect 50430 27806 50482 27858
rect 51662 27806 51714 27858
rect 52334 27806 52386 27858
rect 52782 27806 52834 27858
rect 53454 27806 53506 27858
rect 55022 27806 55074 27858
rect 55582 27806 55634 27858
rect 56814 27806 56866 27858
rect 4734 27694 4786 27746
rect 6862 27694 6914 27746
rect 10334 27694 10386 27746
rect 12462 27694 12514 27746
rect 16606 27694 16658 27746
rect 22542 27694 22594 27746
rect 22990 27694 23042 27746
rect 24110 27694 24162 27746
rect 24558 27694 24610 27746
rect 25566 27694 25618 27746
rect 29598 27694 29650 27746
rect 33966 27694 34018 27746
rect 36094 27694 36146 27746
rect 40910 27694 40962 27746
rect 44494 27694 44546 27746
rect 46286 27694 46338 27746
rect 50766 27694 50818 27746
rect 54238 27694 54290 27746
rect 7310 27582 7362 27634
rect 8990 27582 9042 27634
rect 18958 27582 19010 27634
rect 19294 27582 19346 27634
rect 41246 27582 41298 27634
rect 49086 27582 49138 27634
rect 52222 27582 52274 27634
rect 53230 27582 53282 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 33742 27246 33794 27298
rect 42366 27246 42418 27298
rect 45054 27246 45106 27298
rect 53230 27246 53282 27298
rect 7534 27134 7586 27186
rect 11118 27134 11170 27186
rect 17166 27134 17218 27186
rect 19294 27134 19346 27186
rect 19630 27134 19682 27186
rect 21310 27134 21362 27186
rect 26350 27134 26402 27186
rect 28478 27134 28530 27186
rect 31502 27134 31554 27186
rect 32174 27134 32226 27186
rect 32958 27134 33010 27186
rect 37326 27134 37378 27186
rect 40014 27134 40066 27186
rect 40462 27134 40514 27186
rect 41806 27134 41858 27186
rect 43598 27134 43650 27186
rect 44830 27134 44882 27186
rect 45390 27134 45442 27186
rect 47406 27134 47458 27186
rect 52782 27134 52834 27186
rect 55582 27134 55634 27186
rect 57710 27134 57762 27186
rect 5966 27022 6018 27074
rect 9998 27022 10050 27074
rect 10782 27022 10834 27074
rect 11566 27022 11618 27074
rect 16382 27022 16434 27074
rect 20078 27022 20130 27074
rect 20526 27022 20578 27074
rect 21758 27022 21810 27074
rect 22206 27022 22258 27074
rect 22542 27022 22594 27074
rect 23102 27022 23154 27074
rect 23438 27022 23490 27074
rect 31614 27022 31666 27074
rect 32286 27022 32338 27074
rect 33294 27022 33346 27074
rect 33518 27022 33570 27074
rect 33966 27022 34018 27074
rect 34302 27022 34354 27074
rect 34750 27022 34802 27074
rect 35646 27022 35698 27074
rect 35982 27022 36034 27074
rect 36430 27022 36482 27074
rect 38334 27022 38386 27074
rect 38782 27022 38834 27074
rect 39230 27022 39282 27074
rect 41918 27022 41970 27074
rect 42142 27022 42194 27074
rect 42814 27022 42866 27074
rect 43262 27022 43314 27074
rect 44158 27022 44210 27074
rect 45726 27022 45778 27074
rect 48750 27022 48802 27074
rect 49646 27022 49698 27074
rect 50542 27022 50594 27074
rect 51438 27022 51490 27074
rect 51774 27022 51826 27074
rect 53678 27022 53730 27074
rect 53790 27022 53842 27074
rect 54014 27022 54066 27074
rect 54910 27022 54962 27074
rect 5630 26910 5682 26962
rect 10334 26910 10386 26962
rect 11902 26910 11954 26962
rect 13470 26910 13522 26962
rect 13806 26910 13858 26962
rect 24222 26910 24274 26962
rect 34526 26910 34578 26962
rect 36206 26910 36258 26962
rect 41134 26910 41186 26962
rect 41694 26910 41746 26962
rect 42702 26910 42754 26962
rect 43038 26910 43090 26962
rect 49758 26910 49810 26962
rect 50430 26910 50482 26962
rect 51214 26910 51266 26962
rect 52110 26910 52162 26962
rect 54462 26910 54514 26962
rect 7086 26798 7138 26850
rect 7646 26798 7698 26850
rect 22654 26798 22706 26850
rect 22878 26798 22930 26850
rect 33182 26798 33234 26850
rect 35646 26798 35698 26850
rect 37214 26798 37266 26850
rect 38670 26798 38722 26850
rect 38894 26798 38946 26850
rect 39342 26798 39394 26850
rect 39454 26798 39506 26850
rect 41246 26798 41298 26850
rect 48526 26798 48578 26850
rect 51102 26798 51154 26850
rect 51998 26798 52050 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 10110 26462 10162 26514
rect 15710 26462 15762 26514
rect 22766 26462 22818 26514
rect 24222 26462 24274 26514
rect 36094 26462 36146 26514
rect 36990 26462 37042 26514
rect 42702 26462 42754 26514
rect 43598 26462 43650 26514
rect 44046 26462 44098 26514
rect 46734 26462 46786 26514
rect 48862 26462 48914 26514
rect 7534 26350 7586 26402
rect 10558 26350 10610 26402
rect 13134 26350 13186 26402
rect 21086 26350 21138 26402
rect 21870 26350 21922 26402
rect 22542 26350 22594 26402
rect 22990 26350 23042 26402
rect 29038 26350 29090 26402
rect 29710 26350 29762 26402
rect 32398 26350 32450 26402
rect 34526 26350 34578 26402
rect 39342 26350 39394 26402
rect 44494 26350 44546 26402
rect 47630 26350 47682 26402
rect 49422 26350 49474 26402
rect 53454 26350 53506 26402
rect 53902 26350 53954 26402
rect 6974 26238 7026 26290
rect 7422 26238 7474 26290
rect 10894 26238 10946 26290
rect 12350 26238 12402 26290
rect 18958 26238 19010 26290
rect 19518 26238 19570 26290
rect 20414 26238 20466 26290
rect 20750 26238 20802 26290
rect 21198 26238 21250 26290
rect 21422 26238 21474 26290
rect 21646 26238 21698 26290
rect 22318 26238 22370 26290
rect 23102 26238 23154 26290
rect 23550 26238 23602 26290
rect 24110 26238 24162 26290
rect 24334 26238 24386 26290
rect 25118 26238 25170 26290
rect 25454 26238 25506 26290
rect 25678 26238 25730 26290
rect 28702 26238 28754 26290
rect 29486 26238 29538 26290
rect 31614 26238 31666 26290
rect 32062 26238 32114 26290
rect 33070 26238 33122 26290
rect 33294 26238 33346 26290
rect 33518 26238 33570 26290
rect 33630 26238 33682 26290
rect 34078 26238 34130 26290
rect 34414 26238 34466 26290
rect 35310 26238 35362 26290
rect 35534 26238 35586 26290
rect 35982 26238 36034 26290
rect 36206 26238 36258 26290
rect 36542 26238 36594 26290
rect 40126 26238 40178 26290
rect 40910 26238 40962 26290
rect 41246 26238 41298 26290
rect 41470 26238 41522 26290
rect 41918 26238 41970 26290
rect 44382 26238 44434 26290
rect 48190 26238 48242 26290
rect 49534 26238 49586 26290
rect 49870 26238 49922 26290
rect 50990 26238 51042 26290
rect 51326 26238 51378 26290
rect 51550 26238 51602 26290
rect 52334 26238 52386 26290
rect 53342 26238 53394 26290
rect 54350 26238 54402 26290
rect 54798 26238 54850 26290
rect 15262 26126 15314 26178
rect 18622 26126 18674 26178
rect 20862 26126 20914 26178
rect 23886 26126 23938 26178
rect 25342 26126 25394 26178
rect 26686 26126 26738 26178
rect 33182 26126 33234 26178
rect 35758 26126 35810 26178
rect 37214 26126 37266 26178
rect 41022 26126 41074 26178
rect 51438 26126 51490 26178
rect 52222 26126 52274 26178
rect 6638 26014 6690 26066
rect 26126 26014 26178 26066
rect 26462 26014 26514 26066
rect 32510 26014 32562 26066
rect 34526 26014 34578 26066
rect 50990 26014 51042 26066
rect 52446 26014 52498 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 10670 25678 10722 25730
rect 13582 25678 13634 25730
rect 13918 25678 13970 25730
rect 39566 25678 39618 25730
rect 46510 25678 46562 25730
rect 53902 25678 53954 25730
rect 9886 25566 9938 25618
rect 12798 25566 12850 25618
rect 18398 25566 18450 25618
rect 25678 25566 25730 25618
rect 27806 25566 27858 25618
rect 30494 25566 30546 25618
rect 32622 25566 32674 25618
rect 33966 25566 34018 25618
rect 40126 25566 40178 25618
rect 41246 25566 41298 25618
rect 45278 25566 45330 25618
rect 46958 25566 47010 25618
rect 47294 25566 47346 25618
rect 50878 25566 50930 25618
rect 52894 25566 52946 25618
rect 54014 25566 54066 25618
rect 5966 25454 6018 25506
rect 7086 25454 7138 25506
rect 11454 25454 11506 25506
rect 12238 25454 12290 25506
rect 15598 25454 15650 25506
rect 20302 25454 20354 25506
rect 21646 25454 21698 25506
rect 23550 25454 23602 25506
rect 23998 25454 24050 25506
rect 24334 25454 24386 25506
rect 24894 25454 24946 25506
rect 28590 25454 28642 25506
rect 29710 25454 29762 25506
rect 33070 25454 33122 25506
rect 36206 25454 36258 25506
rect 37102 25454 37154 25506
rect 37998 25454 38050 25506
rect 38222 25454 38274 25506
rect 39902 25454 39954 25506
rect 40014 25454 40066 25506
rect 40798 25454 40850 25506
rect 42254 25454 42306 25506
rect 42814 25454 42866 25506
rect 43150 25454 43202 25506
rect 44942 25454 44994 25506
rect 45726 25454 45778 25506
rect 45950 25454 46002 25506
rect 46062 25454 46114 25506
rect 47406 25454 47458 25506
rect 47630 25454 47682 25506
rect 49198 25454 49250 25506
rect 50654 25454 50706 25506
rect 52782 25454 52834 25506
rect 7758 25342 7810 25394
rect 11230 25342 11282 25394
rect 11902 25342 11954 25394
rect 14142 25342 14194 25394
rect 14702 25342 14754 25394
rect 16270 25342 16322 25394
rect 19294 25342 19346 25394
rect 19854 25342 19906 25394
rect 20750 25342 20802 25394
rect 29374 25342 29426 25394
rect 33854 25342 33906 25394
rect 34638 25342 34690 25394
rect 37774 25342 37826 25394
rect 42590 25342 42642 25394
rect 44158 25342 44210 25394
rect 53342 25342 53394 25394
rect 54462 25342 54514 25394
rect 5630 25230 5682 25282
rect 10334 25230 10386 25282
rect 18734 25230 18786 25282
rect 21982 25230 22034 25282
rect 22654 25230 22706 25282
rect 23102 25230 23154 25282
rect 25342 25230 25394 25282
rect 44270 25230 44322 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 7758 24894 7810 24946
rect 13022 24894 13074 24946
rect 15486 24894 15538 24946
rect 20638 24894 20690 24946
rect 20750 24894 20802 24946
rect 22318 24894 22370 24946
rect 22766 24894 22818 24946
rect 24670 24894 24722 24946
rect 26350 24894 26402 24946
rect 28478 24894 28530 24946
rect 29374 24894 29426 24946
rect 32510 24894 32562 24946
rect 32622 24894 32674 24946
rect 36990 24894 37042 24946
rect 41694 24894 41746 24946
rect 49534 24894 49586 24946
rect 4958 24782 5010 24834
rect 8094 24782 8146 24834
rect 8878 24782 8930 24834
rect 10446 24782 10498 24834
rect 18510 24782 18562 24834
rect 20862 24782 20914 24834
rect 23102 24782 23154 24834
rect 23550 24782 23602 24834
rect 23662 24782 23714 24834
rect 26686 24782 26738 24834
rect 28142 24782 28194 24834
rect 32062 24782 32114 24834
rect 33070 24782 33122 24834
rect 35422 24782 35474 24834
rect 35646 24782 35698 24834
rect 37438 24782 37490 24834
rect 38894 24782 38946 24834
rect 42702 24782 42754 24834
rect 47182 24782 47234 24834
rect 47518 24782 47570 24834
rect 48974 24782 49026 24834
rect 51102 24782 51154 24834
rect 52670 24782 52722 24834
rect 4286 24670 4338 24722
rect 9662 24670 9714 24722
rect 15822 24670 15874 24722
rect 16270 24670 16322 24722
rect 18174 24670 18226 24722
rect 19070 24670 19122 24722
rect 19630 24670 19682 24722
rect 21646 24670 21698 24722
rect 25566 24670 25618 24722
rect 32286 24670 32338 24722
rect 33854 24670 33906 24722
rect 34078 24670 34130 24722
rect 36206 24670 36258 24722
rect 40014 24670 40066 24722
rect 41022 24670 41074 24722
rect 41134 24670 41186 24722
rect 41246 24670 41298 24722
rect 43486 24670 43538 24722
rect 43934 24670 43986 24722
rect 45390 24670 45442 24722
rect 46510 24670 46562 24722
rect 47854 24670 47906 24722
rect 48190 24670 48242 24722
rect 49198 24670 49250 24722
rect 49534 24670 49586 24722
rect 49870 24670 49922 24722
rect 51326 24670 51378 24722
rect 51998 24670 52050 24722
rect 7086 24558 7138 24610
rect 12574 24558 12626 24610
rect 17838 24558 17890 24610
rect 19182 24558 19234 24610
rect 20078 24558 20130 24610
rect 21310 24558 21362 24610
rect 24222 24558 24274 24610
rect 25230 24558 25282 24610
rect 25790 24558 25842 24610
rect 28926 24558 28978 24610
rect 42478 24558 42530 24610
rect 46734 24558 46786 24610
rect 47966 24558 48018 24610
rect 50206 24558 50258 24610
rect 54798 24558 54850 24610
rect 8990 24446 9042 24498
rect 22094 24446 22146 24498
rect 22430 24446 22482 24498
rect 23662 24446 23714 24498
rect 35758 24446 35810 24498
rect 49422 24446 49474 24498
rect 50430 24446 50482 24498
rect 50766 24446 50818 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 11230 24110 11282 24162
rect 11566 24110 11618 24162
rect 14926 24110 14978 24162
rect 35422 24110 35474 24162
rect 43934 24110 43986 24162
rect 47182 24110 47234 24162
rect 49198 24110 49250 24162
rect 7422 23998 7474 24050
rect 8318 23998 8370 24050
rect 8654 23998 8706 24050
rect 9214 23998 9266 24050
rect 23550 23998 23602 24050
rect 29150 23998 29202 24050
rect 32510 23998 32562 24050
rect 33630 23998 33682 24050
rect 34078 23998 34130 24050
rect 34190 23998 34242 24050
rect 36318 23998 36370 24050
rect 37326 23998 37378 24050
rect 43710 23998 43762 24050
rect 53230 23998 53282 24050
rect 53678 23998 53730 24050
rect 7982 23886 8034 23938
rect 12126 23886 12178 23938
rect 17278 23886 17330 23938
rect 17502 23886 17554 23938
rect 19630 23886 19682 23938
rect 19966 23886 20018 23938
rect 21982 23886 22034 23938
rect 22542 23886 22594 23938
rect 23102 23886 23154 23938
rect 24894 23886 24946 23938
rect 25566 23886 25618 23938
rect 32062 23886 32114 23938
rect 33182 23886 33234 23938
rect 35198 23886 35250 23938
rect 35646 23886 35698 23938
rect 37214 23886 37266 23938
rect 37886 23886 37938 23938
rect 38334 23886 38386 23938
rect 40014 23886 40066 23938
rect 41694 23886 41746 23938
rect 42030 23886 42082 23938
rect 44942 23886 44994 23938
rect 45166 23886 45218 23938
rect 45390 23886 45442 23938
rect 45614 23886 45666 23938
rect 45950 23886 46002 23938
rect 46174 23886 46226 23938
rect 46734 23886 46786 23938
rect 47966 23886 48018 23938
rect 50430 23886 50482 23938
rect 50878 23886 50930 23938
rect 51214 23886 51266 23938
rect 51438 23886 51490 23938
rect 4622 23774 4674 23826
rect 7758 23774 7810 23826
rect 12238 23774 12290 23826
rect 15150 23774 15202 23826
rect 15486 23774 15538 23826
rect 17614 23774 17666 23826
rect 17838 23774 17890 23826
rect 18734 23774 18786 23826
rect 21534 23774 21586 23826
rect 23998 23774 24050 23826
rect 31278 23774 31330 23826
rect 33406 23774 33458 23826
rect 33742 23774 33794 23826
rect 34302 23774 34354 23826
rect 34974 23774 35026 23826
rect 35870 23774 35922 23826
rect 37438 23774 37490 23826
rect 39902 23774 39954 23826
rect 41134 23774 41186 23826
rect 42142 23774 42194 23826
rect 42590 23774 42642 23826
rect 46510 23774 46562 23826
rect 47630 23774 47682 23826
rect 47742 23774 47794 23826
rect 48750 23774 48802 23826
rect 49422 23774 49474 23826
rect 50990 23774 51042 23826
rect 51662 23774 51714 23826
rect 51886 23774 51938 23826
rect 52782 23774 52834 23826
rect 4286 23662 4338 23714
rect 6414 23662 6466 23714
rect 8766 23662 8818 23714
rect 13806 23662 13858 23714
rect 14254 23662 14306 23714
rect 14590 23662 14642 23714
rect 16830 23662 16882 23714
rect 18286 23662 18338 23714
rect 22878 23662 22930 23714
rect 22990 23662 23042 23714
rect 35982 23662 36034 23714
rect 43038 23662 43090 23714
rect 44270 23662 44322 23714
rect 45502 23662 45554 23714
rect 46398 23662 46450 23714
rect 48302 23662 48354 23714
rect 48414 23662 48466 23714
rect 48526 23662 48578 23714
rect 49310 23662 49362 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 6526 23326 6578 23378
rect 12910 23326 12962 23378
rect 17726 23326 17778 23378
rect 17950 23326 18002 23378
rect 24446 23326 24498 23378
rect 29374 23326 29426 23378
rect 33966 23326 34018 23378
rect 34302 23326 34354 23378
rect 34526 23326 34578 23378
rect 38558 23326 38610 23378
rect 41806 23326 41858 23378
rect 49198 23326 49250 23378
rect 50878 23326 50930 23378
rect 51886 23326 51938 23378
rect 52334 23326 52386 23378
rect 2382 23214 2434 23266
rect 3950 23214 4002 23266
rect 7422 23214 7474 23266
rect 20078 23214 20130 23266
rect 22206 23214 22258 23266
rect 23102 23214 23154 23266
rect 24334 23214 24386 23266
rect 34190 23214 34242 23266
rect 34750 23214 34802 23266
rect 36430 23214 36482 23266
rect 38782 23214 38834 23266
rect 39678 23214 39730 23266
rect 39790 23214 39842 23266
rect 42590 23214 42642 23266
rect 46062 23214 46114 23266
rect 46510 23214 46562 23266
rect 47518 23214 47570 23266
rect 49646 23214 49698 23266
rect 50766 23214 50818 23266
rect 52446 23214 52498 23266
rect 53006 23214 53058 23266
rect 2718 23102 2770 23154
rect 3278 23102 3330 23154
rect 7646 23102 7698 23154
rect 9662 23102 9714 23154
rect 13246 23102 13298 23154
rect 13806 23102 13858 23154
rect 18062 23102 18114 23154
rect 18622 23102 18674 23154
rect 20750 23102 20802 23154
rect 22654 23102 22706 23154
rect 24670 23102 24722 23154
rect 28590 23102 28642 23154
rect 29150 23102 29202 23154
rect 35086 23102 35138 23154
rect 35646 23102 35698 23154
rect 36542 23102 36594 23154
rect 37774 23102 37826 23154
rect 39006 23102 39058 23154
rect 39454 23102 39506 23154
rect 40238 23102 40290 23154
rect 43598 23102 43650 23154
rect 43822 23102 43874 23154
rect 45390 23102 45442 23154
rect 46286 23102 46338 23154
rect 47070 23102 47122 23154
rect 47966 23102 48018 23154
rect 48638 23102 48690 23154
rect 49086 23102 49138 23154
rect 49310 23102 49362 23154
rect 50094 23102 50146 23154
rect 50542 23102 50594 23154
rect 51326 23102 51378 23154
rect 6078 22990 6130 23042
rect 12574 22990 12626 23042
rect 13470 22990 13522 23042
rect 14590 22990 14642 23042
rect 16718 22990 16770 23042
rect 19854 22990 19906 23042
rect 23438 22990 23490 23042
rect 25342 22990 25394 23042
rect 25678 22990 25730 23042
rect 27806 22990 27858 23042
rect 42142 22990 42194 23042
rect 46174 22990 46226 23042
rect 47406 22990 47458 23042
rect 49758 22990 49810 23042
rect 49982 22990 50034 23042
rect 51774 22990 51826 23042
rect 6862 22878 6914 22930
rect 18510 22878 18562 22930
rect 19630 22878 19682 22930
rect 40462 22878 40514 22930
rect 51102 22878 51154 22930
rect 51662 22878 51714 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 5742 22542 5794 22594
rect 8654 22542 8706 22594
rect 13582 22542 13634 22594
rect 15150 22542 15202 22594
rect 25790 22542 25842 22594
rect 29262 22542 29314 22594
rect 29598 22542 29650 22594
rect 36094 22542 36146 22594
rect 38222 22542 38274 22594
rect 38334 22542 38386 22594
rect 38558 22542 38610 22594
rect 38670 22542 38722 22594
rect 40910 22542 40962 22594
rect 44830 22542 44882 22594
rect 48750 22542 48802 22594
rect 50990 22542 51042 22594
rect 51662 22542 51714 22594
rect 2494 22430 2546 22482
rect 4622 22430 4674 22482
rect 12574 22430 12626 22482
rect 19182 22430 19234 22482
rect 23102 22430 23154 22482
rect 24446 22430 24498 22482
rect 24894 22430 24946 22482
rect 34190 22430 34242 22482
rect 36206 22430 36258 22482
rect 37102 22430 37154 22482
rect 37326 22430 37378 22482
rect 39118 22430 39170 22482
rect 40126 22430 40178 22482
rect 40574 22430 40626 22482
rect 42030 22430 42082 22482
rect 46510 22430 46562 22482
rect 48078 22430 48130 22482
rect 49870 22430 49922 22482
rect 51214 22430 51266 22482
rect 52110 22430 52162 22482
rect 1822 22318 1874 22370
rect 6078 22318 6130 22370
rect 6862 22318 6914 22370
rect 7646 22318 7698 22370
rect 7982 22318 8034 22370
rect 8990 22318 9042 22370
rect 9662 22318 9714 22370
rect 14142 22318 14194 22370
rect 18734 22318 18786 22370
rect 20638 22318 20690 22370
rect 22766 22318 22818 22370
rect 24782 22318 24834 22370
rect 25566 22318 25618 22370
rect 27694 22318 27746 22370
rect 28478 22318 28530 22370
rect 33294 22318 33346 22370
rect 36430 22318 36482 22370
rect 39790 22318 39842 22370
rect 40686 22318 40738 22370
rect 42590 22318 42642 22370
rect 42814 22318 42866 22370
rect 46062 22318 46114 22370
rect 47518 22318 47570 22370
rect 47854 22318 47906 22370
rect 48414 22318 48466 22370
rect 50766 22318 50818 22370
rect 51662 22318 51714 22370
rect 6750 22206 6802 22258
rect 10446 22206 10498 22258
rect 13582 22206 13634 22258
rect 5070 22094 5122 22146
rect 7534 22094 7586 22146
rect 7870 22094 7922 22146
rect 8766 22094 8818 22146
rect 13694 22150 13746 22202
rect 14366 22206 14418 22258
rect 15374 22206 15426 22258
rect 15934 22206 15986 22258
rect 18174 22206 18226 22258
rect 19070 22206 19122 22258
rect 21870 22206 21922 22258
rect 26686 22206 26738 22258
rect 26798 22206 26850 22258
rect 27022 22206 27074 22258
rect 28254 22206 28306 22258
rect 29822 22206 29874 22258
rect 30382 22206 30434 22258
rect 43374 22206 43426 22258
rect 45278 22206 45330 22258
rect 45390 22206 45442 22258
rect 45502 22206 45554 22258
rect 49422 22206 49474 22258
rect 49758 22206 49810 22258
rect 49982 22206 50034 22258
rect 50430 22206 50482 22258
rect 14814 22094 14866 22146
rect 23326 22094 23378 22146
rect 26126 22094 26178 22146
rect 27358 22094 27410 22146
rect 37774 22094 37826 22146
rect 48638 22094 48690 22146
rect 49086 22094 49138 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 8990 21758 9042 21810
rect 10894 21758 10946 21810
rect 27134 21758 27186 21810
rect 29710 21758 29762 21810
rect 30494 21758 30546 21810
rect 35534 21758 35586 21810
rect 38894 21758 38946 21810
rect 47630 21758 47682 21810
rect 48750 21758 48802 21810
rect 49534 21758 49586 21810
rect 7534 21646 7586 21698
rect 7758 21646 7810 21698
rect 8206 21646 8258 21698
rect 9550 21646 9602 21698
rect 11230 21646 11282 21698
rect 11902 21646 11954 21698
rect 12798 21646 12850 21698
rect 14478 21646 14530 21698
rect 19854 21646 19906 21698
rect 19966 21646 20018 21698
rect 21982 21646 22034 21698
rect 23214 21646 23266 21698
rect 23998 21646 24050 21698
rect 24670 21646 24722 21698
rect 25230 21646 25282 21698
rect 26462 21646 26514 21698
rect 29150 21646 29202 21698
rect 30046 21646 30098 21698
rect 31950 21646 32002 21698
rect 33742 21646 33794 21698
rect 34078 21646 34130 21698
rect 34750 21646 34802 21698
rect 36654 21646 36706 21698
rect 41022 21646 41074 21698
rect 46062 21646 46114 21698
rect 47406 21646 47458 21698
rect 50990 21646 51042 21698
rect 1822 21534 1874 21586
rect 8542 21534 8594 21586
rect 8878 21534 8930 21586
rect 9774 21534 9826 21586
rect 9998 21534 10050 21586
rect 10110 21534 10162 21586
rect 12238 21534 12290 21586
rect 12910 21534 12962 21586
rect 13918 21534 13970 21586
rect 14702 21534 14754 21586
rect 16158 21534 16210 21586
rect 16718 21534 16770 21586
rect 20190 21534 20242 21586
rect 20526 21534 20578 21586
rect 20862 21534 20914 21586
rect 22206 21534 22258 21586
rect 22990 21534 23042 21586
rect 23550 21534 23602 21586
rect 24558 21534 24610 21586
rect 25454 21534 25506 21586
rect 26910 21534 26962 21586
rect 32286 21534 32338 21586
rect 33182 21534 33234 21586
rect 35086 21534 35138 21586
rect 35870 21534 35922 21586
rect 39902 21534 39954 21586
rect 40126 21534 40178 21586
rect 40462 21534 40514 21586
rect 42030 21534 42082 21586
rect 43038 21534 43090 21586
rect 46846 21534 46898 21586
rect 47294 21534 47346 21586
rect 47854 21534 47906 21586
rect 48974 21534 49026 21586
rect 49646 21534 49698 21586
rect 50206 21534 50258 21586
rect 2494 21422 2546 21474
rect 4622 21422 4674 21474
rect 5070 21422 5122 21474
rect 7870 21422 7922 21474
rect 8654 21422 8706 21474
rect 9662 21422 9714 21474
rect 15262 21422 15314 21474
rect 17502 21422 17554 21474
rect 18510 21422 18562 21474
rect 26350 21422 26402 21474
rect 40238 21422 40290 21474
rect 42142 21422 42194 21474
rect 43486 21422 43538 21474
rect 43934 21422 43986 21474
rect 48302 21422 48354 21474
rect 53118 21422 53170 21474
rect 13582 21310 13634 21362
rect 20638 21310 20690 21362
rect 21310 21310 21362 21362
rect 22542 21310 22594 21362
rect 23662 21310 23714 21362
rect 25790 21310 25842 21362
rect 29038 21310 29090 21362
rect 33518 21310 33570 21362
rect 49534 21310 49586 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 4174 20974 4226 21026
rect 7646 20974 7698 21026
rect 7982 20974 8034 21026
rect 8542 20974 8594 21026
rect 11790 20974 11842 21026
rect 12350 20974 12402 21026
rect 14366 20974 14418 21026
rect 18958 20974 19010 21026
rect 20526 20974 20578 21026
rect 21646 20974 21698 21026
rect 23326 20974 23378 21026
rect 35086 20974 35138 21026
rect 41806 20974 41858 21026
rect 11230 20862 11282 20914
rect 20414 20862 20466 20914
rect 24222 20862 24274 20914
rect 25006 20862 25058 20914
rect 26350 20862 26402 20914
rect 27470 20862 27522 20914
rect 28590 20862 28642 20914
rect 31838 20862 31890 20914
rect 33966 20862 34018 20914
rect 37214 20862 37266 20914
rect 41246 20862 41298 20914
rect 42814 20862 42866 20914
rect 44046 20862 44098 20914
rect 44270 20862 44322 20914
rect 45614 20862 45666 20914
rect 47742 20862 47794 20914
rect 48302 20862 48354 20914
rect 48638 20862 48690 20914
rect 49870 20862 49922 20914
rect 4958 20750 5010 20802
rect 7982 20750 8034 20802
rect 8542 20750 8594 20802
rect 9102 20750 9154 20802
rect 12350 20750 12402 20802
rect 12910 20750 12962 20802
rect 14366 20750 14418 20802
rect 14926 20750 14978 20802
rect 15598 20750 15650 20802
rect 17390 20750 17442 20802
rect 18062 20750 18114 20802
rect 21534 20750 21586 20802
rect 21758 20750 21810 20802
rect 22318 20750 22370 20802
rect 24558 20750 24610 20802
rect 25678 20750 25730 20802
rect 29150 20750 29202 20802
rect 30718 20750 30770 20802
rect 31054 20750 31106 20802
rect 35422 20750 35474 20802
rect 38446 20750 38498 20802
rect 41582 20750 41634 20802
rect 42030 20750 42082 20802
rect 42366 20750 42418 20802
rect 44942 20750 44994 20802
rect 2382 20638 2434 20690
rect 2718 20638 2770 20690
rect 3838 20638 3890 20690
rect 4734 20638 4786 20690
rect 5966 20638 6018 20690
rect 8878 20638 8930 20690
rect 11566 20638 11618 20690
rect 12686 20638 12738 20690
rect 14702 20638 14754 20690
rect 15262 20638 15314 20690
rect 19182 20638 19234 20690
rect 21310 20638 21362 20690
rect 23214 20638 23266 20690
rect 25454 20638 25506 20690
rect 27022 20638 27074 20690
rect 35646 20638 35698 20690
rect 35982 20638 36034 20690
rect 39118 20638 39170 20690
rect 5630 20526 5682 20578
rect 8990 20526 9042 20578
rect 11678 20526 11730 20578
rect 12798 20526 12850 20578
rect 14814 20526 14866 20578
rect 17614 20526 17666 20578
rect 18286 20526 18338 20578
rect 18622 20526 18674 20578
rect 21982 20526 22034 20578
rect 22206 20526 22258 20578
rect 22766 20526 22818 20578
rect 23774 20526 23826 20578
rect 26686 20526 26738 20578
rect 29486 20526 29538 20578
rect 41582 20526 41634 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 17838 20190 17890 20242
rect 23214 20190 23266 20242
rect 41134 20190 41186 20242
rect 45838 20190 45890 20242
rect 47182 20190 47234 20242
rect 5518 20078 5570 20130
rect 9774 20078 9826 20130
rect 16382 20078 16434 20130
rect 18286 20078 18338 20130
rect 19966 20078 20018 20130
rect 20862 20078 20914 20130
rect 21310 20078 21362 20130
rect 22430 20078 22482 20130
rect 23102 20078 23154 20130
rect 23774 20078 23826 20130
rect 26350 20078 26402 20130
rect 28926 20078 28978 20130
rect 29486 20078 29538 20130
rect 30046 20078 30098 20130
rect 30830 20078 30882 20130
rect 33070 20078 33122 20130
rect 34974 20078 35026 20130
rect 41582 20078 41634 20130
rect 41694 20078 41746 20130
rect 4846 19966 4898 20018
rect 11902 19966 11954 20018
rect 14366 19966 14418 20018
rect 14926 19966 14978 20018
rect 15038 19966 15090 20018
rect 15150 19966 15202 20018
rect 15486 19966 15538 20018
rect 15710 19966 15762 20018
rect 16606 19966 16658 20018
rect 18622 19966 18674 20018
rect 19070 19966 19122 20018
rect 20190 19966 20242 20018
rect 22654 19966 22706 20018
rect 23438 19966 23490 20018
rect 25566 19966 25618 20018
rect 30606 19966 30658 20018
rect 33406 19966 33458 20018
rect 34302 19966 34354 20018
rect 37438 19966 37490 20018
rect 7646 19854 7698 19906
rect 8094 19854 8146 19906
rect 8766 19854 8818 19906
rect 9550 19854 9602 19906
rect 21982 19854 22034 19906
rect 24670 19854 24722 19906
rect 28478 19854 28530 19906
rect 37102 19854 37154 19906
rect 39790 19854 39842 19906
rect 42142 19854 42194 19906
rect 9886 19742 9938 19794
rect 11566 19742 11618 19794
rect 11902 19742 11954 19794
rect 14590 19742 14642 19794
rect 15934 19742 15986 19794
rect 16046 19742 16098 19794
rect 19406 19742 19458 19794
rect 21646 19742 21698 19794
rect 29262 19742 29314 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 6526 19406 6578 19458
rect 6862 19406 6914 19458
rect 10334 19406 10386 19458
rect 14926 19406 14978 19458
rect 16718 19406 16770 19458
rect 30718 19406 30770 19458
rect 18286 19294 18338 19346
rect 20414 19294 20466 19346
rect 24222 19294 24274 19346
rect 25454 19294 25506 19346
rect 32510 19294 32562 19346
rect 34638 19294 34690 19346
rect 37102 19294 37154 19346
rect 7646 19182 7698 19234
rect 9326 19182 9378 19234
rect 10222 19182 10274 19234
rect 10670 19182 10722 19234
rect 11566 19182 11618 19234
rect 11902 19182 11954 19234
rect 14478 19182 14530 19234
rect 14702 19182 14754 19234
rect 15038 19182 15090 19234
rect 15710 19182 15762 19234
rect 16158 19182 16210 19234
rect 16494 19182 16546 19234
rect 17502 19182 17554 19234
rect 21310 19182 21362 19234
rect 25006 19182 25058 19234
rect 26014 19182 26066 19234
rect 26462 19182 26514 19234
rect 29710 19182 29762 19234
rect 30382 19182 30434 19234
rect 31838 19182 31890 19234
rect 35310 19182 35362 19234
rect 35982 19182 36034 19234
rect 2830 19070 2882 19122
rect 3614 19070 3666 19122
rect 7422 19070 7474 19122
rect 8206 19070 8258 19122
rect 8318 19070 8370 19122
rect 8990 19070 9042 19122
rect 9886 19070 9938 19122
rect 11118 19070 11170 19122
rect 11342 19070 11394 19122
rect 22094 19070 22146 19122
rect 25678 19070 25730 19122
rect 26798 19070 26850 19122
rect 29822 19070 29874 19122
rect 35422 19070 35474 19122
rect 2494 18958 2546 19010
rect 3278 18958 3330 19010
rect 5742 18958 5794 19010
rect 7982 18958 8034 19010
rect 9102 18958 9154 19010
rect 10110 18958 10162 19010
rect 11902 18958 11954 19010
rect 24670 18958 24722 19010
rect 27022 18958 27074 19010
rect 36318 18958 36370 19010
rect 37550 18958 37602 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 8654 18622 8706 18674
rect 11454 18622 11506 18674
rect 14142 18622 14194 18674
rect 16382 18622 16434 18674
rect 25566 18622 25618 18674
rect 26350 18622 26402 18674
rect 38670 18622 38722 18674
rect 3054 18510 3106 18562
rect 6526 18510 6578 18562
rect 9550 18510 9602 18562
rect 11230 18510 11282 18562
rect 12910 18510 12962 18562
rect 13582 18510 13634 18562
rect 20862 18510 20914 18562
rect 27246 18510 27298 18562
rect 27694 18510 27746 18562
rect 27918 18510 27970 18562
rect 31054 18510 31106 18562
rect 33742 18510 33794 18562
rect 34078 18510 34130 18562
rect 2270 18398 2322 18450
rect 5630 18398 5682 18450
rect 5966 18398 6018 18450
rect 6638 18398 6690 18450
rect 8430 18398 8482 18450
rect 8990 18398 9042 18450
rect 9886 18398 9938 18450
rect 9998 18398 10050 18450
rect 10334 18398 10386 18450
rect 11006 18398 11058 18450
rect 11566 18398 11618 18450
rect 12350 18398 12402 18450
rect 12798 18398 12850 18450
rect 13022 18398 13074 18450
rect 13358 18398 13410 18450
rect 13806 18398 13858 18450
rect 14142 18398 14194 18450
rect 15934 18398 15986 18450
rect 16158 18398 16210 18450
rect 17390 18398 17442 18450
rect 21198 18398 21250 18450
rect 21646 18398 21698 18450
rect 24334 18398 24386 18450
rect 25454 18398 25506 18450
rect 31838 18398 31890 18450
rect 38222 18398 38274 18450
rect 5182 18286 5234 18338
rect 9662 18286 9714 18338
rect 16046 18286 16098 18338
rect 17950 18286 18002 18338
rect 18398 18286 18450 18338
rect 23774 18286 23826 18338
rect 24110 18286 24162 18338
rect 24670 18286 24722 18338
rect 26798 18286 26850 18338
rect 28926 18286 28978 18338
rect 32286 18286 32338 18338
rect 33182 18286 33234 18338
rect 34862 18286 34914 18338
rect 35310 18286 35362 18338
rect 37438 18286 37490 18338
rect 11566 18174 11618 18226
rect 12462 18174 12514 18226
rect 17502 18174 17554 18226
rect 21198 18174 21250 18226
rect 27582 18174 27634 18226
rect 33518 18174 33570 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 5742 17838 5794 17890
rect 7198 17838 7250 17890
rect 7646 17838 7698 17890
rect 12574 17838 12626 17890
rect 15710 17838 15762 17890
rect 24894 17838 24946 17890
rect 25790 17838 25842 17890
rect 27582 17838 27634 17890
rect 30158 17838 30210 17890
rect 2494 17726 2546 17778
rect 4622 17726 4674 17778
rect 7646 17726 7698 17778
rect 15374 17726 15426 17778
rect 16158 17726 16210 17778
rect 27134 17726 27186 17778
rect 27918 17726 27970 17778
rect 1822 17614 1874 17666
rect 6078 17614 6130 17666
rect 6526 17614 6578 17666
rect 8318 17614 8370 17666
rect 8654 17614 8706 17666
rect 9774 17614 9826 17666
rect 12462 17614 12514 17666
rect 12686 17614 12738 17666
rect 14142 17614 14194 17666
rect 14366 17614 14418 17666
rect 14702 17614 14754 17666
rect 15150 17614 15202 17666
rect 15598 17614 15650 17666
rect 17166 17614 17218 17666
rect 17614 17614 17666 17666
rect 23214 17614 23266 17666
rect 23886 17614 23938 17666
rect 24670 17614 24722 17666
rect 25342 17614 25394 17666
rect 26574 17614 26626 17666
rect 29822 17614 29874 17666
rect 33854 17614 33906 17666
rect 35870 17614 35922 17666
rect 6862 17502 6914 17554
rect 7870 17502 7922 17554
rect 8094 17502 8146 17554
rect 8990 17502 9042 17554
rect 9998 17502 10050 17554
rect 10334 17502 10386 17554
rect 10670 17502 10722 17554
rect 12126 17502 12178 17554
rect 14590 17502 14642 17554
rect 14814 17502 14866 17554
rect 16942 17502 16994 17554
rect 5070 17390 5122 17442
rect 8318 17390 8370 17442
rect 9326 17390 9378 17442
rect 11118 17390 11170 17442
rect 12910 17390 12962 17442
rect 16606 17390 16658 17442
rect 17950 17446 18002 17498
rect 19518 17502 19570 17554
rect 23550 17502 23602 17554
rect 25118 17502 25170 17554
rect 25678 17502 25730 17554
rect 36094 17502 36146 17554
rect 19182 17390 19234 17442
rect 24222 17390 24274 17442
rect 25006 17390 25058 17442
rect 25790 17390 25842 17442
rect 27022 17390 27074 17442
rect 27246 17390 27298 17442
rect 27806 17390 27858 17442
rect 30046 17390 30098 17442
rect 34078 17390 34130 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 6414 17054 6466 17106
rect 6862 17054 6914 17106
rect 7646 17054 7698 17106
rect 8430 17054 8482 17106
rect 8990 17054 9042 17106
rect 9550 17054 9602 17106
rect 9886 17054 9938 17106
rect 10334 17054 10386 17106
rect 11342 17054 11394 17106
rect 16158 17054 16210 17106
rect 21646 17054 21698 17106
rect 25230 17054 25282 17106
rect 26462 17054 26514 17106
rect 27134 17054 27186 17106
rect 27918 17054 27970 17106
rect 36878 17054 36930 17106
rect 2382 16942 2434 16994
rect 8094 16942 8146 16994
rect 14814 16942 14866 16994
rect 15150 16942 15202 16994
rect 15822 16942 15874 16994
rect 16830 16942 16882 16994
rect 17390 16942 17442 16994
rect 19070 16942 19122 16994
rect 21758 16942 21810 16994
rect 23886 16942 23938 16994
rect 26014 16942 26066 16994
rect 27358 16942 27410 16994
rect 28702 16942 28754 16994
rect 30830 16942 30882 16994
rect 31278 16942 31330 16994
rect 31950 16942 32002 16994
rect 32398 16942 32450 16994
rect 34302 16942 34354 16994
rect 2718 16830 2770 16882
rect 6078 16830 6130 16882
rect 6302 16830 6354 16882
rect 6750 16830 6802 16882
rect 11790 16830 11842 16882
rect 12798 16830 12850 16882
rect 13022 16830 13074 16882
rect 13582 16830 13634 16882
rect 14478 16830 14530 16882
rect 15486 16830 15538 16882
rect 16606 16830 16658 16882
rect 17614 16830 17666 16882
rect 18286 16830 18338 16882
rect 21422 16830 21474 16882
rect 22654 16830 22706 16882
rect 25230 16830 25282 16882
rect 25790 16830 25842 16882
rect 26910 16830 26962 16882
rect 27582 16830 27634 16882
rect 28030 16830 28082 16882
rect 28366 16830 28418 16882
rect 30606 16830 30658 16882
rect 33630 16830 33682 16882
rect 7422 16718 7474 16770
rect 7758 16718 7810 16770
rect 10894 16718 10946 16770
rect 11230 16718 11282 16770
rect 12910 16718 12962 16770
rect 13246 16718 13298 16770
rect 14702 16718 14754 16770
rect 21198 16718 21250 16770
rect 27134 16718 27186 16770
rect 36430 16718 36482 16770
rect 14366 16606 14418 16658
rect 25566 16606 25618 16658
rect 28142 16606 28194 16658
rect 31614 16606 31666 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 5742 16270 5794 16322
rect 6078 16270 6130 16322
rect 19518 16270 19570 16322
rect 19854 16270 19906 16322
rect 28142 16270 28194 16322
rect 29598 16270 29650 16322
rect 34190 16270 34242 16322
rect 2494 16158 2546 16210
rect 4622 16158 4674 16210
rect 11118 16158 11170 16210
rect 16046 16158 16098 16210
rect 21534 16158 21586 16210
rect 24222 16158 24274 16210
rect 26238 16158 26290 16210
rect 30830 16158 30882 16210
rect 32958 16158 33010 16210
rect 1822 16046 1874 16098
rect 6862 16046 6914 16098
rect 8206 16046 8258 16098
rect 11902 16046 11954 16098
rect 14254 16046 14306 16098
rect 14814 16046 14866 16098
rect 16382 16046 16434 16098
rect 17502 16046 17554 16098
rect 18062 16046 18114 16098
rect 19070 16046 19122 16098
rect 20526 16046 20578 16098
rect 22766 16046 22818 16098
rect 23438 16046 23490 16098
rect 24334 16046 24386 16098
rect 25678 16046 25730 16098
rect 26686 16046 26738 16098
rect 27022 16046 27074 16098
rect 27246 16046 27298 16098
rect 27918 16046 27970 16098
rect 33630 16046 33682 16098
rect 34526 16046 34578 16098
rect 35870 16046 35922 16098
rect 6750 15934 6802 15986
rect 7422 15934 7474 15986
rect 7646 15934 7698 15986
rect 7758 15934 7810 15986
rect 8990 15934 9042 15986
rect 12238 15934 12290 15986
rect 12462 15934 12514 15986
rect 13918 15934 13970 15986
rect 14590 15934 14642 15986
rect 15262 15934 15314 15986
rect 15598 15934 15650 15986
rect 16718 15934 16770 15986
rect 18286 15934 18338 15986
rect 20414 15934 20466 15986
rect 24558 15934 24610 15986
rect 27470 15934 27522 15986
rect 28366 15934 28418 15986
rect 28590 15934 28642 15986
rect 29822 15934 29874 15986
rect 30382 15934 30434 15986
rect 34750 15934 34802 15986
rect 35086 15934 35138 15986
rect 5070 15822 5122 15874
rect 11566 15822 11618 15874
rect 15934 15822 15986 15874
rect 17166 15822 17218 15874
rect 18734 15822 18786 15874
rect 21982 15822 22034 15874
rect 23102 15822 23154 15874
rect 23774 15822 23826 15874
rect 24110 15822 24162 15874
rect 25006 15822 25058 15874
rect 25342 15822 25394 15874
rect 26126 15822 26178 15874
rect 26350 15822 26402 15874
rect 26686 15822 26738 15874
rect 28142 15822 28194 15874
rect 29262 15822 29314 15874
rect 36094 15822 36146 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 12574 15486 12626 15538
rect 12798 15486 12850 15538
rect 13470 15486 13522 15538
rect 14478 15486 14530 15538
rect 14926 15486 14978 15538
rect 17838 15486 17890 15538
rect 19406 15486 19458 15538
rect 23326 15486 23378 15538
rect 23662 15486 23714 15538
rect 24222 15486 24274 15538
rect 24446 15486 24498 15538
rect 25342 15486 25394 15538
rect 25566 15486 25618 15538
rect 26686 15486 26738 15538
rect 28254 15486 28306 15538
rect 30942 15486 30994 15538
rect 33406 15486 33458 15538
rect 33854 15486 33906 15538
rect 38782 15486 38834 15538
rect 10334 15374 10386 15426
rect 12014 15374 12066 15426
rect 20078 15374 20130 15426
rect 20526 15374 20578 15426
rect 25790 15374 25842 15426
rect 27470 15374 27522 15426
rect 28030 15374 28082 15426
rect 31502 15374 31554 15426
rect 31838 15374 31890 15426
rect 34862 15374 34914 15426
rect 37550 15374 37602 15426
rect 2942 15262 2994 15314
rect 6974 15262 7026 15314
rect 10446 15262 10498 15314
rect 11454 15262 11506 15314
rect 12238 15262 12290 15314
rect 12910 15262 12962 15314
rect 19854 15262 19906 15314
rect 20638 15262 20690 15314
rect 21646 15262 21698 15314
rect 24558 15262 24610 15314
rect 24670 15262 24722 15314
rect 25230 15262 25282 15314
rect 26350 15262 26402 15314
rect 26686 15262 26738 15314
rect 27134 15262 27186 15314
rect 27806 15262 27858 15314
rect 28254 15262 28306 15314
rect 28366 15262 28418 15314
rect 34974 15262 35026 15314
rect 38334 15262 38386 15314
rect 3614 15150 3666 15202
rect 5742 15150 5794 15202
rect 8206 15150 8258 15202
rect 9774 15150 9826 15202
rect 13918 15150 13970 15202
rect 15598 15150 15650 15202
rect 31278 15150 31330 15202
rect 34190 15150 34242 15202
rect 35422 15150 35474 15202
rect 11118 15038 11170 15090
rect 21310 15038 21362 15090
rect 26910 15038 26962 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 11006 14702 11058 14754
rect 11678 14702 11730 14754
rect 15150 14702 15202 14754
rect 26798 14702 26850 14754
rect 27358 14702 27410 14754
rect 36206 14702 36258 14754
rect 9886 14590 9938 14642
rect 10894 14590 10946 14642
rect 15374 14590 15426 14642
rect 22094 14590 22146 14642
rect 24222 14590 24274 14642
rect 24670 14590 24722 14642
rect 5966 14478 6018 14530
rect 7086 14478 7138 14530
rect 12014 14478 12066 14530
rect 13806 14478 13858 14530
rect 16494 14478 16546 14530
rect 16830 14478 16882 14530
rect 21422 14478 21474 14530
rect 25006 14478 25058 14530
rect 26126 14478 26178 14530
rect 26350 14478 26402 14530
rect 27694 14478 27746 14530
rect 28366 14478 28418 14530
rect 30382 14478 30434 14530
rect 35870 14478 35922 14530
rect 3838 14366 3890 14418
rect 4174 14366 4226 14418
rect 7758 14366 7810 14418
rect 10222 14366 10274 14418
rect 10558 14366 10610 14418
rect 12238 14366 12290 14418
rect 12574 14366 12626 14418
rect 14142 14366 14194 14418
rect 15934 14366 15986 14418
rect 25566 14366 25618 14418
rect 28478 14366 28530 14418
rect 35086 14366 35138 14418
rect 35534 14366 35586 14418
rect 13582 14254 13634 14306
rect 14814 14254 14866 14306
rect 17166 14254 17218 14306
rect 30606 14254 30658 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 6190 13918 6242 13970
rect 7982 13918 8034 13970
rect 9102 13918 9154 13970
rect 12798 13918 12850 13970
rect 13470 13918 13522 13970
rect 13806 13918 13858 13970
rect 15934 13918 15986 13970
rect 25342 13918 25394 13970
rect 26574 13918 26626 13970
rect 27134 13918 27186 13970
rect 3054 13806 3106 13858
rect 3726 13806 3778 13858
rect 7198 13806 7250 13858
rect 8318 13806 8370 13858
rect 12910 13806 12962 13858
rect 14478 13806 14530 13858
rect 14702 13806 14754 13858
rect 17390 13806 17442 13858
rect 19182 13806 19234 13858
rect 27694 13806 27746 13858
rect 31726 13806 31778 13858
rect 34302 13806 34354 13858
rect 3278 13694 3330 13746
rect 4062 13694 4114 13746
rect 6526 13694 6578 13746
rect 7310 13694 7362 13746
rect 9998 13694 10050 13746
rect 17726 13694 17778 13746
rect 19406 13694 19458 13746
rect 20862 13694 20914 13746
rect 21198 13694 21250 13746
rect 26014 13694 26066 13746
rect 26462 13694 26514 13746
rect 26798 13694 26850 13746
rect 27134 13694 27186 13746
rect 27918 13694 27970 13746
rect 32510 13694 32562 13746
rect 33182 13694 33234 13746
rect 33518 13694 33570 13746
rect 33966 13694 34018 13746
rect 5294 13582 5346 13634
rect 10670 13582 10722 13634
rect 18286 13582 18338 13634
rect 22318 13582 22370 13634
rect 24446 13582 24498 13634
rect 27470 13582 27522 13634
rect 29598 13582 29650 13634
rect 12798 13470 12850 13522
rect 14142 13470 14194 13522
rect 18622 13470 18674 13522
rect 20526 13470 20578 13522
rect 20862 13470 20914 13522
rect 26350 13470 26402 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 5742 13134 5794 13186
rect 19742 13134 19794 13186
rect 22094 13134 22146 13186
rect 22990 13134 23042 13186
rect 25566 13134 25618 13186
rect 27358 13134 27410 13186
rect 27918 13134 27970 13186
rect 30382 13134 30434 13186
rect 35198 13134 35250 13186
rect 35534 13134 35586 13186
rect 2830 13022 2882 13074
rect 4958 13022 5010 13074
rect 8542 13022 8594 13074
rect 11678 13022 11730 13074
rect 12462 13022 12514 13074
rect 19406 13022 19458 13074
rect 23438 13022 23490 13074
rect 26238 13022 26290 13074
rect 26910 13022 26962 13074
rect 32734 13022 32786 13074
rect 2046 12910 2098 12962
rect 6078 12910 6130 12962
rect 8878 12910 8930 12962
rect 13918 12910 13970 12962
rect 16606 12910 16658 12962
rect 20078 12910 20130 12962
rect 21982 12910 22034 12962
rect 22318 12910 22370 12962
rect 22766 12910 22818 12962
rect 23326 12910 23378 12962
rect 24222 12910 24274 12962
rect 24334 12910 24386 12962
rect 24446 12910 24498 12962
rect 25118 12910 25170 12962
rect 25342 12910 25394 12962
rect 25678 12910 25730 12962
rect 26462 12910 26514 12962
rect 27358 12910 27410 12962
rect 29374 12910 29426 12962
rect 29598 12910 29650 12962
rect 29710 12910 29762 12962
rect 30718 12910 30770 12962
rect 31502 12910 31554 12962
rect 33182 12910 33234 12962
rect 6414 12798 6466 12850
rect 6862 12798 6914 12850
rect 9550 12798 9602 12850
rect 14142 12798 14194 12850
rect 14478 12798 14530 12850
rect 17278 12798 17330 12850
rect 20302 12798 20354 12850
rect 21646 12798 21698 12850
rect 23550 12798 23602 12850
rect 23886 12798 23938 12850
rect 25006 12798 25058 12850
rect 26126 12798 26178 12850
rect 26798 12798 26850 12850
rect 27022 12798 27074 12850
rect 28030 12798 28082 12850
rect 28254 12798 28306 12850
rect 29150 12798 29202 12850
rect 31278 12798 31330 12850
rect 35758 12798 35810 12850
rect 36318 12798 36370 12850
rect 12798 12686 12850 12738
rect 13582 12686 13634 12738
rect 20750 12686 20802 12738
rect 22430 12686 22482 12738
rect 24670 12686 24722 12738
rect 29934 12686 29986 12738
rect 33406 12686 33458 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 5070 12350 5122 12402
rect 9886 12350 9938 12402
rect 16830 12350 16882 12402
rect 18062 12350 18114 12402
rect 21646 12350 21698 12402
rect 22990 12350 23042 12402
rect 23438 12350 23490 12402
rect 25790 12350 25842 12402
rect 29262 12350 29314 12402
rect 29934 12350 29986 12402
rect 39678 12350 39730 12402
rect 2494 12238 2546 12290
rect 6078 12238 6130 12290
rect 10558 12238 10610 12290
rect 10894 12238 10946 12290
rect 12910 12238 12962 12290
rect 13358 12238 13410 12290
rect 16494 12238 16546 12290
rect 18958 12238 19010 12290
rect 24110 12238 24162 12290
rect 24446 12238 24498 12290
rect 29598 12238 29650 12290
rect 33854 12238 33906 12290
rect 1822 12126 1874 12178
rect 5406 12126 5458 12178
rect 6190 12126 6242 12178
rect 10222 12126 10274 12178
rect 12350 12126 12402 12178
rect 18398 12126 18450 12178
rect 19182 12126 19234 12178
rect 27022 12126 27074 12178
rect 27918 12126 27970 12178
rect 33070 12126 33122 12178
rect 39118 12126 39170 12178
rect 4622 12014 4674 12066
rect 12686 12014 12738 12066
rect 19742 12014 19794 12066
rect 21534 12014 21586 12066
rect 22878 12014 22930 12066
rect 25342 12014 25394 12066
rect 26350 12014 26402 12066
rect 26910 12014 26962 12066
rect 27470 12014 27522 12066
rect 35982 12014 36034 12066
rect 36318 12014 36370 12066
rect 38446 12014 38498 12066
rect 23774 11902 23826 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 15150 11566 15202 11618
rect 19854 11566 19906 11618
rect 27582 11566 27634 11618
rect 30382 11566 30434 11618
rect 33294 11566 33346 11618
rect 33630 11566 33682 11618
rect 35534 11566 35586 11618
rect 4846 11454 4898 11506
rect 8542 11454 8594 11506
rect 8990 11454 9042 11506
rect 10334 11454 10386 11506
rect 12462 11454 12514 11506
rect 12910 11454 12962 11506
rect 16382 11454 16434 11506
rect 18510 11454 18562 11506
rect 23438 11454 23490 11506
rect 24334 11454 24386 11506
rect 24558 11454 24610 11506
rect 37102 11454 37154 11506
rect 5630 11342 5682 11394
rect 9550 11342 9602 11394
rect 14814 11342 14866 11394
rect 15710 11342 15762 11394
rect 20302 11342 20354 11394
rect 23998 11342 24050 11394
rect 25454 11342 25506 11394
rect 25902 11342 25954 11394
rect 26462 11342 26514 11394
rect 26686 11342 26738 11394
rect 29598 11342 29650 11394
rect 6414 11230 6466 11282
rect 14030 11230 14082 11282
rect 14590 11230 14642 11282
rect 20638 11230 20690 11282
rect 27246 11230 27298 11282
rect 27694 11230 27746 11282
rect 29262 11230 29314 11282
rect 30606 11230 30658 11282
rect 30942 11230 30994 11282
rect 33854 11230 33906 11282
rect 34302 11230 34354 11282
rect 35758 11230 35810 11282
rect 36318 11230 36370 11282
rect 19070 11118 19122 11170
rect 19518 11118 19570 11170
rect 26126 11118 26178 11170
rect 29374 11118 29426 11170
rect 30046 11118 30098 11170
rect 35198 11118 35250 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 6302 10782 6354 10834
rect 13134 10782 13186 10834
rect 17838 10782 17890 10834
rect 18958 10782 19010 10834
rect 29598 10782 29650 10834
rect 29934 10782 29986 10834
rect 30270 10782 30322 10834
rect 35982 10782 36034 10834
rect 7982 10670 8034 10722
rect 12462 10670 12514 10722
rect 14030 10670 14082 10722
rect 16270 10670 16322 10722
rect 18174 10670 18226 10722
rect 24334 10670 24386 10722
rect 26462 10670 26514 10722
rect 30830 10670 30882 10722
rect 35646 10670 35698 10722
rect 6638 10558 6690 10610
rect 7086 10558 7138 10610
rect 7422 10558 7474 10610
rect 8206 10558 8258 10610
rect 12574 10558 12626 10610
rect 14366 10558 14418 10610
rect 16606 10558 16658 10610
rect 18398 10558 18450 10610
rect 19070 10558 19122 10610
rect 20078 10558 20130 10610
rect 24670 10558 24722 10610
rect 25678 10558 25730 10610
rect 30718 10558 30770 10610
rect 31502 10558 31554 10610
rect 15486 10446 15538 10498
rect 19294 10446 19346 10498
rect 20750 10446 20802 10498
rect 22878 10446 22930 10498
rect 23326 10446 23378 10498
rect 25342 10446 25394 10498
rect 28590 10446 28642 10498
rect 11454 10334 11506 10386
rect 11790 10334 11842 10386
rect 31838 10334 31890 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 12462 9998 12514 10050
rect 12798 9998 12850 10050
rect 26462 9998 26514 10050
rect 14254 9886 14306 9938
rect 16382 9886 16434 9938
rect 16942 9886 16994 9938
rect 17950 9886 18002 9938
rect 20078 9886 20130 9938
rect 25006 9886 25058 9938
rect 26014 9886 26066 9938
rect 6638 9774 6690 9826
rect 7646 9774 7698 9826
rect 8094 9774 8146 9826
rect 13470 9774 13522 9826
rect 17278 9774 17330 9826
rect 20414 9774 20466 9826
rect 22318 9774 22370 9826
rect 26798 9774 26850 9826
rect 27358 9774 27410 9826
rect 29934 9774 29986 9826
rect 31054 9774 31106 9826
rect 7310 9662 7362 9714
rect 8318 9662 8370 9714
rect 11902 9662 11954 9714
rect 12238 9662 12290 9714
rect 20750 9662 20802 9714
rect 22542 9662 22594 9714
rect 23102 9662 23154 9714
rect 27582 9662 27634 9714
rect 6862 9550 6914 9602
rect 21982 9550 22034 9602
rect 25566 9550 25618 9602
rect 30158 9550 30210 9602
rect 31278 9550 31330 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 14366 9214 14418 9266
rect 18398 9214 18450 9266
rect 20526 9214 20578 9266
rect 28590 9214 28642 9266
rect 33182 9214 33234 9266
rect 6862 9102 6914 9154
rect 13134 9102 13186 9154
rect 15486 9102 15538 9154
rect 18958 9102 19010 9154
rect 19518 9102 19570 9154
rect 25790 9102 25842 9154
rect 27582 9102 27634 9154
rect 31390 9102 31442 9154
rect 6078 8990 6130 9042
rect 9550 8990 9602 9042
rect 12910 8990 12962 9042
rect 15374 8990 15426 9042
rect 24558 8990 24610 9042
rect 26014 8990 26066 9042
rect 26686 8990 26738 9042
rect 27022 8990 27074 9042
rect 27806 8990 27858 9042
rect 32174 8990 32226 9042
rect 8990 8878 9042 8930
rect 10334 8878 10386 8930
rect 12462 8878 12514 8930
rect 13694 8878 13746 8930
rect 20078 8878 20130 8930
rect 21310 8878 21362 8930
rect 21758 8878 21810 8930
rect 23886 8878 23938 8930
rect 25566 8878 25618 8930
rect 27246 8878 27298 8930
rect 28478 8878 28530 8930
rect 29262 8878 29314 8930
rect 14702 8766 14754 8818
rect 18734 8766 18786 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 9214 8318 9266 8370
rect 13582 8318 13634 8370
rect 22430 8318 22482 8370
rect 25230 8318 25282 8370
rect 26462 8318 26514 8370
rect 28590 8318 28642 8370
rect 30718 8318 30770 8370
rect 32846 8318 32898 8370
rect 10670 8206 10722 8258
rect 13918 8206 13970 8258
rect 18286 8206 18338 8258
rect 18510 8206 18562 8258
rect 19182 8206 19234 8258
rect 19630 8206 19682 8258
rect 20078 8206 20130 8258
rect 20414 8206 20466 8258
rect 21870 8206 21922 8258
rect 22318 8206 22370 8258
rect 22990 8206 23042 8258
rect 23662 8206 23714 8258
rect 23998 8206 24050 8258
rect 24670 8206 24722 8258
rect 25678 8206 25730 8258
rect 33630 8206 33682 8258
rect 34190 8206 34242 8258
rect 10334 8094 10386 8146
rect 14142 8094 14194 8146
rect 14702 8094 14754 8146
rect 17726 8094 17778 8146
rect 18846 8094 18898 8146
rect 22878 8094 22930 8146
rect 24446 8094 24498 8146
rect 12686 7982 12738 8034
rect 20750 7982 20802 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 19182 7646 19234 7698
rect 24110 7646 24162 7698
rect 24670 7646 24722 7698
rect 25342 7646 25394 7698
rect 26798 7646 26850 7698
rect 13358 7534 13410 7586
rect 16494 7534 16546 7586
rect 18510 7534 18562 7586
rect 20974 7534 21026 7586
rect 27358 7534 27410 7586
rect 27918 7534 27970 7586
rect 12574 7422 12626 7474
rect 13246 7422 13298 7474
rect 16830 7422 16882 7474
rect 17502 7422 17554 7474
rect 17838 7422 17890 7474
rect 18286 7422 18338 7474
rect 20302 7422 20354 7474
rect 23998 7422 24050 7474
rect 24222 7422 24274 7474
rect 27134 7422 27186 7474
rect 23102 7310 23154 7362
rect 12238 7198 12290 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 14366 6862 14418 6914
rect 23550 6862 23602 6914
rect 12910 6750 12962 6802
rect 16382 6750 16434 6802
rect 18510 6750 18562 6802
rect 22766 6750 22818 6802
rect 24894 6750 24946 6802
rect 10110 6638 10162 6690
rect 13582 6638 13634 6690
rect 14814 6638 14866 6690
rect 15710 6638 15762 6690
rect 18958 6638 19010 6690
rect 23214 6638 23266 6690
rect 23998 6638 24050 6690
rect 28590 6638 28642 6690
rect 10782 6526 10834 6578
rect 15038 6526 15090 6578
rect 24334 6526 24386 6578
rect 26910 6526 26962 6578
rect 28478 6526 28530 6578
rect 14030 6414 14082 6466
rect 22206 6414 22258 6466
rect 27246 6414 27298 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 11230 6078 11282 6130
rect 14926 6078 14978 6130
rect 26350 6078 26402 6130
rect 26798 6078 26850 6130
rect 13470 5966 13522 6018
rect 13806 5966 13858 6018
rect 16046 5966 16098 6018
rect 16830 5966 16882 6018
rect 18286 5966 18338 6018
rect 18510 5966 18562 6018
rect 22542 5966 22594 6018
rect 24334 5966 24386 6018
rect 27918 5966 27970 6018
rect 11454 5854 11506 5906
rect 15262 5854 15314 5906
rect 15934 5854 15986 5906
rect 16494 5854 16546 5906
rect 17614 5854 17666 5906
rect 17950 5854 18002 5906
rect 21870 5854 21922 5906
rect 22654 5854 22706 5906
rect 23550 5854 23602 5906
rect 24222 5854 24274 5906
rect 27134 5854 27186 5906
rect 27582 5854 27634 5906
rect 25342 5742 25394 5794
rect 25790 5742 25842 5794
rect 26238 5742 26290 5794
rect 21534 5630 21586 5682
rect 23214 5630 23266 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 16270 5182 16322 5234
rect 17278 5182 17330 5234
rect 19406 5182 19458 5234
rect 19854 5182 19906 5234
rect 25006 5182 25058 5234
rect 28254 5182 28306 5234
rect 16606 5070 16658 5122
rect 20526 5070 20578 5122
rect 21534 5070 21586 5122
rect 22094 5070 22146 5122
rect 22878 5070 22930 5122
rect 25342 5070 25394 5122
rect 21758 4958 21810 5010
rect 26126 4958 26178 5010
rect 20750 4846 20802 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 12238 4510 12290 4562
rect 24222 4510 24274 4562
rect 25678 4510 25730 4562
rect 26014 4510 26066 4562
rect 13358 4398 13410 4450
rect 27470 4398 27522 4450
rect 12574 4286 12626 4338
rect 20862 4286 20914 4338
rect 26238 4286 26290 4338
rect 26686 4286 26738 4338
rect 15486 4174 15538 4226
rect 21646 4174 21698 4226
rect 23774 4174 23826 4226
rect 29598 4174 29650 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 26238 3726 26290 3778
rect 26574 3726 26626 3778
rect 27246 3502 27298 3554
rect 27134 3390 27186 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 4032 59200 4144 60000
rect 4480 59200 4592 60000
rect 4928 59200 5040 60000
rect 5376 59200 5488 60000
rect 5824 59200 5936 60000
rect 6272 59200 6384 60000
rect 6720 59200 6832 60000
rect 7168 59200 7280 60000
rect 7616 59200 7728 60000
rect 8064 59200 8176 60000
rect 8512 59200 8624 60000
rect 8960 59200 9072 60000
rect 9408 59200 9520 60000
rect 9856 59200 9968 60000
rect 10304 59200 10416 60000
rect 10752 59200 10864 60000
rect 11200 59200 11312 60000
rect 11648 59200 11760 60000
rect 12096 59200 12208 60000
rect 12544 59200 12656 60000
rect 12992 59200 13104 60000
rect 13440 59200 13552 60000
rect 13888 59200 14000 60000
rect 14336 59200 14448 60000
rect 14784 59200 14896 60000
rect 15232 59200 15344 60000
rect 15680 59200 15792 60000
rect 16128 59200 16240 60000
rect 16576 59200 16688 60000
rect 17024 59200 17136 60000
rect 17472 59200 17584 60000
rect 17920 59200 18032 60000
rect 18368 59200 18480 60000
rect 18816 59200 18928 60000
rect 19264 59200 19376 60000
rect 19712 59200 19824 60000
rect 20160 59200 20272 60000
rect 20608 59200 20720 60000
rect 21056 59200 21168 60000
rect 21504 59200 21616 60000
rect 21952 59200 22064 60000
rect 22400 59200 22512 60000
rect 22848 59200 22960 60000
rect 23296 59200 23408 60000
rect 23744 59200 23856 60000
rect 24192 59200 24304 60000
rect 24640 59200 24752 60000
rect 25088 59200 25200 60000
rect 25536 59200 25648 60000
rect 25984 59200 26096 60000
rect 26432 59200 26544 60000
rect 26880 59200 26992 60000
rect 27328 59200 27440 60000
rect 27776 59200 27888 60000
rect 28224 59200 28336 60000
rect 28672 59200 28784 60000
rect 29120 59200 29232 60000
rect 29568 59200 29680 60000
rect 30016 59200 30128 60000
rect 30464 59200 30576 60000
rect 30912 59200 31024 60000
rect 31360 59200 31472 60000
rect 31808 59200 31920 60000
rect 32256 59200 32368 60000
rect 32704 59200 32816 60000
rect 33152 59200 33264 60000
rect 33600 59200 33712 60000
rect 34048 59200 34160 60000
rect 34496 59200 34608 60000
rect 34944 59200 35056 60000
rect 35392 59200 35504 60000
rect 35840 59200 35952 60000
rect 36288 59200 36400 60000
rect 36736 59200 36848 60000
rect 37184 59200 37296 60000
rect 37632 59200 37744 60000
rect 38080 59200 38192 60000
rect 38528 59200 38640 60000
rect 38976 59200 39088 60000
rect 39424 59200 39536 60000
rect 39872 59200 39984 60000
rect 40320 59200 40432 60000
rect 40768 59200 40880 60000
rect 41216 59200 41328 60000
rect 41664 59200 41776 60000
rect 42112 59200 42224 60000
rect 42560 59200 42672 60000
rect 43008 59200 43120 60000
rect 43456 59200 43568 60000
rect 43904 59200 44016 60000
rect 44352 59200 44464 60000
rect 44800 59200 44912 60000
rect 45248 59200 45360 60000
rect 45696 59200 45808 60000
rect 46144 59200 46256 60000
rect 46592 59200 46704 60000
rect 47040 59200 47152 60000
rect 47488 59200 47600 60000
rect 47936 59200 48048 60000
rect 48384 59200 48496 60000
rect 48832 59200 48944 60000
rect 49280 59200 49392 60000
rect 49728 59200 49840 60000
rect 50176 59200 50288 60000
rect 50624 59200 50736 60000
rect 51072 59200 51184 60000
rect 51520 59200 51632 60000
rect 51968 59200 52080 60000
rect 52416 59200 52528 60000
rect 52864 59200 52976 60000
rect 53312 59200 53424 60000
rect 53760 59200 53872 60000
rect 54208 59200 54320 60000
rect 54656 59200 54768 60000
rect 55104 59200 55216 60000
rect 55552 59200 55664 60000
rect 1820 55298 1876 55310
rect 1820 55246 1822 55298
rect 1874 55246 1876 55298
rect 1820 53730 1876 55246
rect 2492 55186 2548 55198
rect 2492 55134 2494 55186
rect 2546 55134 2548 55186
rect 2492 54738 2548 55134
rect 2492 54686 2494 54738
rect 2546 54686 2548 54738
rect 2492 54674 2548 54686
rect 1820 53678 1822 53730
rect 1874 53678 1876 53730
rect 1820 50594 1876 53678
rect 2380 54626 2436 54638
rect 2380 54574 2382 54626
rect 2434 54574 2436 54626
rect 2380 52724 2436 54574
rect 2604 54516 2660 54526
rect 2940 54516 2996 54526
rect 2604 54514 2996 54516
rect 2604 54462 2606 54514
rect 2658 54462 2942 54514
rect 2994 54462 2996 54514
rect 2604 54460 2996 54462
rect 2604 54450 2660 54460
rect 2940 54450 2996 54460
rect 3388 54514 3444 54526
rect 3388 54462 3390 54514
rect 3442 54462 3444 54514
rect 3276 54402 3332 54414
rect 3276 54350 3278 54402
rect 3330 54350 3332 54402
rect 2492 53620 2548 53630
rect 2492 53618 2772 53620
rect 2492 53566 2494 53618
rect 2546 53566 2772 53618
rect 2492 53564 2772 53566
rect 2492 53554 2548 53564
rect 2716 53170 2772 53564
rect 2716 53118 2718 53170
rect 2770 53118 2772 53170
rect 2716 53106 2772 53118
rect 2940 52948 2996 52958
rect 3276 52948 3332 54350
rect 2940 52946 3332 52948
rect 2940 52894 2942 52946
rect 2994 52894 3278 52946
rect 3330 52894 3332 52946
rect 2940 52892 3332 52894
rect 3388 52948 3444 54462
rect 4060 53844 4116 59200
rect 4508 56308 4564 59200
rect 5404 56420 5460 59200
rect 5852 57540 5908 59200
rect 5852 57484 6244 57540
rect 4956 56364 5460 56420
rect 4620 56308 4676 56318
rect 4508 56252 4620 56308
rect 4620 56214 4676 56252
rect 4956 56306 5012 56364
rect 4956 56254 4958 56306
rect 5010 56254 5012 56306
rect 4956 56242 5012 56254
rect 5516 56308 5572 56318
rect 5516 56194 5572 56252
rect 5516 56142 5518 56194
rect 5570 56142 5572 56194
rect 5516 56130 5572 56142
rect 5852 56196 5908 56206
rect 5852 56102 5908 56140
rect 6188 55970 6244 57484
rect 6748 56308 6804 59200
rect 6972 56308 7028 56318
rect 6748 56306 7028 56308
rect 6748 56254 6974 56306
rect 7026 56254 7028 56306
rect 6748 56252 7028 56254
rect 6972 56242 7028 56252
rect 6188 55918 6190 55970
rect 6242 55918 6244 55970
rect 6188 55906 6244 55918
rect 7196 55972 7252 59200
rect 8092 56308 8148 59200
rect 8204 56308 8260 56318
rect 8092 56306 8260 56308
rect 8092 56254 8206 56306
rect 8258 56254 8260 56306
rect 8092 56252 8260 56254
rect 8204 56242 8260 56252
rect 8428 56196 8484 56206
rect 7420 55972 7476 55982
rect 7196 55970 7476 55972
rect 7196 55918 7422 55970
rect 7474 55918 7476 55970
rect 7196 55916 7476 55918
rect 7420 55906 7476 55916
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 8428 55468 8484 56140
rect 8540 55972 8596 59200
rect 9436 56308 9492 59200
rect 9660 56308 9716 56318
rect 9436 56306 9716 56308
rect 9436 56254 9662 56306
rect 9714 56254 9716 56306
rect 9436 56252 9716 56254
rect 9660 56242 9716 56252
rect 8652 55972 8708 55982
rect 8540 55970 8708 55972
rect 8540 55918 8654 55970
rect 8706 55918 8708 55970
rect 8540 55916 8708 55918
rect 9884 55972 9940 59200
rect 10780 56308 10836 59200
rect 11004 56308 11060 56318
rect 10780 56306 11060 56308
rect 10780 56254 11006 56306
rect 11058 56254 11060 56306
rect 10780 56252 11060 56254
rect 11004 56242 11060 56252
rect 10108 55972 10164 55982
rect 9884 55970 10164 55972
rect 9884 55918 10110 55970
rect 10162 55918 10164 55970
rect 9884 55916 10164 55918
rect 11228 55972 11284 59200
rect 12124 56308 12180 59200
rect 12572 56642 12628 59200
rect 12572 56590 12574 56642
rect 12626 56590 12628 56642
rect 12572 56578 12628 56590
rect 13132 56642 13188 56654
rect 13132 56590 13134 56642
rect 13186 56590 13188 56642
rect 12348 56308 12404 56318
rect 12124 56306 12404 56308
rect 12124 56254 12350 56306
rect 12402 56254 12404 56306
rect 12124 56252 12404 56254
rect 12348 56242 12404 56252
rect 11452 55972 11508 55982
rect 11228 55970 11508 55972
rect 11228 55918 11454 55970
rect 11506 55918 11508 55970
rect 11228 55916 11508 55918
rect 8652 55906 8708 55916
rect 10108 55906 10164 55916
rect 11452 55906 11508 55916
rect 13132 55970 13188 56590
rect 13468 56308 13524 59200
rect 13692 56308 13748 56318
rect 13468 56306 13748 56308
rect 13468 56254 13694 56306
rect 13746 56254 13748 56306
rect 13468 56252 13748 56254
rect 13692 56242 13748 56252
rect 13132 55918 13134 55970
rect 13186 55918 13188 55970
rect 13132 55906 13188 55918
rect 13916 55972 13972 59200
rect 14700 56308 14756 56318
rect 14812 56308 14868 59200
rect 14700 56306 14868 56308
rect 14700 56254 14702 56306
rect 14754 56254 14868 56306
rect 14700 56252 14868 56254
rect 15148 57090 15204 57102
rect 15148 57038 15150 57090
rect 15202 57038 15204 57090
rect 15148 56306 15204 57038
rect 15148 56254 15150 56306
rect 15202 56254 15204 56306
rect 14700 56242 14756 56252
rect 15148 56242 15204 56254
rect 14812 56084 14868 56094
rect 14140 55972 14196 55982
rect 13916 55970 14196 55972
rect 13916 55918 14142 55970
rect 14194 55918 14196 55970
rect 13916 55916 14196 55918
rect 14140 55906 14196 55916
rect 4620 55410 4676 55422
rect 4620 55358 4622 55410
rect 4674 55358 4676 55410
rect 4620 54740 4676 55358
rect 5852 55410 5908 55422
rect 8428 55412 8708 55468
rect 5852 55358 5854 55410
rect 5906 55358 5908 55410
rect 4172 54684 4676 54740
rect 5068 55074 5124 55086
rect 5068 55022 5070 55074
rect 5122 55022 5124 55074
rect 4172 53844 4228 54684
rect 4396 54516 4452 54526
rect 4284 54514 4452 54516
rect 4284 54462 4398 54514
rect 4450 54462 4452 54514
rect 4284 54460 4452 54462
rect 4284 53956 4340 54460
rect 4396 54450 4452 54460
rect 4956 54402 5012 54414
rect 4956 54350 4958 54402
rect 5010 54350 5012 54402
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4284 53900 4676 53956
rect 4172 53788 4340 53844
rect 4060 53778 4116 53788
rect 3500 53172 3556 53182
rect 3500 53170 4228 53172
rect 3500 53118 3502 53170
rect 3554 53118 4228 53170
rect 3500 53116 4228 53118
rect 3500 53106 3556 53116
rect 3612 52948 3668 52958
rect 3388 52946 3668 52948
rect 3388 52894 3614 52946
rect 3666 52894 3668 52946
rect 3388 52892 3668 52894
rect 2940 52882 2996 52892
rect 3276 52836 3332 52892
rect 3276 52770 3332 52780
rect 2604 52724 2660 52734
rect 2380 52722 3108 52724
rect 2380 52670 2606 52722
rect 2658 52670 3108 52722
rect 2380 52668 3108 52670
rect 2604 52658 2660 52668
rect 2492 51940 2548 51950
rect 2492 50706 2548 51884
rect 2492 50654 2494 50706
rect 2546 50654 2548 50706
rect 2492 50642 2548 50654
rect 1820 50542 1822 50594
rect 1874 50542 1876 50594
rect 1820 49810 1876 50542
rect 1820 49758 1822 49810
rect 1874 49758 1876 49810
rect 1820 47458 1876 49758
rect 2492 49698 2548 49710
rect 2492 49646 2494 49698
rect 2546 49646 2548 49698
rect 2492 48804 2548 49646
rect 2492 48738 2548 48748
rect 3052 48356 3108 52668
rect 3612 52052 3668 52892
rect 3612 51986 3668 51996
rect 3836 52948 3892 52958
rect 3836 50820 3892 52892
rect 4172 52162 4228 53116
rect 4172 52110 4174 52162
rect 4226 52110 4228 52162
rect 4172 52098 4228 52110
rect 4284 52946 4340 53788
rect 4396 53058 4452 53900
rect 4620 53842 4676 53900
rect 4620 53790 4622 53842
rect 4674 53790 4676 53842
rect 4620 53778 4676 53790
rect 4396 53006 4398 53058
rect 4450 53006 4452 53058
rect 4396 52994 4452 53006
rect 4284 52894 4286 52946
rect 4338 52894 4340 52946
rect 4284 52164 4340 52894
rect 4508 52948 4564 52958
rect 4508 52854 4564 52892
rect 4956 52948 5012 54350
rect 4956 52882 5012 52892
rect 5068 53506 5124 55022
rect 5852 54516 5908 55358
rect 7980 55188 8036 55198
rect 7644 55186 8036 55188
rect 7644 55134 7982 55186
rect 8034 55134 8036 55186
rect 7644 55132 8036 55134
rect 7532 54626 7588 54638
rect 7532 54574 7534 54626
rect 7586 54574 7588 54626
rect 6524 54516 6580 54526
rect 6972 54516 7028 54526
rect 7308 54516 7364 54526
rect 5852 54514 6692 54516
rect 5852 54462 6526 54514
rect 6578 54462 6692 54514
rect 5852 54460 6692 54462
rect 6524 54450 6580 54460
rect 5068 53454 5070 53506
rect 5122 53454 5124 53506
rect 4956 52722 5012 52734
rect 4956 52670 4958 52722
rect 5010 52670 5012 52722
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4396 52388 4452 52398
rect 4396 52294 4452 52332
rect 4956 52276 5012 52670
rect 4956 52210 5012 52220
rect 4620 52164 4676 52174
rect 4284 52108 4452 52164
rect 4396 52052 4452 52108
rect 4620 52162 4788 52164
rect 4620 52110 4622 52162
rect 4674 52110 4788 52162
rect 4620 52108 4788 52110
rect 4620 52098 4676 52108
rect 4284 51940 4340 51950
rect 4396 51940 4452 51996
rect 4396 51884 4676 51940
rect 4284 51846 4340 51884
rect 4620 51490 4676 51884
rect 4620 51438 4622 51490
rect 4674 51438 4676 51490
rect 4620 51426 4676 51438
rect 4732 51156 4788 52108
rect 4732 51100 5012 51156
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 3836 50754 3892 50764
rect 4620 50820 4676 50830
rect 4620 50706 4676 50764
rect 4620 50654 4622 50706
rect 4674 50654 4676 50706
rect 4620 50642 4676 50654
rect 4956 50708 5012 51100
rect 4060 50596 4116 50606
rect 4060 50428 4116 50540
rect 4060 50372 4228 50428
rect 4172 49250 4228 50372
rect 4620 49700 4676 49710
rect 4620 49698 4900 49700
rect 4620 49646 4622 49698
rect 4674 49646 4900 49698
rect 4620 49644 4900 49646
rect 4620 49634 4676 49644
rect 4844 49476 4900 49644
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4844 49410 4900 49420
rect 4476 49354 4740 49364
rect 4956 49252 5012 50652
rect 4172 49198 4174 49250
rect 4226 49198 4228 49250
rect 4172 49186 4228 49198
rect 4844 49250 5012 49252
rect 4844 49198 4958 49250
rect 5010 49198 5012 49250
rect 4844 49196 5012 49198
rect 3948 49140 4004 49150
rect 3948 48914 4004 49084
rect 4060 49028 4116 49038
rect 4508 49028 4564 49038
rect 4060 49026 4564 49028
rect 4060 48974 4062 49026
rect 4114 48974 4510 49026
rect 4562 48974 4564 49026
rect 4060 48972 4564 48974
rect 4060 48962 4116 48972
rect 4508 48962 4564 48972
rect 4732 49028 4788 49038
rect 4732 48934 4788 48972
rect 3948 48862 3950 48914
rect 4002 48862 4004 48914
rect 3948 48850 4004 48862
rect 4620 48804 4676 48814
rect 4620 48710 4676 48748
rect 4844 48580 4900 49196
rect 4956 49186 5012 49196
rect 5068 50370 5124 53454
rect 6188 52836 6244 52846
rect 5852 51938 5908 51950
rect 5852 51886 5854 51938
rect 5906 51886 5908 51938
rect 5852 50596 5908 51886
rect 6188 51378 6244 52780
rect 6412 52388 6468 52398
rect 6300 52276 6356 52286
rect 6300 52162 6356 52220
rect 6300 52110 6302 52162
rect 6354 52110 6356 52162
rect 6300 52098 6356 52110
rect 6412 52162 6468 52332
rect 6412 52110 6414 52162
rect 6466 52110 6468 52162
rect 6412 52098 6468 52110
rect 6636 52164 6692 54460
rect 6972 54514 7364 54516
rect 6972 54462 6974 54514
rect 7026 54462 7310 54514
rect 7362 54462 7364 54514
rect 6972 54460 7364 54462
rect 6972 54450 7028 54460
rect 7308 54450 7364 54460
rect 6748 54402 6804 54414
rect 6748 54350 6750 54402
rect 6802 54350 6804 54402
rect 6748 52276 6804 54350
rect 7532 52612 7588 54574
rect 7644 54402 7700 55132
rect 7980 55122 8036 55132
rect 7644 54350 7646 54402
rect 7698 54350 7700 54402
rect 7644 54338 7700 54350
rect 6748 52164 6804 52220
rect 6972 52556 7588 52612
rect 8092 53060 8148 53070
rect 6860 52164 6916 52174
rect 6748 52162 6916 52164
rect 6748 52110 6862 52162
rect 6914 52110 6916 52162
rect 6748 52108 6916 52110
rect 6636 52070 6692 52108
rect 6860 52098 6916 52108
rect 6188 51326 6190 51378
rect 6242 51326 6244 51378
rect 6188 51314 6244 51326
rect 6748 51378 6804 51390
rect 6748 51326 6750 51378
rect 6802 51326 6804 51378
rect 6076 51266 6132 51278
rect 6076 51214 6078 51266
rect 6130 51214 6132 51266
rect 5964 50596 6020 50606
rect 5852 50540 5964 50596
rect 5964 50502 6020 50540
rect 5068 50318 5070 50370
rect 5122 50318 5124 50370
rect 5068 49700 5124 50318
rect 5628 50370 5684 50382
rect 5628 50318 5630 50370
rect 5682 50318 5684 50370
rect 5404 49810 5460 49822
rect 5404 49758 5406 49810
rect 5458 49758 5460 49810
rect 5404 49700 5460 49758
rect 5068 49698 5460 49700
rect 5068 49646 5070 49698
rect 5122 49646 5460 49698
rect 5068 49644 5460 49646
rect 4284 48524 4900 48580
rect 4956 48916 5012 48926
rect 4284 48466 4340 48524
rect 4284 48414 4286 48466
rect 4338 48414 4340 48466
rect 4284 48402 4340 48414
rect 4956 48356 5012 48860
rect 2828 48244 2884 48254
rect 2492 48242 2884 48244
rect 2492 48190 2830 48242
rect 2882 48190 2884 48242
rect 2492 48188 2884 48190
rect 2492 47570 2548 48188
rect 2828 48178 2884 48188
rect 3052 48242 3108 48300
rect 4620 48300 5012 48356
rect 3052 48190 3054 48242
rect 3106 48190 3108 48242
rect 3052 48178 3108 48190
rect 4060 48244 4116 48254
rect 4060 48150 4116 48188
rect 4620 48130 4676 48300
rect 4956 48132 5012 48142
rect 4620 48078 4622 48130
rect 4674 48078 4676 48130
rect 4620 48066 4676 48078
rect 4844 48076 4956 48132
rect 2716 48020 2772 48030
rect 2492 47518 2494 47570
rect 2546 47518 2548 47570
rect 2492 47506 2548 47518
rect 2604 48018 2772 48020
rect 2604 47966 2718 48018
rect 2770 47966 2772 48018
rect 2604 47964 2772 47966
rect 1820 47406 1822 47458
rect 1874 47406 1876 47458
rect 1820 46004 1876 47406
rect 2492 46788 2548 46798
rect 2604 46788 2660 47964
rect 2716 47954 2772 47964
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4620 47572 4676 47582
rect 4284 47570 4676 47572
rect 4284 47518 4622 47570
rect 4674 47518 4676 47570
rect 4284 47516 4676 47518
rect 2492 46786 2660 46788
rect 2492 46734 2494 46786
rect 2546 46734 2660 46786
rect 2492 46732 2660 46734
rect 3948 46786 4004 46798
rect 3948 46734 3950 46786
rect 4002 46734 4004 46786
rect 2492 46722 2548 46732
rect 3164 46674 3220 46686
rect 3164 46622 3166 46674
rect 3218 46622 3220 46674
rect 3164 46452 3220 46622
rect 3388 46676 3444 46686
rect 3724 46676 3780 46686
rect 3388 46674 3780 46676
rect 3388 46622 3390 46674
rect 3442 46622 3726 46674
rect 3778 46622 3780 46674
rect 3388 46620 3780 46622
rect 3388 46610 3444 46620
rect 3724 46610 3780 46620
rect 3388 46452 3444 46462
rect 3164 46396 3388 46452
rect 3388 46386 3444 46396
rect 1820 45890 1876 45948
rect 1820 45838 1822 45890
rect 1874 45838 1876 45890
rect 1820 43538 1876 45838
rect 2492 45780 2548 45790
rect 2380 45778 2548 45780
rect 2380 45726 2494 45778
rect 2546 45726 2548 45778
rect 2380 45724 2548 45726
rect 2268 45220 2324 45230
rect 2268 44322 2324 45164
rect 2380 44436 2436 45724
rect 2492 45714 2548 45724
rect 2604 45332 2660 45342
rect 2604 45330 2884 45332
rect 2604 45278 2606 45330
rect 2658 45278 2884 45330
rect 2604 45276 2884 45278
rect 2604 45266 2660 45276
rect 2492 45220 2548 45230
rect 2492 45126 2548 45164
rect 2716 45108 2772 45118
rect 2492 44436 2548 44446
rect 2380 44434 2548 44436
rect 2380 44382 2494 44434
rect 2546 44382 2548 44434
rect 2380 44380 2548 44382
rect 2492 44370 2548 44380
rect 2268 44270 2270 44322
rect 2322 44270 2324 44322
rect 2268 44258 2324 44270
rect 2716 44322 2772 45052
rect 2716 44270 2718 44322
rect 2770 44270 2772 44322
rect 2716 44258 2772 44270
rect 2828 44322 2884 45276
rect 3500 45220 3556 45230
rect 3164 45108 3220 45118
rect 3164 45106 3332 45108
rect 3164 45054 3166 45106
rect 3218 45054 3332 45106
rect 3164 45052 3332 45054
rect 3164 45042 3220 45052
rect 3276 44548 3332 45052
rect 3388 44548 3444 44558
rect 3276 44492 3388 44548
rect 3388 44482 3444 44492
rect 2828 44270 2830 44322
rect 2882 44270 2884 44322
rect 2828 44258 2884 44270
rect 3388 44322 3444 44334
rect 3388 44270 3390 44322
rect 3442 44270 3444 44322
rect 3276 44210 3332 44222
rect 3276 44158 3278 44210
rect 3330 44158 3332 44210
rect 3276 43708 3332 44158
rect 2492 43652 3332 43708
rect 2492 43650 2548 43652
rect 2492 43598 2494 43650
rect 2546 43598 2548 43650
rect 2492 43586 2548 43598
rect 1820 43486 1822 43538
rect 1874 43486 1876 43538
rect 1820 43474 1876 43486
rect 3388 43540 3444 44270
rect 3388 43474 3444 43484
rect 3500 44324 3556 45164
rect 3948 45108 4004 46734
rect 4060 46674 4116 46686
rect 4060 46622 4062 46674
rect 4114 46622 4116 46674
rect 4060 45220 4116 46622
rect 4284 46452 4340 47516
rect 4620 47506 4676 47516
rect 4284 46116 4340 46396
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4284 46060 4564 46116
rect 4060 45154 4116 45164
rect 4508 45218 4564 46060
rect 4508 45166 4510 45218
rect 4562 45166 4564 45218
rect 4508 45154 4564 45166
rect 4620 46002 4676 46014
rect 4620 45950 4622 46002
rect 4674 45950 4676 46002
rect 3948 45042 4004 45052
rect 4620 45108 4676 45950
rect 4620 45042 4676 45052
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 3612 44548 3668 44558
rect 4172 44548 4228 44558
rect 3612 44546 4228 44548
rect 3612 44494 3614 44546
rect 3666 44494 4174 44546
rect 4226 44494 4228 44546
rect 3612 44492 4228 44494
rect 3612 44482 3668 44492
rect 4172 44482 4228 44492
rect 3724 44324 3780 44334
rect 4508 44324 4564 44334
rect 3500 44322 3780 44324
rect 3500 44270 3726 44322
rect 3778 44270 3780 44322
rect 3500 44268 3780 44270
rect 3388 42980 3444 42990
rect 3500 42980 3556 44268
rect 3724 44258 3780 44268
rect 3836 44322 4564 44324
rect 3836 44270 4510 44322
rect 4562 44270 4564 44322
rect 3836 44268 4564 44270
rect 3388 42978 3556 42980
rect 3388 42926 3390 42978
rect 3442 42926 3556 42978
rect 3388 42924 3556 42926
rect 3612 44100 3668 44110
rect 3388 42914 3444 42924
rect 2828 41972 2884 41982
rect 2828 41878 2884 41916
rect 3388 41972 3444 41982
rect 3612 41972 3668 44044
rect 3388 41970 3668 41972
rect 3388 41918 3390 41970
rect 3442 41918 3668 41970
rect 3388 41916 3668 41918
rect 3724 42980 3780 42990
rect 3836 42980 3892 44268
rect 4508 44258 4564 44268
rect 4844 44324 4900 48076
rect 4956 48066 5012 48076
rect 5068 47234 5124 49644
rect 5628 49028 5684 50318
rect 5964 50372 6020 50382
rect 5628 48962 5684 48972
rect 5740 50148 5796 50158
rect 5740 49140 5796 50092
rect 5740 47460 5796 49084
rect 5852 49026 5908 49038
rect 5852 48974 5854 49026
rect 5906 48974 5908 49026
rect 5852 48916 5908 48974
rect 5852 48850 5908 48860
rect 5964 48804 6020 50316
rect 6076 49252 6132 51214
rect 6748 50820 6804 51326
rect 6748 50754 6804 50764
rect 6636 50708 6692 50718
rect 6188 50594 6244 50606
rect 6188 50542 6190 50594
rect 6242 50542 6244 50594
rect 6188 50148 6244 50542
rect 6524 50484 6580 50494
rect 6188 50082 6244 50092
rect 6300 50482 6580 50484
rect 6300 50430 6526 50482
rect 6578 50430 6580 50482
rect 6300 50428 6580 50430
rect 6188 49924 6244 49934
rect 6300 49924 6356 50428
rect 6524 50418 6580 50428
rect 6636 50428 6692 50652
rect 6860 50596 6916 50606
rect 6860 50502 6916 50540
rect 6636 50372 6916 50428
rect 6188 49922 6356 49924
rect 6188 49870 6190 49922
rect 6242 49870 6356 49922
rect 6188 49868 6356 49870
rect 6188 49858 6244 49868
rect 6076 49196 6244 49252
rect 6076 49028 6132 49038
rect 6076 48934 6132 48972
rect 5964 48748 6132 48804
rect 5964 47460 6020 47470
rect 5740 47458 6020 47460
rect 5740 47406 5966 47458
rect 6018 47406 6020 47458
rect 5740 47404 6020 47406
rect 5964 47394 6020 47404
rect 6076 47346 6132 48748
rect 6076 47294 6078 47346
rect 6130 47294 6132 47346
rect 6076 47282 6132 47294
rect 5068 47182 5070 47234
rect 5122 47182 5124 47234
rect 5068 46004 5124 47182
rect 5068 45666 5124 45948
rect 5068 45614 5070 45666
rect 5122 45614 5124 45666
rect 5068 45556 5124 45614
rect 5628 45890 5684 45902
rect 5628 45838 5630 45890
rect 5682 45838 5684 45890
rect 5068 45500 5572 45556
rect 4956 45108 5012 45118
rect 5404 45108 5460 45118
rect 4956 45014 5012 45052
rect 5180 45106 5460 45108
rect 5180 45054 5406 45106
rect 5458 45054 5460 45106
rect 5180 45052 5460 45054
rect 4956 44324 5012 44334
rect 4844 44322 5012 44324
rect 4844 44270 4958 44322
rect 5010 44270 5012 44322
rect 4844 44268 5012 44270
rect 3724 42978 3892 42980
rect 3724 42926 3726 42978
rect 3778 42926 3892 42978
rect 3724 42924 3892 42926
rect 3724 41972 3780 42924
rect 3836 42644 3892 42924
rect 4284 44098 4340 44110
rect 4284 44046 4286 44098
rect 4338 44046 4340 44098
rect 4284 43316 4340 44046
rect 4844 43988 4900 44268
rect 4956 44258 5012 44268
rect 5068 44100 5124 44110
rect 5068 44006 5124 44044
rect 4732 43932 4900 43988
rect 4620 43764 4676 43774
rect 4620 43426 4676 43708
rect 4620 43374 4622 43426
rect 4674 43374 4676 43426
rect 4620 43316 4676 43374
rect 4732 43428 4788 43932
rect 4956 43764 5012 43774
rect 4732 43362 4788 43372
rect 4844 43652 4900 43662
rect 4284 43260 4676 43316
rect 3948 42868 4004 42878
rect 4284 42868 4340 43260
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 3948 42866 4340 42868
rect 3948 42814 3950 42866
rect 4002 42814 4340 42866
rect 3948 42812 4340 42814
rect 4732 42868 4788 42878
rect 4844 42868 4900 43596
rect 4956 43650 5012 43708
rect 5068 43764 5124 43774
rect 5180 43764 5236 45052
rect 5404 45042 5460 45052
rect 5516 44324 5572 45500
rect 5628 45330 5684 45838
rect 6188 45890 6244 49196
rect 6860 49250 6916 50372
rect 6860 49198 6862 49250
rect 6914 49198 6916 49250
rect 6860 49186 6916 49198
rect 6748 48914 6804 48926
rect 6748 48862 6750 48914
rect 6802 48862 6804 48914
rect 6412 48804 6468 48814
rect 6524 48804 6580 48814
rect 6412 48802 6524 48804
rect 6412 48750 6414 48802
rect 6466 48750 6524 48802
rect 6412 48748 6524 48750
rect 6412 48738 6468 48748
rect 6524 47068 6580 48748
rect 6748 48354 6804 48862
rect 6748 48302 6750 48354
rect 6802 48302 6804 48354
rect 6748 48290 6804 48302
rect 6972 48356 7028 52556
rect 7532 52388 7588 52398
rect 7196 52164 7252 52174
rect 7084 51938 7140 51950
rect 7084 51886 7086 51938
rect 7138 51886 7140 51938
rect 7084 50594 7140 51886
rect 7196 51490 7252 52108
rect 7196 51438 7198 51490
rect 7250 51438 7252 51490
rect 7196 51426 7252 51438
rect 7532 52050 7588 52332
rect 7980 52276 8036 52286
rect 8092 52276 8148 53004
rect 7980 52274 8148 52276
rect 7980 52222 7982 52274
rect 8034 52222 8148 52274
rect 7980 52220 8148 52222
rect 7980 52210 8036 52220
rect 7532 51998 7534 52050
rect 7586 51998 7588 52050
rect 7084 50542 7086 50594
rect 7138 50542 7140 50594
rect 7084 50530 7140 50542
rect 7532 50482 7588 51998
rect 8092 50596 8148 52220
rect 8540 53060 8596 53070
rect 8540 52162 8596 53004
rect 8540 52110 8542 52162
rect 8594 52110 8596 52162
rect 8540 52098 8596 52110
rect 8092 50594 8372 50596
rect 8092 50542 8094 50594
rect 8146 50542 8372 50594
rect 8092 50540 8372 50542
rect 8092 50530 8148 50540
rect 7532 50430 7534 50482
rect 7586 50430 7588 50482
rect 7420 50372 7476 50382
rect 7420 50278 7476 50316
rect 7532 49700 7588 50430
rect 8316 50428 8372 50540
rect 8316 50372 8484 50428
rect 8316 49700 8372 49710
rect 7532 49698 8372 49700
rect 7532 49646 8318 49698
rect 8370 49646 8372 49698
rect 7532 49644 8372 49646
rect 8316 49634 8372 49644
rect 7084 49252 7140 49262
rect 7084 49250 7364 49252
rect 7084 49198 7086 49250
rect 7138 49198 7364 49250
rect 7084 49196 7364 49198
rect 7084 49186 7140 49196
rect 7308 49140 7364 49196
rect 7756 49140 7812 49150
rect 7308 49138 7812 49140
rect 7308 49086 7758 49138
rect 7810 49086 7812 49138
rect 7308 49084 7812 49086
rect 7756 49074 7812 49084
rect 7196 49026 7252 49038
rect 7196 48974 7198 49026
rect 7250 48974 7252 49026
rect 6972 48290 7028 48300
rect 7084 48916 7140 48926
rect 7084 48468 7140 48860
rect 7196 48804 7252 48974
rect 7644 48916 7700 48926
rect 7644 48822 7700 48860
rect 7868 48804 7924 48814
rect 7196 48738 7252 48748
rect 7756 48802 7924 48804
rect 7756 48750 7870 48802
rect 7922 48750 7924 48802
rect 7756 48748 7924 48750
rect 7756 48468 7812 48748
rect 7868 48738 7924 48748
rect 8428 48804 8484 50372
rect 8652 49028 8708 55412
rect 14812 55410 14868 56028
rect 14812 55358 14814 55410
rect 14866 55358 14868 55410
rect 14812 55346 14868 55358
rect 15148 55972 15204 55982
rect 8764 55298 8820 55310
rect 8764 55246 8766 55298
rect 8818 55246 8820 55298
rect 8764 55076 8820 55246
rect 15148 55300 15204 55916
rect 15260 55524 15316 59200
rect 15596 57092 15652 57102
rect 15596 56306 15652 57036
rect 15596 56254 15598 56306
rect 15650 56254 15652 56306
rect 15596 56242 15652 56254
rect 15708 56308 15764 59200
rect 16156 57540 16212 59200
rect 16044 57484 16212 57540
rect 16044 57090 16100 57484
rect 16604 57428 16660 59200
rect 16044 57038 16046 57090
rect 16098 57038 16100 57090
rect 16044 57026 16100 57038
rect 16156 57372 16660 57428
rect 15932 56308 15988 56318
rect 15764 56306 15988 56308
rect 15764 56254 15934 56306
rect 15986 56254 15988 56306
rect 15764 56252 15988 56254
rect 15708 56214 15764 56252
rect 15932 56242 15988 56252
rect 15484 55524 15540 55534
rect 15260 55522 15540 55524
rect 15260 55470 15486 55522
rect 15538 55470 15540 55522
rect 15260 55468 15540 55470
rect 15484 55458 15540 55468
rect 16156 55522 16212 57372
rect 16156 55470 16158 55522
rect 16210 55470 16212 55522
rect 16156 55458 16212 55470
rect 16268 56194 16324 56206
rect 16268 56142 16270 56194
rect 16322 56142 16324 56194
rect 15260 55300 15316 55310
rect 15148 55298 15316 55300
rect 15148 55246 15262 55298
rect 15314 55246 15316 55298
rect 15148 55244 15316 55246
rect 15260 55234 15316 55244
rect 9212 55076 9268 55086
rect 8764 55074 9268 55076
rect 8764 55022 9214 55074
rect 9266 55022 9268 55074
rect 8764 55020 9268 55022
rect 9212 54516 9268 55020
rect 9212 54450 9268 54460
rect 9996 54516 10052 54526
rect 9324 53844 9380 53854
rect 9212 52052 9268 52062
rect 9212 51958 9268 51996
rect 8764 51156 8820 51166
rect 8764 50706 8820 51100
rect 8764 50654 8766 50706
rect 8818 50654 8820 50706
rect 8764 50642 8820 50654
rect 9324 50428 9380 53788
rect 9548 53844 9604 53854
rect 9996 53844 10052 54460
rect 12124 54516 12180 54526
rect 12460 54516 12516 54526
rect 12180 54514 12516 54516
rect 12180 54462 12462 54514
rect 12514 54462 12516 54514
rect 12180 54460 12516 54462
rect 12124 54422 12180 54460
rect 12460 54450 12516 54460
rect 16268 54514 16324 56142
rect 17052 56196 17108 59200
rect 17500 57092 17556 59200
rect 17500 57026 17556 57036
rect 17276 56196 17332 56206
rect 17052 56194 17332 56196
rect 17052 56142 17278 56194
rect 17330 56142 17332 56194
rect 17052 56140 17332 56142
rect 17052 55972 17108 56140
rect 17276 56130 17332 56140
rect 17612 56194 17668 56206
rect 17612 56142 17614 56194
rect 17666 56142 17668 56194
rect 17052 55906 17108 55916
rect 16492 55412 16548 55422
rect 16492 55298 16548 55356
rect 16492 55246 16494 55298
rect 16546 55246 16548 55298
rect 16492 55234 16548 55246
rect 16604 55300 16660 55310
rect 17164 55300 17220 55310
rect 16604 55186 16660 55244
rect 16940 55298 17220 55300
rect 16940 55246 17166 55298
rect 17218 55246 17220 55298
rect 16940 55244 17220 55246
rect 16604 55134 16606 55186
rect 16658 55134 16660 55186
rect 16604 55122 16660 55134
rect 16828 55188 16884 55198
rect 16828 55094 16884 55132
rect 16828 54740 16884 54750
rect 16940 54740 16996 55244
rect 17164 55234 17220 55244
rect 17388 55298 17444 55310
rect 17388 55246 17390 55298
rect 17442 55246 17444 55298
rect 16828 54738 16996 54740
rect 16828 54686 16830 54738
rect 16882 54686 16996 54738
rect 16828 54684 16996 54686
rect 17052 55074 17108 55086
rect 17052 55022 17054 55074
rect 17106 55022 17108 55074
rect 16828 54674 16884 54684
rect 16268 54462 16270 54514
rect 16322 54462 16324 54514
rect 13244 54404 13300 54414
rect 15372 54404 15428 54414
rect 13244 54402 13412 54404
rect 13244 54350 13246 54402
rect 13298 54350 13412 54402
rect 13244 54348 13412 54350
rect 13244 54338 13300 54348
rect 12908 53956 12964 53966
rect 9548 53842 10052 53844
rect 9548 53790 9550 53842
rect 9602 53790 10052 53842
rect 9548 53788 10052 53790
rect 9548 53060 9604 53788
rect 9996 53730 10052 53788
rect 9996 53678 9998 53730
rect 10050 53678 10052 53730
rect 9996 53666 10052 53678
rect 10668 53844 10724 53854
rect 10668 53730 10724 53788
rect 10668 53678 10670 53730
rect 10722 53678 10724 53730
rect 10668 53666 10724 53678
rect 12796 53842 12852 53854
rect 12796 53790 12798 53842
rect 12850 53790 12852 53842
rect 9548 52994 9604 53004
rect 11452 52948 11508 52958
rect 11452 52854 11508 52892
rect 12460 52946 12516 52958
rect 12460 52894 12462 52946
rect 12514 52894 12516 52946
rect 10332 52834 10388 52846
rect 10332 52782 10334 52834
rect 10386 52782 10388 52834
rect 10332 51492 10388 52782
rect 10892 52836 10948 52846
rect 10892 52742 10948 52780
rect 12012 52836 12068 52846
rect 12068 52780 12180 52836
rect 12012 52742 12068 52780
rect 10332 51426 10388 51436
rect 10556 52722 10612 52734
rect 10556 52670 10558 52722
rect 10610 52670 10612 52722
rect 10556 51380 10612 52670
rect 11564 52722 11620 52734
rect 11564 52670 11566 52722
rect 11618 52670 11620 52722
rect 11340 52274 11396 52286
rect 11340 52222 11342 52274
rect 11394 52222 11396 52274
rect 11340 51492 11396 52222
rect 11564 52276 11620 52670
rect 11564 52210 11620 52220
rect 11004 51380 11060 51390
rect 10556 51378 11060 51380
rect 10556 51326 10558 51378
rect 10610 51326 11006 51378
rect 11058 51326 11060 51378
rect 10556 51324 11060 51326
rect 10108 51156 10164 51166
rect 10108 51062 10164 51100
rect 10220 51154 10276 51166
rect 10220 51102 10222 51154
rect 10274 51102 10276 51154
rect 10220 51044 10276 51102
rect 10220 50978 10276 50988
rect 10444 51154 10500 51166
rect 10444 51102 10446 51154
rect 10498 51102 10500 51154
rect 9996 50484 10052 50494
rect 9324 50372 9492 50428
rect 8652 48962 8708 48972
rect 8764 49698 8820 49710
rect 8764 49646 8766 49698
rect 8818 49646 8820 49698
rect 8764 48804 8820 49646
rect 8428 48802 8820 48804
rect 8428 48750 8430 48802
rect 8482 48750 8820 48802
rect 8428 48748 8820 48750
rect 7084 48412 7812 48468
rect 7084 47458 7140 48412
rect 7868 48356 7924 48366
rect 7868 48262 7924 48300
rect 7532 48244 7588 48254
rect 8092 48244 8148 48254
rect 7532 48242 7700 48244
rect 7532 48190 7534 48242
rect 7586 48190 7700 48242
rect 7532 48188 7700 48190
rect 7532 48178 7588 48188
rect 7084 47406 7086 47458
rect 7138 47406 7140 47458
rect 7084 47394 7140 47406
rect 7532 47346 7588 47358
rect 7532 47294 7534 47346
rect 7586 47294 7588 47346
rect 6972 47236 7028 47246
rect 6860 47234 7028 47236
rect 6860 47182 6974 47234
rect 7026 47182 7028 47234
rect 6860 47180 7028 47182
rect 6860 47068 6916 47180
rect 6972 47170 7028 47180
rect 6524 47012 6692 47068
rect 6860 47012 7140 47068
rect 6412 46786 6468 46798
rect 6412 46734 6414 46786
rect 6466 46734 6468 46786
rect 6412 46676 6468 46734
rect 6412 46610 6468 46620
rect 6188 45838 6190 45890
rect 6242 45838 6244 45890
rect 6188 45826 6244 45838
rect 6300 46450 6356 46462
rect 6300 46398 6302 46450
rect 6354 46398 6356 46450
rect 5852 45780 5908 45790
rect 5852 45686 5908 45724
rect 6300 45444 6356 46398
rect 6636 46450 6692 47012
rect 6636 46398 6638 46450
rect 6690 46398 6692 46450
rect 5628 45278 5630 45330
rect 5682 45278 5684 45330
rect 5628 45266 5684 45278
rect 5740 45388 6356 45444
rect 6412 46114 6468 46126
rect 6412 46062 6414 46114
rect 6466 46062 6468 46114
rect 5628 44324 5684 44334
rect 5516 44322 5684 44324
rect 5516 44270 5630 44322
rect 5682 44270 5684 44322
rect 5516 44268 5684 44270
rect 5068 43762 5236 43764
rect 5068 43710 5070 43762
rect 5122 43710 5236 43762
rect 5068 43708 5236 43710
rect 5292 44100 5348 44110
rect 5068 43698 5124 43708
rect 4956 43598 4958 43650
rect 5010 43598 5012 43650
rect 4956 43586 5012 43598
rect 5292 43540 5348 44044
rect 5628 43764 5684 44268
rect 5628 43698 5684 43708
rect 5068 43484 5348 43540
rect 5516 43540 5572 43550
rect 5068 43428 5124 43484
rect 4732 42866 4900 42868
rect 4732 42814 4734 42866
rect 4786 42814 4900 42866
rect 4732 42812 4900 42814
rect 4956 43372 5124 43428
rect 3948 42802 4004 42812
rect 4732 42802 4788 42812
rect 3836 42588 4452 42644
rect 4396 42194 4452 42588
rect 4396 42142 4398 42194
rect 4450 42142 4452 42194
rect 4396 42130 4452 42142
rect 3164 41860 3220 41870
rect 3164 41766 3220 41804
rect 2828 41748 2884 41758
rect 2492 41746 2884 41748
rect 2492 41694 2830 41746
rect 2882 41694 2884 41746
rect 2492 41692 2884 41694
rect 2492 41298 2548 41692
rect 2828 41682 2884 41692
rect 2492 41246 2494 41298
rect 2546 41246 2548 41298
rect 2492 41234 2548 41246
rect 1820 41186 1876 41198
rect 1820 41134 1822 41186
rect 1874 41134 1876 41186
rect 1820 38834 1876 41134
rect 2492 40628 2548 40638
rect 2492 38946 2548 40572
rect 3388 39284 3444 41916
rect 3724 41906 3780 41916
rect 3836 41970 3892 41982
rect 3836 41918 3838 41970
rect 3890 41918 3892 41970
rect 3836 41412 3892 41918
rect 4060 41972 4116 41982
rect 4060 41878 4116 41916
rect 4732 41972 4788 41982
rect 4956 41972 5012 43372
rect 5516 42644 5572 43484
rect 5740 43538 5796 45388
rect 5964 45218 6020 45230
rect 5964 45166 5966 45218
rect 6018 45166 6020 45218
rect 5964 44436 6020 45166
rect 6412 45220 6468 46062
rect 6412 45154 6468 45164
rect 6524 45780 6580 45790
rect 5964 44370 6020 44380
rect 6412 44210 6468 44222
rect 6412 44158 6414 44210
rect 6466 44158 6468 44210
rect 6412 43876 6468 44158
rect 5852 43820 6468 43876
rect 5852 43762 5908 43820
rect 5852 43710 5854 43762
rect 5906 43710 5908 43762
rect 5852 43698 5908 43710
rect 5740 43486 5742 43538
rect 5794 43486 5796 43538
rect 5740 43474 5796 43486
rect 5628 43428 5684 43438
rect 5628 43092 5684 43372
rect 5852 43316 5908 43326
rect 5852 43222 5908 43260
rect 5628 43036 5908 43092
rect 5852 42754 5908 43036
rect 6524 42866 6580 45724
rect 6636 45444 6692 46398
rect 7084 45890 7140 47012
rect 7084 45838 7086 45890
rect 7138 45838 7140 45890
rect 7084 45826 7140 45838
rect 7532 46676 7588 47294
rect 6636 45388 6804 45444
rect 6636 43540 6692 43550
rect 6636 43446 6692 43484
rect 6748 42980 6804 45388
rect 7308 44436 7364 44446
rect 7532 44436 7588 46620
rect 7364 44380 7588 44436
rect 7644 46564 7700 48188
rect 8092 48150 8148 48188
rect 8092 47460 8148 47470
rect 8428 47460 8484 48748
rect 8652 48244 8708 48254
rect 8652 48150 8708 48188
rect 8764 48132 8820 48142
rect 8764 48038 8820 48076
rect 8988 48020 9044 48030
rect 8988 47926 9044 47964
rect 8876 47572 8932 47582
rect 8876 47478 8932 47516
rect 8092 47458 8484 47460
rect 8092 47406 8094 47458
rect 8146 47406 8484 47458
rect 8092 47404 8484 47406
rect 7756 46564 7812 46574
rect 7644 46562 7812 46564
rect 7644 46510 7758 46562
rect 7810 46510 7812 46562
rect 7644 46508 7812 46510
rect 7644 45892 7700 46508
rect 7756 46498 7812 46508
rect 7980 45892 8036 45902
rect 8092 45892 8148 47404
rect 7644 45890 8148 45892
rect 7644 45838 7982 45890
rect 8034 45838 8148 45890
rect 7644 45836 8148 45838
rect 7644 45666 7700 45836
rect 7980 45826 8036 45836
rect 7644 45614 7646 45666
rect 7698 45614 7700 45666
rect 7196 42980 7252 42990
rect 6748 42978 7252 42980
rect 6748 42926 7198 42978
rect 7250 42926 7252 42978
rect 6748 42924 7252 42926
rect 7196 42914 7252 42924
rect 6524 42814 6526 42866
rect 6578 42814 6580 42866
rect 6524 42802 6580 42814
rect 5852 42702 5854 42754
rect 5906 42702 5908 42754
rect 5852 42690 5908 42702
rect 6636 42754 6692 42766
rect 6636 42702 6638 42754
rect 6690 42702 6692 42754
rect 5628 42644 5684 42654
rect 5516 42588 5628 42644
rect 5628 42550 5684 42588
rect 6300 42642 6356 42654
rect 6300 42590 6302 42642
rect 6354 42590 6356 42642
rect 4732 41878 4788 41916
rect 4844 41970 5012 41972
rect 4844 41918 4958 41970
rect 5010 41918 5012 41970
rect 4844 41916 5012 41918
rect 3948 41860 4004 41870
rect 3948 41766 4004 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4844 41412 4900 41916
rect 4956 41906 5012 41916
rect 5068 42530 5124 42542
rect 5068 42478 5070 42530
rect 5122 42478 5124 42530
rect 3836 41356 4900 41412
rect 4620 41298 4676 41356
rect 4620 41246 4622 41298
rect 4674 41246 4676 41298
rect 4620 41234 4676 41246
rect 5068 41298 5124 42478
rect 5292 41972 5348 41982
rect 5292 41878 5348 41916
rect 5964 41972 6020 41982
rect 5852 41858 5908 41870
rect 5852 41806 5854 41858
rect 5906 41806 5908 41858
rect 5628 41746 5684 41758
rect 5628 41694 5630 41746
rect 5682 41694 5684 41746
rect 5628 41412 5684 41694
rect 5068 41246 5070 41298
rect 5122 41246 5124 41298
rect 4508 40628 4564 40638
rect 4508 40534 4564 40572
rect 4844 40404 4900 40414
rect 4620 40292 4676 40302
rect 4620 40198 4676 40236
rect 4844 40290 4900 40348
rect 4844 40238 4846 40290
rect 4898 40238 4900 40290
rect 4844 40226 4900 40238
rect 4508 40180 4564 40190
rect 4284 40178 4564 40180
rect 4284 40126 4510 40178
rect 4562 40126 4564 40178
rect 4284 40124 4564 40126
rect 4284 39620 4340 40124
rect 4508 40114 4564 40124
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5068 39730 5124 41246
rect 5516 41356 5628 41412
rect 5516 40292 5572 41356
rect 5628 41346 5684 41356
rect 5852 41076 5908 41806
rect 5964 41186 6020 41916
rect 5964 41134 5966 41186
rect 6018 41134 6020 41186
rect 5964 41122 6020 41134
rect 6188 41188 6244 41198
rect 6188 41094 6244 41132
rect 5516 40226 5572 40236
rect 5628 40292 5684 40302
rect 5852 40292 5908 41020
rect 5628 40290 5908 40292
rect 5628 40238 5630 40290
rect 5682 40238 5908 40290
rect 5628 40236 5908 40238
rect 5964 40292 6020 40302
rect 5628 40226 5684 40236
rect 5068 39678 5070 39730
rect 5122 39678 5124 39730
rect 4284 39564 4452 39620
rect 3388 39218 3444 39228
rect 4060 39394 4116 39406
rect 4060 39342 4062 39394
rect 4114 39342 4116 39394
rect 2492 38894 2494 38946
rect 2546 38894 2548 38946
rect 2492 38882 2548 38894
rect 1820 38782 1822 38834
rect 1874 38782 1876 38834
rect 1820 38052 1876 38782
rect 4060 38668 4116 39342
rect 1820 37958 1876 37996
rect 3836 38612 4116 38668
rect 4172 39394 4228 39406
rect 4172 39342 4174 39394
rect 4226 39342 4228 39394
rect 2492 37940 2548 37950
rect 2492 37846 2548 37884
rect 3500 37940 3556 37950
rect 3500 37490 3556 37884
rect 3500 37438 3502 37490
rect 3554 37438 3556 37490
rect 3500 37426 3556 37438
rect 3724 37492 3780 37502
rect 3724 37378 3780 37436
rect 3724 37326 3726 37378
rect 3778 37326 3780 37378
rect 3724 37314 3780 37326
rect 3388 37268 3444 37278
rect 3388 37174 3444 37212
rect 3836 37268 3892 38612
rect 3948 37380 4004 37390
rect 4172 37380 4228 39342
rect 4284 39396 4340 39406
rect 4284 39302 4340 39340
rect 4396 38668 4452 39564
rect 4732 39618 4788 39630
rect 4732 39566 4734 39618
rect 4786 39566 4788 39618
rect 4732 39284 4788 39566
rect 4732 39218 4788 39228
rect 4844 38948 4900 38958
rect 4284 38612 4452 38668
rect 4620 38722 4676 38734
rect 4620 38670 4622 38722
rect 4674 38670 4676 38722
rect 4620 38668 4676 38670
rect 4844 38668 4900 38892
rect 4620 38612 4900 38668
rect 4284 37492 4340 38612
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4620 38164 4676 38174
rect 4620 38070 4676 38108
rect 4396 37492 4452 37502
rect 4284 37490 4452 37492
rect 4284 37438 4398 37490
rect 4450 37438 4452 37490
rect 4284 37436 4452 37438
rect 4396 37426 4452 37436
rect 4620 37492 4676 37502
rect 3948 37378 4228 37380
rect 3948 37326 3950 37378
rect 4002 37326 4228 37378
rect 3948 37324 4228 37326
rect 4620 37378 4676 37436
rect 4620 37326 4622 37378
rect 4674 37326 4676 37378
rect 3948 37314 4004 37324
rect 4620 37314 4676 37326
rect 4844 37378 4900 38612
rect 5068 37828 5124 39678
rect 5516 39620 5572 39630
rect 5292 39618 5572 39620
rect 5292 39566 5518 39618
rect 5570 39566 5572 39618
rect 5292 39564 5572 39566
rect 5068 37734 5124 37772
rect 5180 39396 5236 39406
rect 5180 38946 5236 39340
rect 5180 38894 5182 38946
rect 5234 38894 5236 38946
rect 5180 37492 5236 38894
rect 5292 38948 5348 39564
rect 5516 39554 5572 39564
rect 5852 39394 5908 39406
rect 5852 39342 5854 39394
rect 5906 39342 5908 39394
rect 5852 39172 5908 39342
rect 5740 39116 5908 39172
rect 5964 39172 6020 40236
rect 6188 39844 6244 39854
rect 6300 39844 6356 42590
rect 6412 42644 6468 42654
rect 6412 41410 6468 42588
rect 6412 41358 6414 41410
rect 6466 41358 6468 41410
rect 6412 40404 6468 41358
rect 6524 41074 6580 41086
rect 6524 41022 6526 41074
rect 6578 41022 6580 41074
rect 6524 40516 6580 41022
rect 6636 41076 6692 42702
rect 6972 42756 7028 42766
rect 7308 42756 7364 44380
rect 7420 43652 7476 43662
rect 7644 43652 7700 45614
rect 8764 45778 8820 45790
rect 8764 45726 8766 45778
rect 8818 45726 8820 45778
rect 8652 45220 8708 45230
rect 8652 45126 8708 45164
rect 8764 44548 8820 45726
rect 8764 44482 8820 44492
rect 8988 45218 9044 45230
rect 8988 45166 8990 45218
rect 9042 45166 9044 45218
rect 8540 44436 8596 44446
rect 8540 44342 8596 44380
rect 8988 43876 9044 45166
rect 8988 43810 9044 43820
rect 9100 44098 9156 44110
rect 9100 44046 9102 44098
rect 9154 44046 9156 44098
rect 7476 43596 7700 43652
rect 7420 43426 7476 43596
rect 7420 43374 7422 43426
rect 7474 43374 7476 43426
rect 7420 43362 7476 43374
rect 9100 43540 9156 44046
rect 6972 42754 7364 42756
rect 6972 42702 6974 42754
rect 7026 42702 7364 42754
rect 6972 42700 7364 42702
rect 7532 43316 7588 43326
rect 7532 42978 7588 43260
rect 7532 42926 7534 42978
rect 7586 42926 7588 42978
rect 6972 42690 7028 42700
rect 6860 41412 6916 41422
rect 6860 41318 6916 41356
rect 6972 41188 7028 41198
rect 6972 41094 7028 41132
rect 6636 41010 6692 41020
rect 7084 41076 7140 41086
rect 7084 40982 7140 41020
rect 6524 40450 6580 40460
rect 6412 40338 6468 40348
rect 6188 39842 6356 39844
rect 6188 39790 6190 39842
rect 6242 39790 6356 39842
rect 6188 39788 6356 39790
rect 6188 39778 6244 39788
rect 6076 39396 6132 39406
rect 6412 39396 6468 39406
rect 6076 39302 6132 39340
rect 6188 39394 6468 39396
rect 6188 39342 6414 39394
rect 6466 39342 6468 39394
rect 6188 39340 6468 39342
rect 5964 39116 6132 39172
rect 5516 38948 5572 38958
rect 5292 38854 5348 38892
rect 5404 38892 5516 38948
rect 5404 38834 5460 38892
rect 5516 38882 5572 38892
rect 5404 38782 5406 38834
rect 5458 38782 5460 38834
rect 5404 38770 5460 38782
rect 5740 38668 5796 39116
rect 5852 38948 5908 38958
rect 6076 38948 6132 39116
rect 5852 38946 6132 38948
rect 5852 38894 5854 38946
rect 5906 38894 6132 38946
rect 5852 38892 6132 38894
rect 6188 39058 6244 39340
rect 6412 39330 6468 39340
rect 6748 39394 6804 39406
rect 6748 39342 6750 39394
rect 6802 39342 6804 39394
rect 6188 39006 6190 39058
rect 6242 39006 6244 39058
rect 6188 38948 6244 39006
rect 5852 38882 5908 38892
rect 6188 38882 6244 38892
rect 6524 39060 6580 39070
rect 6524 38834 6580 39004
rect 6748 38948 6804 39342
rect 6524 38782 6526 38834
rect 6578 38782 6580 38834
rect 6524 38770 6580 38782
rect 6636 38892 6804 38948
rect 6860 39396 6916 39406
rect 6636 38668 6692 38892
rect 6860 38836 6916 39340
rect 5180 37398 5236 37436
rect 5516 38612 5796 38668
rect 6524 38612 6692 38668
rect 6748 38780 6860 38836
rect 6748 38722 6804 38780
rect 6860 38770 6916 38780
rect 6972 39284 7028 39294
rect 6972 38834 7028 39228
rect 7532 39060 7588 42926
rect 8652 43316 8708 43326
rect 8652 42866 8708 43260
rect 8652 42814 8654 42866
rect 8706 42814 8708 42866
rect 8652 42802 8708 42814
rect 7868 42756 7924 42766
rect 7756 42754 7924 42756
rect 7756 42702 7870 42754
rect 7922 42702 7924 42754
rect 7756 42700 7924 42702
rect 7644 41860 7700 41870
rect 7756 41860 7812 42700
rect 7868 42690 7924 42700
rect 8876 42084 8932 42094
rect 8764 41972 8820 41982
rect 8764 41878 8820 41916
rect 7644 41858 7812 41860
rect 7644 41806 7646 41858
rect 7698 41806 7812 41858
rect 7644 41804 7812 41806
rect 7644 41794 7700 41804
rect 7756 41300 7812 41804
rect 7756 41298 8148 41300
rect 7756 41246 7758 41298
rect 7810 41246 8148 41298
rect 7756 41244 8148 41246
rect 7756 41234 7812 41244
rect 8092 41188 8148 41244
rect 8876 41298 8932 42028
rect 9100 41972 9156 43484
rect 9100 41906 9156 41916
rect 8876 41246 8878 41298
rect 8930 41246 8932 41298
rect 8876 41234 8932 41246
rect 8092 41186 8484 41188
rect 8092 41134 8094 41186
rect 8146 41134 8484 41186
rect 8092 41132 8484 41134
rect 8092 41122 8148 41132
rect 8428 40628 8484 41132
rect 8988 40628 9044 40638
rect 8428 40572 8988 40628
rect 7756 40516 7812 40526
rect 7756 40422 7812 40460
rect 8428 40402 8484 40572
rect 8428 40350 8430 40402
rect 8482 40350 8484 40402
rect 8428 40338 8484 40350
rect 8764 39732 8820 40572
rect 8988 40534 9044 40572
rect 8764 39730 8932 39732
rect 8764 39678 8766 39730
rect 8818 39678 8932 39730
rect 8764 39676 8932 39678
rect 8764 39666 8820 39676
rect 7644 39060 7700 39070
rect 7588 39058 7700 39060
rect 7588 39006 7646 39058
rect 7698 39006 7700 39058
rect 7588 39004 7700 39006
rect 7532 38966 7588 39004
rect 7644 38994 7700 39004
rect 6972 38782 6974 38834
rect 7026 38782 7028 38834
rect 6972 38770 7028 38782
rect 7420 38836 7476 38846
rect 7420 38742 7476 38780
rect 8764 38836 8820 38846
rect 6748 38670 6750 38722
rect 6802 38670 6804 38722
rect 6748 38658 6804 38670
rect 7532 38722 7588 38734
rect 7532 38670 7534 38722
rect 7586 38670 7588 38722
rect 7532 38668 7588 38670
rect 6860 38612 7588 38668
rect 5516 38164 5572 38612
rect 4844 37326 4846 37378
rect 4898 37326 4900 37378
rect 4844 37314 4900 37326
rect 5516 37378 5572 38108
rect 5964 38050 6020 38062
rect 5964 37998 5966 38050
rect 6018 37998 6020 38050
rect 5964 37828 6020 37998
rect 5964 37762 6020 37772
rect 5516 37326 5518 37378
rect 5570 37326 5572 37378
rect 5516 37314 5572 37326
rect 6524 37490 6580 38612
rect 6524 37438 6526 37490
rect 6578 37438 6580 37490
rect 3836 37202 3892 37212
rect 4284 37268 4340 37278
rect 4284 37174 4340 37212
rect 6524 37268 6580 37438
rect 6636 37938 6692 37950
rect 6636 37886 6638 37938
rect 6690 37886 6692 37938
rect 6636 37490 6692 37886
rect 6636 37438 6638 37490
rect 6690 37438 6692 37490
rect 6636 37426 6692 37438
rect 6748 37380 6804 37390
rect 6860 37380 6916 38612
rect 8764 38162 8820 38780
rect 8764 38110 8766 38162
rect 8818 38110 8820 38162
rect 8764 38098 8820 38110
rect 6748 37378 6916 37380
rect 6748 37326 6750 37378
rect 6802 37326 6916 37378
rect 6748 37324 6916 37326
rect 8428 37828 8484 37838
rect 6748 37314 6804 37324
rect 6524 37202 6580 37212
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5740 29426 5796 29438
rect 5740 29374 5742 29426
rect 5794 29374 5796 29426
rect 4284 29316 4340 29326
rect 4060 27860 4116 27870
rect 4284 27860 4340 29260
rect 5740 29316 5796 29374
rect 5740 29250 5796 29260
rect 6412 29316 6468 29326
rect 8316 29316 8372 29326
rect 8428 29316 8484 37772
rect 8876 37828 8932 39676
rect 8876 37762 8932 37772
rect 9212 37828 9268 37838
rect 9212 37734 9268 37772
rect 9436 32788 9492 50372
rect 9996 49810 10052 50428
rect 9996 49758 9998 49810
rect 10050 49758 10052 49810
rect 9996 49746 10052 49758
rect 10444 49812 10500 51102
rect 10556 50034 10612 51324
rect 11004 51314 11060 51324
rect 11340 51378 11396 51436
rect 11676 52052 11732 52062
rect 11676 51490 11732 51996
rect 11676 51438 11678 51490
rect 11730 51438 11732 51490
rect 11676 51426 11732 51438
rect 11340 51326 11342 51378
rect 11394 51326 11396 51378
rect 11340 51314 11396 51326
rect 12124 51378 12180 52780
rect 12460 52276 12516 52894
rect 12796 52948 12852 53790
rect 12908 53058 12964 53900
rect 12908 53006 12910 53058
rect 12962 53006 12964 53058
rect 12908 52994 12964 53006
rect 12460 52210 12516 52220
rect 12572 52388 12628 52398
rect 12572 52162 12628 52332
rect 12572 52110 12574 52162
rect 12626 52110 12628 52162
rect 12572 52098 12628 52110
rect 12796 52162 12852 52892
rect 12796 52110 12798 52162
rect 12850 52110 12852 52162
rect 12796 51490 12852 52110
rect 12796 51438 12798 51490
rect 12850 51438 12852 51490
rect 12796 51426 12852 51438
rect 12908 52162 12964 52174
rect 12908 52110 12910 52162
rect 12962 52110 12964 52162
rect 12124 51326 12126 51378
rect 12178 51326 12180 51378
rect 12124 51314 12180 51326
rect 11340 51156 11396 51166
rect 11340 51062 11396 51100
rect 11788 51156 11844 51166
rect 12012 51156 12068 51166
rect 11788 51154 11956 51156
rect 11788 51102 11790 51154
rect 11842 51102 11956 51154
rect 11788 51100 11956 51102
rect 11788 51090 11844 51100
rect 10892 50706 10948 50718
rect 10892 50654 10894 50706
rect 10946 50654 10948 50706
rect 10892 50484 10948 50654
rect 10892 50418 10948 50428
rect 11228 50594 11284 50606
rect 11228 50542 11230 50594
rect 11282 50542 11284 50594
rect 10556 49982 10558 50034
rect 10610 49982 10612 50034
rect 10556 49970 10612 49982
rect 11004 49812 11060 49822
rect 10444 49810 11060 49812
rect 10444 49758 11006 49810
rect 11058 49758 11060 49810
rect 10444 49756 11060 49758
rect 11004 49746 11060 49756
rect 11228 49810 11284 50542
rect 11788 50484 11844 50494
rect 11788 50390 11844 50428
rect 11228 49758 11230 49810
rect 11282 49758 11284 49810
rect 11228 49700 11284 49758
rect 11228 49634 11284 49644
rect 11676 49700 11732 49710
rect 11676 49606 11732 49644
rect 10220 49588 10276 49598
rect 10892 49588 10948 49598
rect 10220 49586 10948 49588
rect 10220 49534 10222 49586
rect 10274 49534 10894 49586
rect 10946 49534 10948 49586
rect 10220 49532 10948 49534
rect 9772 49026 9828 49038
rect 9996 49028 10052 49038
rect 9772 48974 9774 49026
rect 9826 48974 9828 49026
rect 9660 48914 9716 48926
rect 9660 48862 9662 48914
rect 9714 48862 9716 48914
rect 9660 47572 9716 48862
rect 9772 48916 9828 48974
rect 9772 48850 9828 48860
rect 9884 49026 10052 49028
rect 9884 48974 9998 49026
rect 10050 48974 10052 49026
rect 9884 48972 10052 48974
rect 9772 48244 9828 48254
rect 9772 48150 9828 48188
rect 9884 48132 9940 48972
rect 9996 48962 10052 48972
rect 10220 49028 10276 49532
rect 10892 49522 10948 49532
rect 11788 49028 11844 49038
rect 10220 49026 10388 49028
rect 10220 48974 10222 49026
rect 10274 48974 10388 49026
rect 10220 48972 10388 48974
rect 10220 48962 10276 48972
rect 10332 48466 10388 48972
rect 11004 48804 11060 48814
rect 10332 48414 10334 48466
rect 10386 48414 10388 48466
rect 10332 48402 10388 48414
rect 10892 48802 11060 48804
rect 10892 48750 11006 48802
rect 11058 48750 11060 48802
rect 10892 48748 11060 48750
rect 9884 48066 9940 48076
rect 10892 48244 10948 48748
rect 11004 48738 11060 48748
rect 11340 48804 11396 48814
rect 11340 48802 11508 48804
rect 11340 48750 11342 48802
rect 11394 48750 11508 48802
rect 11340 48748 11508 48750
rect 11340 48738 11396 48748
rect 11340 48468 11396 48478
rect 11340 48244 11396 48412
rect 9660 47506 9716 47516
rect 9996 48020 10052 48030
rect 9996 45332 10052 47964
rect 10892 47348 10948 48188
rect 11004 48242 11396 48244
rect 11004 48190 11342 48242
rect 11394 48190 11396 48242
rect 11004 48188 11396 48190
rect 11004 47570 11060 48188
rect 11340 48178 11396 48188
rect 11452 48356 11508 48748
rect 11676 48356 11732 48366
rect 11452 48300 11676 48356
rect 11452 47908 11508 48300
rect 11676 48130 11732 48300
rect 11676 48078 11678 48130
rect 11730 48078 11732 48130
rect 11676 48066 11732 48078
rect 11004 47518 11006 47570
rect 11058 47518 11060 47570
rect 11004 47506 11060 47518
rect 11228 47852 11508 47908
rect 10892 47292 11172 47348
rect 11004 46674 11060 46686
rect 11004 46622 11006 46674
rect 11058 46622 11060 46674
rect 10556 46562 10612 46574
rect 10556 46510 10558 46562
rect 10610 46510 10612 46562
rect 10556 46116 10612 46510
rect 10556 46050 10612 46060
rect 10668 46452 10724 46462
rect 11004 46452 11060 46622
rect 10668 46450 11060 46452
rect 10668 46398 10670 46450
rect 10722 46398 11060 46450
rect 10668 46396 11060 46398
rect 9996 45330 10388 45332
rect 9996 45278 9998 45330
rect 10050 45278 10388 45330
rect 9996 45276 10388 45278
rect 9996 45266 10052 45276
rect 10108 44548 10164 44558
rect 10332 44548 10388 45276
rect 10556 45220 10612 45230
rect 10556 44994 10612 45164
rect 10668 45106 10724 46396
rect 10892 46116 10948 46126
rect 10892 46002 10948 46060
rect 10892 45950 10894 46002
rect 10946 45950 10948 46002
rect 10892 45938 10948 45950
rect 11116 46004 11172 47292
rect 11228 46674 11284 47852
rect 11228 46622 11230 46674
rect 11282 46622 11284 46674
rect 11228 46610 11284 46622
rect 11564 46676 11620 46686
rect 11564 46582 11620 46620
rect 11788 46564 11844 48972
rect 11900 48916 11956 51100
rect 12012 51062 12068 51100
rect 12908 50708 12964 52110
rect 12908 50642 12964 50652
rect 13132 52164 13188 52174
rect 13356 52164 13412 54348
rect 15148 54402 15428 54404
rect 15148 54350 15374 54402
rect 15426 54350 15428 54402
rect 15148 54348 15428 54350
rect 13468 53956 13524 53966
rect 13468 53862 13524 53900
rect 13580 53844 13636 53854
rect 13580 53750 13636 53788
rect 13692 53506 13748 53518
rect 13692 53454 13694 53506
rect 13746 53454 13748 53506
rect 13468 52946 13524 52958
rect 13468 52894 13470 52946
rect 13522 52894 13524 52946
rect 13468 52836 13524 52894
rect 13468 52770 13524 52780
rect 13580 52834 13636 52846
rect 13580 52782 13582 52834
rect 13634 52782 13636 52834
rect 13356 52108 13524 52164
rect 13132 51490 13188 52108
rect 13132 51438 13134 51490
rect 13186 51438 13188 51490
rect 12572 50596 12628 50606
rect 12572 50502 12628 50540
rect 12348 50484 12404 50494
rect 12348 50390 12404 50428
rect 12572 50372 12628 50382
rect 12460 50316 12572 50372
rect 12348 50036 12404 50046
rect 12460 50036 12516 50316
rect 12572 50306 12628 50316
rect 12908 50370 12964 50382
rect 12908 50318 12910 50370
rect 12962 50318 12964 50370
rect 12348 50034 12516 50036
rect 12348 49982 12350 50034
rect 12402 49982 12516 50034
rect 12348 49980 12516 49982
rect 12348 49970 12404 49980
rect 12236 49924 12292 49934
rect 12236 49830 12292 49868
rect 12572 49810 12628 49822
rect 12572 49758 12574 49810
rect 12626 49758 12628 49810
rect 11900 48850 11956 48860
rect 12124 49028 12180 49038
rect 12124 48356 12180 48972
rect 12124 48354 12516 48356
rect 12124 48302 12126 48354
rect 12178 48302 12516 48354
rect 12124 48300 12516 48302
rect 12124 48290 12180 48300
rect 12348 48020 12404 48030
rect 12124 47572 12180 47582
rect 12124 46786 12180 47516
rect 12124 46734 12126 46786
rect 12178 46734 12180 46786
rect 12124 46722 12180 46734
rect 12012 46674 12068 46686
rect 12012 46622 12014 46674
rect 12066 46622 12068 46674
rect 11788 46508 11956 46564
rect 11452 46450 11508 46462
rect 11452 46398 11454 46450
rect 11506 46398 11508 46450
rect 11452 46340 11508 46398
rect 11788 46340 11844 46350
rect 11340 46284 11788 46340
rect 11228 46004 11284 46014
rect 11116 45948 11228 46004
rect 11228 45938 11284 45948
rect 10668 45054 10670 45106
rect 10722 45054 10724 45106
rect 10668 45042 10724 45054
rect 11004 45106 11060 45118
rect 11004 45054 11006 45106
rect 11058 45054 11060 45106
rect 10556 44942 10558 44994
rect 10610 44942 10612 44994
rect 10556 44930 10612 44942
rect 10668 44884 10724 44894
rect 10444 44548 10500 44558
rect 10668 44548 10724 44828
rect 10332 44546 10500 44548
rect 10332 44494 10446 44546
rect 10498 44494 10500 44546
rect 10332 44492 10500 44494
rect 10108 44454 10164 44492
rect 10444 44482 10500 44492
rect 10556 44492 10724 44548
rect 11004 44548 11060 45054
rect 10220 44436 10276 44446
rect 10220 44342 10276 44380
rect 9548 44098 9604 44110
rect 9548 44046 9550 44098
rect 9602 44046 9604 44098
rect 9548 43652 9604 44046
rect 10332 43876 10388 43886
rect 10220 43652 10276 43662
rect 9548 43586 9604 43596
rect 10108 43650 10276 43652
rect 10108 43598 10222 43650
rect 10274 43598 10276 43650
rect 10108 43596 10276 43598
rect 9884 43428 9940 43438
rect 10108 43428 10164 43596
rect 10220 43586 10276 43596
rect 10332 43650 10388 43820
rect 10332 43598 10334 43650
rect 10386 43598 10388 43650
rect 10332 43586 10388 43598
rect 9884 43426 10164 43428
rect 9884 43374 9886 43426
rect 9938 43374 10164 43426
rect 9884 43372 10164 43374
rect 9884 43362 9940 43372
rect 10108 43092 10164 43372
rect 10220 43428 10276 43438
rect 10220 43314 10276 43372
rect 10220 43262 10222 43314
rect 10274 43262 10276 43314
rect 10220 43250 10276 43262
rect 10220 43092 10276 43102
rect 10108 43036 10220 43092
rect 10220 43026 10276 43036
rect 9660 41972 9716 41982
rect 9660 41858 9716 41916
rect 9660 41806 9662 41858
rect 9714 41806 9716 41858
rect 9660 41748 9716 41806
rect 9660 41692 10164 41748
rect 9548 40628 9604 40638
rect 9548 40402 9604 40572
rect 9548 40350 9550 40402
rect 9602 40350 9604 40402
rect 9548 40338 9604 40350
rect 9660 38388 9716 38398
rect 9660 38162 9716 38332
rect 9660 38110 9662 38162
rect 9714 38110 9716 38162
rect 9660 38098 9716 38110
rect 10108 38052 10164 41692
rect 10332 40516 10388 40526
rect 10332 40422 10388 40460
rect 10108 37986 10164 37996
rect 10556 34916 10612 44492
rect 11004 44482 11060 44492
rect 11116 45108 11172 45118
rect 10668 44324 10724 44334
rect 11116 44324 11172 45052
rect 10668 44230 10724 44268
rect 10780 44322 11172 44324
rect 10780 44270 11118 44322
rect 11170 44270 11172 44322
rect 10780 44268 11172 44270
rect 10780 42866 10836 44268
rect 11116 44258 11172 44268
rect 11228 44996 11284 45006
rect 11228 44210 11284 44940
rect 11228 44158 11230 44210
rect 11282 44158 11284 44210
rect 11228 44100 11284 44158
rect 11004 44044 11284 44100
rect 10892 43652 10948 43662
rect 10892 43558 10948 43596
rect 10780 42814 10782 42866
rect 10834 42814 10836 42866
rect 10780 42802 10836 42814
rect 11004 41972 11060 44044
rect 11116 43876 11172 43886
rect 11116 43650 11172 43820
rect 11116 43598 11118 43650
rect 11170 43598 11172 43650
rect 11116 43586 11172 43598
rect 11228 43652 11284 43662
rect 11340 43652 11396 46284
rect 11788 46002 11844 46284
rect 11788 45950 11790 46002
rect 11842 45950 11844 46002
rect 11788 45938 11844 45950
rect 11788 44996 11844 45006
rect 11788 44902 11844 44940
rect 11452 44548 11508 44558
rect 11452 44322 11508 44492
rect 11788 44436 11844 44446
rect 11788 44342 11844 44380
rect 11452 44270 11454 44322
rect 11506 44270 11508 44322
rect 11452 44258 11508 44270
rect 11284 43596 11396 43652
rect 11228 43558 11284 43596
rect 11340 42868 11396 43596
rect 11676 44100 11732 44110
rect 11452 43538 11508 43550
rect 11676 43540 11732 44044
rect 11452 43486 11454 43538
rect 11506 43486 11508 43538
rect 11452 43204 11508 43486
rect 11452 43138 11508 43148
rect 11564 43484 11732 43540
rect 11788 43876 11844 43886
rect 11788 43538 11844 43820
rect 11788 43486 11790 43538
rect 11842 43486 11844 43538
rect 11564 42980 11620 43484
rect 11788 43474 11844 43486
rect 11676 43316 11732 43326
rect 11676 43222 11732 43260
rect 11676 42980 11732 42990
rect 11564 42978 11732 42980
rect 11564 42926 11678 42978
rect 11730 42926 11732 42978
rect 11564 42924 11732 42926
rect 11676 42914 11732 42924
rect 11452 42868 11508 42878
rect 11116 42866 11508 42868
rect 11116 42814 11454 42866
rect 11506 42814 11508 42866
rect 11116 42812 11508 42814
rect 11116 42194 11172 42812
rect 11116 42142 11118 42194
rect 11170 42142 11172 42194
rect 11116 42130 11172 42142
rect 11340 41972 11396 41982
rect 11004 41970 11396 41972
rect 11004 41918 11342 41970
rect 11394 41918 11396 41970
rect 11004 41916 11396 41918
rect 11004 41298 11060 41916
rect 11340 41906 11396 41916
rect 11452 41972 11508 42812
rect 11452 41906 11508 41916
rect 11004 41246 11006 41298
rect 11058 41246 11060 41298
rect 11004 41234 11060 41246
rect 11900 41300 11956 46508
rect 12012 45108 12068 46622
rect 12348 45330 12404 47964
rect 12460 46116 12516 48300
rect 12572 47348 12628 49758
rect 12908 49812 12964 50318
rect 13132 49924 13188 51438
rect 13468 51490 13524 52108
rect 13468 51438 13470 51490
rect 13522 51438 13524 51490
rect 13468 51426 13524 51438
rect 13580 51380 13636 52782
rect 13692 52500 13748 53454
rect 13692 52434 13748 52444
rect 13804 52946 13860 52958
rect 13804 52894 13806 52946
rect 13858 52894 13860 52946
rect 13692 52162 13748 52174
rect 13692 52110 13694 52162
rect 13746 52110 13748 52162
rect 13692 51604 13748 52110
rect 13804 52164 13860 52894
rect 14028 52946 14084 52958
rect 14028 52894 14030 52946
rect 14082 52894 14084 52946
rect 13804 52070 13860 52108
rect 13916 52836 13972 52846
rect 13916 52162 13972 52780
rect 13916 52110 13918 52162
rect 13970 52110 13972 52162
rect 13916 52098 13972 52110
rect 14028 51604 14084 52894
rect 14812 52388 14868 52398
rect 14812 52276 14868 52332
rect 15148 52276 15204 54348
rect 15372 54338 15428 54348
rect 16268 54292 16324 54462
rect 16268 54226 16324 54236
rect 16492 54290 16548 54302
rect 16492 54238 16494 54290
rect 16546 54238 16548 54290
rect 16492 53956 16548 54238
rect 16492 53890 16548 53900
rect 16828 53508 16884 53518
rect 16828 53414 16884 53452
rect 16604 52834 16660 52846
rect 16604 52782 16606 52834
rect 16658 52782 16660 52834
rect 16492 52724 16548 52734
rect 15820 52722 16548 52724
rect 15820 52670 16494 52722
rect 16546 52670 16548 52722
rect 15820 52668 16548 52670
rect 14812 52220 15204 52276
rect 14812 52162 14868 52220
rect 14812 52110 14814 52162
rect 14866 52110 14868 52162
rect 14812 52098 14868 52110
rect 13692 51548 14084 51604
rect 14364 51938 14420 51950
rect 14364 51886 14366 51938
rect 14418 51886 14420 51938
rect 13804 51380 13860 51390
rect 13580 51378 13860 51380
rect 13580 51326 13806 51378
rect 13858 51326 13860 51378
rect 13580 51324 13860 51326
rect 13804 51314 13860 51324
rect 13580 51156 13636 51166
rect 13580 51154 13748 51156
rect 13580 51102 13582 51154
rect 13634 51102 13748 51154
rect 13580 51100 13748 51102
rect 13580 51090 13636 51100
rect 13692 51044 13748 51100
rect 13468 50708 13524 50718
rect 13468 50428 13524 50652
rect 13692 50428 13748 50988
rect 13468 50372 13636 50428
rect 13692 50372 13860 50428
rect 13132 49858 13188 49868
rect 12908 49746 12964 49756
rect 13244 49810 13300 49822
rect 13244 49758 13246 49810
rect 13298 49758 13300 49810
rect 13244 48804 13300 49758
rect 13468 49810 13524 49822
rect 13468 49758 13470 49810
rect 13522 49758 13524 49810
rect 13468 49252 13524 49758
rect 13244 48738 13300 48748
rect 13356 49196 13524 49252
rect 12908 48244 12964 48254
rect 12684 48018 12740 48030
rect 12684 47966 12686 48018
rect 12738 47966 12740 48018
rect 12684 47796 12740 47966
rect 12684 47730 12740 47740
rect 12908 47570 12964 48188
rect 12908 47518 12910 47570
rect 12962 47518 12964 47570
rect 12908 47506 12964 47518
rect 13356 48020 13412 49196
rect 13468 49028 13524 49038
rect 13580 49028 13636 50372
rect 13804 50036 13860 50372
rect 13916 50372 13972 51548
rect 14028 51380 14084 51390
rect 14028 51286 14084 51324
rect 14364 51380 14420 51886
rect 15036 51938 15092 51950
rect 15036 51886 15038 51938
rect 15090 51886 15092 51938
rect 14364 51314 14420 51324
rect 14476 51492 14532 51502
rect 14476 51378 14532 51436
rect 14476 51326 14478 51378
rect 14530 51326 14532 51378
rect 14364 51154 14420 51166
rect 14364 51102 14366 51154
rect 14418 51102 14420 51154
rect 14364 50596 14420 51102
rect 14364 50530 14420 50540
rect 13916 50306 13972 50316
rect 13804 49980 14308 50036
rect 13804 49812 13860 49822
rect 13804 49698 13860 49756
rect 14140 49810 14196 49822
rect 14140 49758 14142 49810
rect 14194 49758 14196 49810
rect 13804 49646 13806 49698
rect 13858 49646 13860 49698
rect 13804 49634 13860 49646
rect 13916 49700 13972 49710
rect 13468 49026 13636 49028
rect 13468 48974 13470 49026
rect 13522 48974 13636 49026
rect 13468 48972 13636 48974
rect 13468 48962 13524 48972
rect 13356 47460 13412 47964
rect 13580 47684 13636 47694
rect 13580 47590 13636 47628
rect 13468 47460 13524 47470
rect 13356 47458 13524 47460
rect 13356 47406 13470 47458
rect 13522 47406 13524 47458
rect 13356 47404 13524 47406
rect 12572 47282 12628 47292
rect 12796 47234 12852 47246
rect 12796 47182 12798 47234
rect 12850 47182 12852 47234
rect 12796 46674 12852 47182
rect 13468 47124 13524 47404
rect 13468 47058 13524 47068
rect 13580 47234 13636 47246
rect 13580 47182 13582 47234
rect 13634 47182 13636 47234
rect 12796 46622 12798 46674
rect 12850 46622 12852 46674
rect 12796 46610 12852 46622
rect 12908 47012 12964 47022
rect 12460 45892 12516 46060
rect 12572 45892 12628 45902
rect 12460 45890 12628 45892
rect 12460 45838 12574 45890
rect 12626 45838 12628 45890
rect 12460 45836 12628 45838
rect 12572 45826 12628 45836
rect 12908 45778 12964 46956
rect 13580 47012 13636 47182
rect 13356 46786 13412 46798
rect 13356 46734 13358 46786
rect 13410 46734 13412 46786
rect 13132 46676 13188 46686
rect 13132 46582 13188 46620
rect 13356 46676 13412 46734
rect 13356 46610 13412 46620
rect 12908 45726 12910 45778
rect 12962 45726 12964 45778
rect 12908 45714 12964 45726
rect 12348 45278 12350 45330
rect 12402 45278 12404 45330
rect 12348 45266 12404 45278
rect 12012 45014 12068 45052
rect 12572 45108 12628 45118
rect 12572 44548 12628 45052
rect 12572 44322 12628 44492
rect 12572 44270 12574 44322
rect 12626 44270 12628 44322
rect 12572 44258 12628 44270
rect 12908 44996 12964 45006
rect 12236 44210 12292 44222
rect 12236 44158 12238 44210
rect 12290 44158 12292 44210
rect 12012 44100 12068 44110
rect 12236 44100 12292 44158
rect 12068 44044 12292 44100
rect 12348 44100 12404 44110
rect 12012 44034 12068 44044
rect 12348 43876 12404 44044
rect 12012 43820 12404 43876
rect 12012 43538 12068 43820
rect 12908 43762 12964 44940
rect 13468 44436 13524 44446
rect 13244 44212 13300 44222
rect 12908 43710 12910 43762
rect 12962 43710 12964 43762
rect 12012 43486 12014 43538
rect 12066 43486 12068 43538
rect 12012 43474 12068 43486
rect 12236 43652 12852 43708
rect 12908 43698 12964 43710
rect 13020 43988 13076 43998
rect 12236 43538 12292 43652
rect 12796 43650 12852 43652
rect 12796 43598 12798 43650
rect 12850 43598 12852 43650
rect 12796 43586 12852 43598
rect 12236 43486 12238 43538
rect 12290 43486 12292 43538
rect 12236 43474 12292 43486
rect 12684 43538 12740 43550
rect 12684 43486 12686 43538
rect 12738 43486 12740 43538
rect 12684 43204 12740 43486
rect 12684 43138 12740 43148
rect 12908 42980 12964 42990
rect 13020 42980 13076 43932
rect 13132 43540 13188 43550
rect 13132 43446 13188 43484
rect 12908 42978 13076 42980
rect 12908 42926 12910 42978
rect 12962 42926 13076 42978
rect 12908 42924 13076 42926
rect 12908 42914 12964 42924
rect 12796 42756 12852 42766
rect 12796 42662 12852 42700
rect 12012 42532 12068 42542
rect 12012 42438 12068 42476
rect 12684 42532 12740 42542
rect 13244 42532 13300 44156
rect 13356 43652 13412 43662
rect 13356 43538 13412 43596
rect 13356 43486 13358 43538
rect 13410 43486 13412 43538
rect 13356 43474 13412 43486
rect 12684 42530 13300 42532
rect 12684 42478 12686 42530
rect 12738 42478 13300 42530
rect 12684 42476 13300 42478
rect 13356 42754 13412 42766
rect 13356 42702 13358 42754
rect 13410 42702 13412 42754
rect 13356 42532 13412 42702
rect 12684 42466 12740 42476
rect 13356 42466 13412 42476
rect 13468 42308 13524 44380
rect 13580 44322 13636 46956
rect 13916 47236 13972 49644
rect 14140 48914 14196 49758
rect 14140 48862 14142 48914
rect 14194 48862 14196 48914
rect 14140 48850 14196 48862
rect 14140 48354 14196 48366
rect 14140 48302 14142 48354
rect 14194 48302 14196 48354
rect 14140 47796 14196 48302
rect 14140 47730 14196 47740
rect 13916 46786 13972 47180
rect 13916 46734 13918 46786
rect 13970 46734 13972 46786
rect 13692 46674 13748 46686
rect 13692 46622 13694 46674
rect 13746 46622 13748 46674
rect 13692 46564 13748 46622
rect 13692 46498 13748 46508
rect 13916 46228 13972 46734
rect 14028 47458 14084 47470
rect 14028 47406 14030 47458
rect 14082 47406 14084 47458
rect 14028 46450 14084 47406
rect 14140 47348 14196 47358
rect 14140 47254 14196 47292
rect 14028 46398 14030 46450
rect 14082 46398 14084 46450
rect 14028 46386 14084 46398
rect 14140 47124 14196 47134
rect 13692 46172 13972 46228
rect 13692 46002 13748 46172
rect 13692 45950 13694 46002
rect 13746 45950 13748 46002
rect 13692 45938 13748 45950
rect 14140 45890 14196 47068
rect 14140 45838 14142 45890
rect 14194 45838 14196 45890
rect 14140 45826 14196 45838
rect 14252 44548 14308 49980
rect 14364 49812 14420 49822
rect 14364 49718 14420 49756
rect 14364 47012 14420 47022
rect 14364 46674 14420 46956
rect 14364 46622 14366 46674
rect 14418 46622 14420 46674
rect 14364 46610 14420 46622
rect 14476 46564 14532 51326
rect 15036 51044 15092 51886
rect 14812 50988 15092 51044
rect 15148 51044 15204 52220
rect 15708 52276 15764 52286
rect 15484 52164 15540 52174
rect 15484 52070 15540 52108
rect 15372 51492 15428 51502
rect 15372 51398 15428 51436
rect 15260 51378 15316 51390
rect 15260 51326 15262 51378
rect 15314 51326 15316 51378
rect 15260 51268 15316 51326
rect 15596 51380 15652 51390
rect 15596 51286 15652 51324
rect 15260 51202 15316 51212
rect 15148 50988 15428 51044
rect 14700 50706 14756 50718
rect 14700 50654 14702 50706
rect 14754 50654 14756 50706
rect 14588 49586 14644 49598
rect 14588 49534 14590 49586
rect 14642 49534 14644 49586
rect 14588 47796 14644 49534
rect 14700 48244 14756 50654
rect 14812 50372 14868 50988
rect 15148 50820 15204 50830
rect 15036 50596 15092 50606
rect 15036 50502 15092 50540
rect 14924 50484 14980 50494
rect 14924 50390 14980 50428
rect 15148 50372 15204 50764
rect 14812 49924 14868 50316
rect 15036 50316 15204 50372
rect 15372 50594 15428 50988
rect 15372 50542 15374 50594
rect 15426 50542 15428 50594
rect 14812 49868 14980 49924
rect 14812 49588 14868 49598
rect 14812 49494 14868 49532
rect 14924 48916 14980 49868
rect 15036 49810 15092 50316
rect 15372 50260 15428 50542
rect 15708 50484 15764 52220
rect 15820 51490 15876 52668
rect 16492 52658 16548 52668
rect 15820 51438 15822 51490
rect 15874 51438 15876 51490
rect 15820 51426 15876 51438
rect 15932 52500 15988 52510
rect 15932 51044 15988 52444
rect 16156 52052 16212 52062
rect 16156 52050 16324 52052
rect 16156 51998 16158 52050
rect 16210 51998 16324 52050
rect 16156 51996 16324 51998
rect 16156 51986 16212 51996
rect 16268 51602 16324 51996
rect 16268 51550 16270 51602
rect 16322 51550 16324 51602
rect 16268 51538 16324 51550
rect 16156 51380 16212 51390
rect 16380 51380 16436 51390
rect 16212 51378 16436 51380
rect 16212 51326 16382 51378
rect 16434 51326 16436 51378
rect 16212 51324 16436 51326
rect 16156 51314 16212 51324
rect 16044 51268 16100 51278
rect 16044 51174 16100 51212
rect 16268 51154 16324 51166
rect 16268 51102 16270 51154
rect 16322 51102 16324 51154
rect 16268 51044 16324 51102
rect 15932 50988 16324 51044
rect 15820 50484 15876 50494
rect 15708 50482 15876 50484
rect 15708 50430 15822 50482
rect 15874 50430 15876 50482
rect 15708 50428 15876 50430
rect 15820 50418 15876 50428
rect 15372 50204 16212 50260
rect 16156 50034 16212 50204
rect 16156 49982 16158 50034
rect 16210 49982 16212 50034
rect 16156 49970 16212 49982
rect 15036 49758 15038 49810
rect 15090 49758 15092 49810
rect 15036 49746 15092 49758
rect 15932 49922 15988 49934
rect 15932 49870 15934 49922
rect 15986 49870 15988 49922
rect 15484 49586 15540 49598
rect 15484 49534 15486 49586
rect 15538 49534 15540 49586
rect 14924 48850 14980 48860
rect 15148 48914 15204 48926
rect 15148 48862 15150 48914
rect 15202 48862 15204 48914
rect 15148 48468 15204 48862
rect 15148 48402 15204 48412
rect 15260 48804 15316 48814
rect 14700 48150 14756 48188
rect 14588 47730 14644 47740
rect 14812 48130 14868 48142
rect 14812 48078 14814 48130
rect 14866 48078 14868 48130
rect 14476 46498 14532 46508
rect 14588 46900 14644 46910
rect 14588 46004 14644 46844
rect 14476 46002 14644 46004
rect 14476 45950 14590 46002
rect 14642 45950 14644 46002
rect 14476 45948 14644 45950
rect 14476 45444 14532 45948
rect 14588 45938 14644 45948
rect 14476 45330 14532 45388
rect 14476 45278 14478 45330
rect 14530 45278 14532 45330
rect 14476 45266 14532 45278
rect 14700 45780 14756 45790
rect 14700 45330 14756 45724
rect 14700 45278 14702 45330
rect 14754 45278 14756 45330
rect 14700 45266 14756 45278
rect 14364 45108 14420 45118
rect 14364 45014 14420 45052
rect 13916 44492 14308 44548
rect 13580 44270 13582 44322
rect 13634 44270 13636 44322
rect 13580 44258 13636 44270
rect 13692 44324 13748 44334
rect 13692 44230 13748 44268
rect 13804 44100 13860 44110
rect 13804 44006 13860 44044
rect 13916 43708 13972 44492
rect 13804 43652 13972 43708
rect 14028 44322 14084 44334
rect 14252 44324 14308 44334
rect 14028 44270 14030 44322
rect 14082 44270 14084 44322
rect 14028 43764 14084 44270
rect 14140 44322 14308 44324
rect 14140 44270 14254 44322
rect 14306 44270 14308 44322
rect 14140 44268 14308 44270
rect 14140 44212 14196 44268
rect 14252 44258 14308 44268
rect 14476 44324 14532 44334
rect 14140 44146 14196 44156
rect 14364 44212 14420 44222
rect 14028 43698 14084 43708
rect 13804 43650 13860 43652
rect 13804 43598 13806 43650
rect 13858 43598 13860 43650
rect 13804 43586 13860 43598
rect 13692 43540 13748 43550
rect 13692 43446 13748 43484
rect 13916 43540 13972 43550
rect 13916 43538 14308 43540
rect 13916 43486 13918 43538
rect 13970 43486 14308 43538
rect 13916 43484 14308 43486
rect 13916 43474 13972 43484
rect 13692 43204 13748 43214
rect 13692 42754 13748 43148
rect 14252 43092 14308 43484
rect 14364 43538 14420 44156
rect 14476 43988 14532 44268
rect 14476 43922 14532 43932
rect 14700 44098 14756 44110
rect 14700 44046 14702 44098
rect 14754 44046 14756 44098
rect 14700 43876 14756 44046
rect 14812 43876 14868 48078
rect 15148 46676 15204 46686
rect 14924 46674 15204 46676
rect 14924 46622 15150 46674
rect 15202 46622 15204 46674
rect 14924 46620 15204 46622
rect 14924 46114 14980 46620
rect 15148 46228 15204 46620
rect 15148 46162 15204 46172
rect 14924 46062 14926 46114
rect 14978 46062 14980 46114
rect 14924 46050 14980 46062
rect 15036 46004 15092 46014
rect 15036 45910 15092 45948
rect 15036 45444 15092 45454
rect 15036 44322 15092 45388
rect 15148 45332 15204 45342
rect 15260 45332 15316 48748
rect 15484 47460 15540 49534
rect 15820 49588 15876 49598
rect 15820 49494 15876 49532
rect 15596 48356 15652 48366
rect 15932 48356 15988 49870
rect 15652 48300 15988 48356
rect 15596 48262 15652 48300
rect 15484 47404 15988 47460
rect 15596 47234 15652 47246
rect 15596 47182 15598 47234
rect 15650 47182 15652 47234
rect 15484 46786 15540 46798
rect 15484 46734 15486 46786
rect 15538 46734 15540 46786
rect 15484 46004 15540 46734
rect 15484 45938 15540 45948
rect 15148 45330 15316 45332
rect 15148 45278 15150 45330
rect 15202 45278 15316 45330
rect 15148 45276 15316 45278
rect 15148 45266 15204 45276
rect 15036 44270 15038 44322
rect 15090 44270 15092 44322
rect 15036 44258 15092 44270
rect 15372 45218 15428 45230
rect 15372 45166 15374 45218
rect 15426 45166 15428 45218
rect 14924 44212 14980 44222
rect 15372 44212 15428 45166
rect 15484 45106 15540 45118
rect 15484 45054 15486 45106
rect 15538 45054 15540 45106
rect 15484 44546 15540 45054
rect 15484 44494 15486 44546
rect 15538 44494 15540 44546
rect 15484 44482 15540 44494
rect 15484 44212 15540 44222
rect 15372 44156 15484 44212
rect 14924 44118 14980 44156
rect 15484 44118 15540 44156
rect 15148 43876 15204 43886
rect 14812 43820 14980 43876
rect 14700 43810 14756 43820
rect 14364 43486 14366 43538
rect 14418 43486 14420 43538
rect 14364 43474 14420 43486
rect 14812 43426 14868 43438
rect 14812 43374 14814 43426
rect 14866 43374 14868 43426
rect 14252 43036 14532 43092
rect 14028 42868 14084 42878
rect 14476 42868 14532 43036
rect 14700 42868 14756 42878
rect 14476 42866 14756 42868
rect 14476 42814 14702 42866
rect 14754 42814 14756 42866
rect 14476 42812 14756 42814
rect 13692 42702 13694 42754
rect 13746 42702 13748 42754
rect 13692 42690 13748 42702
rect 13916 42756 13972 42766
rect 14028 42756 14084 42812
rect 14700 42802 14756 42812
rect 14812 42868 14868 43374
rect 14812 42802 14868 42812
rect 13916 42754 14084 42756
rect 13916 42702 13918 42754
rect 13970 42702 14084 42754
rect 13916 42700 14084 42702
rect 13916 42690 13972 42700
rect 13804 42530 13860 42542
rect 13804 42478 13806 42530
rect 13858 42478 13860 42530
rect 13468 42252 13748 42308
rect 12236 41972 12292 41982
rect 12236 41878 12292 41916
rect 13468 41860 13524 41870
rect 13356 41636 13412 41646
rect 11900 41298 12292 41300
rect 11900 41246 11902 41298
rect 11954 41246 12292 41298
rect 11900 41244 12292 41246
rect 11900 41234 11956 41244
rect 12236 41186 12292 41244
rect 12236 41134 12238 41186
rect 12290 41134 12292 41186
rect 11452 39732 11508 39742
rect 11452 39638 11508 39676
rect 12236 39732 12292 41134
rect 12572 40964 12628 40974
rect 12572 40870 12628 40908
rect 13132 40514 13188 40526
rect 13132 40462 13134 40514
rect 13186 40462 13188 40514
rect 12796 40402 12852 40414
rect 12796 40350 12798 40402
rect 12850 40350 12852 40402
rect 12236 39618 12292 39676
rect 12236 39566 12238 39618
rect 12290 39566 12292 39618
rect 12236 39554 12292 39566
rect 12460 40292 12516 40302
rect 12796 40292 12852 40350
rect 13132 40404 13188 40462
rect 13132 40338 13188 40348
rect 12460 40290 12852 40292
rect 12460 40238 12462 40290
rect 12514 40238 12852 40290
rect 12460 40236 12852 40238
rect 12460 39620 12516 40236
rect 12684 39732 12740 39742
rect 12572 39620 12628 39630
rect 12460 39618 12628 39620
rect 12460 39566 12574 39618
rect 12626 39566 12628 39618
rect 12460 39564 12628 39566
rect 12572 39554 12628 39564
rect 11900 39060 11956 39070
rect 11788 37940 11844 37950
rect 11788 37846 11844 37884
rect 11788 37380 11844 37390
rect 11900 37380 11956 39004
rect 12684 38388 12740 39676
rect 13020 39508 13076 39518
rect 13020 39414 13076 39452
rect 12684 38322 12740 38332
rect 12796 38722 12852 38734
rect 12796 38670 12798 38722
rect 12850 38670 12852 38722
rect 11788 37378 11956 37380
rect 11788 37326 11790 37378
rect 11842 37326 11956 37378
rect 11788 37324 11956 37326
rect 12572 38052 12628 38062
rect 12796 38052 12852 38670
rect 12572 38050 12852 38052
rect 12572 37998 12574 38050
rect 12626 37998 12852 38050
rect 12572 37996 12852 37998
rect 11788 37314 11844 37324
rect 11116 37268 11172 37278
rect 11116 37174 11172 37212
rect 12572 37268 12628 37996
rect 12572 35812 12628 37212
rect 12908 36258 12964 36270
rect 12908 36206 12910 36258
rect 12962 36206 12964 36258
rect 12908 35812 12964 36206
rect 12012 35756 12964 35812
rect 12012 35698 12068 35756
rect 12012 35646 12014 35698
rect 12066 35646 12068 35698
rect 12012 35634 12068 35646
rect 12684 35586 12740 35598
rect 12684 35534 12686 35586
rect 12738 35534 12740 35586
rect 12684 35140 12740 35534
rect 12908 35364 12964 35756
rect 13244 35364 13300 35374
rect 12908 35308 13244 35364
rect 13244 35298 13300 35308
rect 12684 35074 12740 35084
rect 10556 34850 10612 34860
rect 9436 32722 9492 32732
rect 11788 33124 11844 33134
rect 11788 30548 11844 33068
rect 13356 32676 13412 41580
rect 13468 41410 13524 41804
rect 13692 41860 13748 42252
rect 13804 42084 13860 42478
rect 13804 42018 13860 42028
rect 13916 41860 13972 41870
rect 13692 41858 13972 41860
rect 13692 41806 13918 41858
rect 13970 41806 13972 41858
rect 13692 41804 13972 41806
rect 13468 41358 13470 41410
rect 13522 41358 13524 41410
rect 13468 41346 13524 41358
rect 13580 41410 13636 41422
rect 13580 41358 13582 41410
rect 13634 41358 13636 41410
rect 13580 40516 13636 41358
rect 13580 40450 13636 40460
rect 13692 41186 13748 41804
rect 13916 41794 13972 41804
rect 13916 41636 13972 41646
rect 14028 41636 14084 42700
rect 14140 42756 14196 42766
rect 14140 42662 14196 42700
rect 14364 42642 14420 42654
rect 14364 42590 14366 42642
rect 14418 42590 14420 42642
rect 14364 42532 14420 42590
rect 14812 42642 14868 42654
rect 14812 42590 14814 42642
rect 14866 42590 14868 42642
rect 14812 42532 14868 42590
rect 14364 42476 14868 42532
rect 14364 42196 14420 42206
rect 14364 42102 14420 42140
rect 14476 42084 14532 42094
rect 14476 41990 14532 42028
rect 14812 41972 14868 42476
rect 14924 42084 14980 43820
rect 14924 41990 14980 42028
rect 15148 43538 15204 43820
rect 15148 43486 15150 43538
rect 15202 43486 15204 43538
rect 14700 41916 14868 41972
rect 13972 41580 14084 41636
rect 14364 41746 14420 41758
rect 14364 41694 14366 41746
rect 14418 41694 14420 41746
rect 13916 41570 13972 41580
rect 14252 41300 14308 41310
rect 14252 41206 14308 41244
rect 14028 41188 14084 41198
rect 13692 41134 13694 41186
rect 13746 41134 13748 41186
rect 13692 39956 13748 41134
rect 13916 41186 14084 41188
rect 13916 41134 14030 41186
rect 14082 41134 14084 41186
rect 13916 41132 14084 41134
rect 13916 40628 13972 41132
rect 14028 41122 14084 41132
rect 14364 40740 14420 41694
rect 14364 40674 14420 40684
rect 14476 41298 14532 41310
rect 14476 41246 14478 41298
rect 14530 41246 14532 41298
rect 13916 40562 13972 40572
rect 14476 40626 14532 41246
rect 14476 40574 14478 40626
rect 14530 40574 14532 40626
rect 14476 40562 14532 40574
rect 14588 40628 14644 40638
rect 14700 40628 14756 41916
rect 14812 41748 14868 41758
rect 14812 41298 14868 41692
rect 14812 41246 14814 41298
rect 14866 41246 14868 41298
rect 14812 41234 14868 41246
rect 15036 41188 15092 41198
rect 14924 41186 15092 41188
rect 14924 41134 15038 41186
rect 15090 41134 15092 41186
rect 14924 41132 15092 41134
rect 14924 41076 14980 41132
rect 15036 41122 15092 41132
rect 14588 40626 14756 40628
rect 14588 40574 14590 40626
rect 14642 40574 14756 40626
rect 14588 40572 14756 40574
rect 14812 40740 14868 40750
rect 14588 40562 14644 40572
rect 13916 40404 13972 40414
rect 13916 40310 13972 40348
rect 14700 40402 14756 40414
rect 14700 40350 14702 40402
rect 14754 40350 14756 40402
rect 13692 39890 13748 39900
rect 14588 39506 14644 39518
rect 14588 39454 14590 39506
rect 14642 39454 14644 39506
rect 13916 39396 13972 39406
rect 13804 38948 13860 38958
rect 13804 38854 13860 38892
rect 13692 37828 13748 37838
rect 13692 37826 13860 37828
rect 13692 37774 13694 37826
rect 13746 37774 13860 37826
rect 13692 37772 13860 37774
rect 13692 37762 13748 37772
rect 13692 37268 13748 37278
rect 13692 36482 13748 37212
rect 13804 36708 13860 37772
rect 13916 37154 13972 39340
rect 14588 39396 14644 39454
rect 14588 39330 14644 39340
rect 14700 39284 14756 40350
rect 14700 39218 14756 39228
rect 14812 39060 14868 40684
rect 14924 39506 14980 41020
rect 15148 40628 15204 43486
rect 15260 43652 15316 43662
rect 15372 43652 15428 43662
rect 15316 43650 15428 43652
rect 15316 43598 15374 43650
rect 15426 43598 15428 43650
rect 15316 43596 15428 43598
rect 15260 42868 15316 43596
rect 15372 43586 15428 43596
rect 15596 42980 15652 47182
rect 15708 47012 15764 47022
rect 15708 46898 15764 46956
rect 15708 46846 15710 46898
rect 15762 46846 15764 46898
rect 15708 46834 15764 46846
rect 15820 46452 15876 46462
rect 15820 46358 15876 46396
rect 15932 46228 15988 47404
rect 16044 47012 16100 47022
rect 16268 47012 16324 50988
rect 16380 50428 16436 51324
rect 16604 50820 16660 52782
rect 16828 51378 16884 51390
rect 16828 51326 16830 51378
rect 16882 51326 16884 51378
rect 16828 51156 16884 51326
rect 16828 51090 16884 51100
rect 16604 50754 16660 50764
rect 16380 50372 16548 50428
rect 16492 49924 16548 50372
rect 16492 49858 16548 49868
rect 16380 49812 16436 49822
rect 16380 49718 16436 49756
rect 16716 49138 16772 49150
rect 16716 49086 16718 49138
rect 16770 49086 16772 49138
rect 16604 49028 16660 49038
rect 16604 48934 16660 48972
rect 16604 48804 16660 48814
rect 16492 47684 16548 47694
rect 16492 47348 16548 47628
rect 16492 47282 16548 47292
rect 16044 46674 16100 46956
rect 16044 46622 16046 46674
rect 16098 46622 16100 46674
rect 16044 46610 16100 46622
rect 16156 46956 16324 47012
rect 15708 45780 15764 45790
rect 15708 45686 15764 45724
rect 15820 45780 15876 45790
rect 15932 45780 15988 46172
rect 15820 45778 15988 45780
rect 15820 45726 15822 45778
rect 15874 45726 15988 45778
rect 15820 45724 15988 45726
rect 15820 45714 15876 45724
rect 16044 45668 16100 45678
rect 16044 45574 16100 45612
rect 16156 45444 16212 46956
rect 16380 46900 16436 46910
rect 16380 46898 16548 46900
rect 16380 46846 16382 46898
rect 16434 46846 16548 46898
rect 16380 46844 16548 46846
rect 16380 46834 16436 46844
rect 16268 46788 16324 46798
rect 16268 46694 16324 46732
rect 16380 46564 16436 46574
rect 16380 46450 16436 46508
rect 16380 46398 16382 46450
rect 16434 46398 16436 46450
rect 16380 46386 16436 46398
rect 16492 46116 16548 46844
rect 16604 46340 16660 48748
rect 16716 47460 16772 49086
rect 16828 48692 16884 48702
rect 16828 48242 16884 48636
rect 16828 48190 16830 48242
rect 16882 48190 16884 48242
rect 16828 47908 16884 48190
rect 16828 47842 16884 47852
rect 16716 47394 16772 47404
rect 16716 47236 16772 47246
rect 16716 46788 16772 47180
rect 16716 46722 16772 46732
rect 17052 46340 17108 55022
rect 17388 54516 17444 55246
rect 17612 55300 17668 56142
rect 17948 55524 18004 59200
rect 18396 56644 18452 59200
rect 18508 56644 18564 56654
rect 18396 56642 18564 56644
rect 18396 56590 18510 56642
rect 18562 56590 18564 56642
rect 18396 56588 18564 56590
rect 18508 56578 18564 56588
rect 18844 56420 18900 59200
rect 18284 56364 18900 56420
rect 18956 56642 19012 56654
rect 18956 56590 18958 56642
rect 19010 56590 19012 56642
rect 18284 56306 18340 56364
rect 18284 56254 18286 56306
rect 18338 56254 18340 56306
rect 18284 56242 18340 56254
rect 17948 55458 18004 55468
rect 18620 56194 18676 56206
rect 18620 56142 18622 56194
rect 18674 56142 18676 56194
rect 18508 55412 18564 55422
rect 18508 55318 18564 55356
rect 17612 55234 17668 55244
rect 17836 55298 17892 55310
rect 17836 55246 17838 55298
rect 17890 55246 17892 55298
rect 17164 53956 17220 53966
rect 17164 53862 17220 53900
rect 17388 53842 17444 54460
rect 17836 55076 17892 55246
rect 18284 55300 18340 55310
rect 17836 54514 17892 55020
rect 17948 55186 18004 55198
rect 17948 55134 17950 55186
rect 18002 55134 18004 55186
rect 17948 54740 18004 55134
rect 18284 55188 18340 55244
rect 18284 55186 18564 55188
rect 18284 55134 18286 55186
rect 18338 55134 18564 55186
rect 18284 55132 18564 55134
rect 18284 55122 18340 55132
rect 17948 54674 18004 54684
rect 17836 54462 17838 54514
rect 17890 54462 17892 54514
rect 17836 54450 17892 54462
rect 18284 54514 18340 54526
rect 18284 54462 18286 54514
rect 18338 54462 18340 54514
rect 17388 53790 17390 53842
rect 17442 53790 17444 53842
rect 17388 53778 17444 53790
rect 17500 54292 17556 54302
rect 17500 53730 17556 54236
rect 18284 54292 18340 54462
rect 17500 53678 17502 53730
rect 17554 53678 17556 53730
rect 17500 53666 17556 53678
rect 17836 53730 17892 53742
rect 17836 53678 17838 53730
rect 17890 53678 17892 53730
rect 17836 53508 17892 53678
rect 17724 52836 17780 52846
rect 17724 52742 17780 52780
rect 17836 52164 17892 53452
rect 18172 53060 18228 53070
rect 18284 53060 18340 54236
rect 18172 53058 18340 53060
rect 18172 53006 18174 53058
rect 18226 53006 18340 53058
rect 18172 53004 18340 53006
rect 18172 52994 18228 53004
rect 18508 52946 18564 55132
rect 18620 54514 18676 56142
rect 18956 56194 19012 56590
rect 18956 56142 18958 56194
rect 19010 56142 19012 56194
rect 18956 55300 19012 56142
rect 19292 55972 19348 59200
rect 19740 56868 19796 59200
rect 20188 57204 20244 59200
rect 20188 57148 20468 57204
rect 19740 56812 20132 56868
rect 20076 56644 20132 56812
rect 20076 56588 20244 56644
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 20188 56308 20244 56588
rect 20076 56252 20244 56308
rect 19852 56194 19908 56206
rect 19852 56142 19854 56194
rect 19906 56142 19908 56194
rect 19404 55972 19460 55982
rect 19292 55970 19460 55972
rect 19292 55918 19406 55970
rect 19458 55918 19460 55970
rect 19292 55916 19460 55918
rect 19404 55906 19460 55916
rect 19180 55524 19236 55534
rect 19180 55430 19236 55468
rect 19852 55412 19908 56142
rect 19852 55346 19908 55356
rect 20076 56082 20132 56252
rect 20076 56030 20078 56082
rect 20130 56030 20132 56082
rect 20076 55410 20132 56030
rect 20076 55358 20078 55410
rect 20130 55358 20132 55410
rect 20076 55346 20132 55358
rect 18956 55234 19012 55244
rect 20188 55300 20244 55310
rect 19628 55188 19684 55198
rect 18844 55076 18900 55086
rect 18900 55020 19348 55076
rect 18844 54982 18900 55020
rect 19180 54740 19236 54750
rect 18620 54462 18622 54514
rect 18674 54462 18676 54514
rect 18620 53956 18676 54462
rect 18620 53890 18676 53900
rect 19068 54514 19124 54526
rect 19068 54462 19070 54514
rect 19122 54462 19124 54514
rect 18620 53620 18676 53630
rect 18620 53618 18900 53620
rect 18620 53566 18622 53618
rect 18674 53566 18900 53618
rect 18620 53564 18900 53566
rect 18620 53554 18676 53564
rect 18844 53170 18900 53564
rect 18844 53118 18846 53170
rect 18898 53118 18900 53170
rect 18844 53106 18900 53118
rect 18508 52894 18510 52946
rect 18562 52894 18564 52946
rect 18508 52882 18564 52894
rect 18732 52836 18788 52846
rect 18788 52780 19012 52836
rect 18732 52742 18788 52780
rect 17948 52722 18004 52734
rect 17948 52670 17950 52722
rect 18002 52670 18004 52722
rect 17948 52388 18004 52670
rect 17948 52332 18116 52388
rect 17948 52164 18004 52174
rect 17836 52108 17948 52164
rect 17948 52098 18004 52108
rect 17388 51492 17444 51502
rect 17388 51398 17444 51436
rect 17612 51268 17668 51278
rect 17612 51174 17668 51212
rect 17948 51154 18004 51166
rect 17948 51102 17950 51154
rect 18002 51102 18004 51154
rect 17948 50428 18004 51102
rect 17836 50372 18004 50428
rect 17836 50034 17892 50372
rect 17836 49982 17838 50034
rect 17890 49982 17892 50034
rect 17836 49970 17892 49982
rect 17276 49924 17332 49934
rect 17276 49810 17332 49868
rect 17276 49758 17278 49810
rect 17330 49758 17332 49810
rect 17276 49746 17332 49758
rect 17612 49810 17668 49822
rect 17612 49758 17614 49810
rect 17666 49758 17668 49810
rect 17164 49028 17220 49038
rect 17164 48934 17220 48972
rect 17500 48468 17556 48478
rect 17500 48374 17556 48412
rect 17276 48244 17332 48254
rect 17276 48150 17332 48188
rect 17164 47346 17220 47358
rect 17164 47294 17166 47346
rect 17218 47294 17220 47346
rect 17164 47012 17220 47294
rect 17164 46946 17220 46956
rect 17388 46450 17444 46462
rect 17388 46398 17390 46450
rect 17442 46398 17444 46450
rect 17052 46284 17332 46340
rect 16604 46274 16660 46284
rect 16492 46050 16548 46060
rect 17164 46116 17220 46126
rect 17164 46022 17220 46060
rect 17052 45780 17108 45790
rect 15820 45388 16212 45444
rect 16828 45724 17052 45780
rect 15596 42924 15764 42980
rect 15260 42812 15652 42868
rect 15260 42196 15316 42812
rect 15596 42754 15652 42812
rect 15596 42702 15598 42754
rect 15650 42702 15652 42754
rect 15596 42690 15652 42702
rect 15484 42642 15540 42654
rect 15484 42590 15486 42642
rect 15538 42590 15540 42642
rect 15260 42130 15316 42140
rect 15372 42420 15428 42430
rect 15372 41972 15428 42364
rect 15484 42196 15540 42590
rect 15484 42140 15652 42196
rect 15484 41972 15540 41982
rect 15372 41970 15540 41972
rect 15372 41918 15486 41970
rect 15538 41918 15540 41970
rect 15372 41916 15540 41918
rect 15260 41748 15316 41758
rect 15260 41410 15316 41692
rect 15260 41358 15262 41410
rect 15314 41358 15316 41410
rect 15260 41346 15316 41358
rect 15372 41188 15428 41916
rect 15484 41906 15540 41916
rect 15596 41412 15652 42140
rect 15596 41346 15652 41356
rect 15372 41122 15428 41132
rect 15484 41076 15540 41086
rect 15372 40964 15428 40974
rect 15260 40628 15316 40638
rect 15148 40572 15260 40628
rect 15036 40404 15092 40414
rect 15148 40404 15204 40572
rect 15036 40402 15204 40404
rect 15036 40350 15038 40402
rect 15090 40350 15204 40402
rect 15036 40348 15204 40350
rect 15036 40338 15092 40348
rect 14924 39454 14926 39506
rect 14978 39454 14980 39506
rect 14924 39442 14980 39454
rect 14476 39004 14868 39060
rect 15148 39284 15204 39294
rect 15148 39058 15204 39228
rect 15260 39172 15316 40572
rect 15372 40292 15428 40908
rect 15484 40516 15540 41020
rect 15708 41076 15764 42924
rect 15820 42866 15876 45388
rect 16828 45330 16884 45724
rect 17052 45686 17108 45724
rect 16828 45278 16830 45330
rect 16882 45278 16884 45330
rect 16828 45266 16884 45278
rect 17164 45666 17220 45678
rect 17164 45614 17166 45666
rect 17218 45614 17220 45666
rect 17164 45332 17220 45614
rect 17164 45266 17220 45276
rect 17276 45108 17332 46284
rect 17276 45042 17332 45052
rect 15932 44994 15988 45006
rect 15932 44942 15934 44994
rect 15986 44942 15988 44994
rect 15932 44212 15988 44942
rect 16716 44994 16772 45006
rect 16716 44942 16718 44994
rect 16770 44942 16772 44994
rect 15932 44118 15988 44156
rect 16380 44884 16436 44894
rect 16380 43650 16436 44828
rect 16492 44546 16548 44558
rect 16492 44494 16494 44546
rect 16546 44494 16548 44546
rect 16492 44436 16548 44494
rect 16604 44436 16660 44446
rect 16492 44434 16660 44436
rect 16492 44382 16606 44434
rect 16658 44382 16660 44434
rect 16492 44380 16660 44382
rect 16604 44370 16660 44380
rect 16380 43598 16382 43650
rect 16434 43598 16436 43650
rect 16380 43586 16436 43598
rect 16492 44098 16548 44110
rect 16492 44046 16494 44098
rect 16546 44046 16548 44098
rect 16268 43540 16324 43550
rect 16268 43446 16324 43484
rect 16156 43426 16212 43438
rect 16156 43374 16158 43426
rect 16210 43374 16212 43426
rect 15820 42814 15822 42866
rect 15874 42814 15876 42866
rect 15820 42802 15876 42814
rect 16044 42980 16100 42990
rect 16044 42420 16100 42924
rect 16156 42644 16212 43374
rect 16268 42756 16324 42766
rect 16268 42662 16324 42700
rect 16156 42578 16212 42588
rect 16044 42354 16100 42364
rect 16492 42196 16548 44046
rect 16604 43538 16660 43550
rect 16604 43486 16606 43538
rect 16658 43486 16660 43538
rect 16604 42868 16660 43486
rect 16716 43316 16772 44942
rect 17388 44772 17444 46398
rect 17612 46228 17668 49758
rect 17724 49698 17780 49710
rect 17724 49646 17726 49698
rect 17778 49646 17780 49698
rect 17724 48354 17780 49646
rect 17836 48914 17892 48926
rect 17836 48862 17838 48914
rect 17890 48862 17892 48914
rect 17836 48468 17892 48862
rect 17836 48402 17892 48412
rect 17724 48302 17726 48354
rect 17778 48302 17780 48354
rect 17724 48290 17780 48302
rect 17948 48242 18004 48254
rect 17948 48190 17950 48242
rect 18002 48190 18004 48242
rect 17948 48132 18004 48190
rect 17948 48066 18004 48076
rect 17836 47908 17892 47918
rect 17836 47458 17892 47852
rect 17836 47406 17838 47458
rect 17890 47406 17892 47458
rect 17836 47394 17892 47406
rect 17724 46788 17780 46798
rect 17724 46674 17780 46732
rect 17724 46622 17726 46674
rect 17778 46622 17780 46674
rect 17724 46610 17780 46622
rect 17948 46676 18004 46686
rect 17612 46172 17892 46228
rect 17724 45892 17780 45902
rect 17388 44706 17444 44716
rect 17500 45836 17724 45892
rect 16716 43250 16772 43260
rect 16828 44660 16884 44670
rect 16604 42802 16660 42812
rect 16716 42644 16772 42654
rect 15932 42140 16548 42196
rect 16604 42588 16716 42644
rect 15932 41412 15988 42140
rect 16044 41972 16100 41982
rect 16268 41972 16324 41982
rect 16044 41970 16268 41972
rect 16044 41918 16046 41970
rect 16098 41918 16268 41970
rect 16044 41916 16268 41918
rect 16044 41906 16100 41916
rect 16268 41878 16324 41916
rect 16492 41972 16548 41982
rect 16604 41972 16660 42588
rect 16716 42578 16772 42588
rect 16492 41970 16660 41972
rect 16492 41918 16494 41970
rect 16546 41918 16660 41970
rect 16492 41916 16660 41918
rect 16492 41906 16548 41916
rect 16380 41860 16436 41870
rect 16380 41766 16436 41804
rect 16268 41636 16324 41646
rect 16044 41412 16100 41422
rect 15932 41356 16044 41412
rect 16044 41346 16100 41356
rect 16156 41300 16212 41338
rect 16156 41234 16212 41244
rect 15708 41010 15764 41020
rect 16156 41076 16212 41086
rect 15484 40402 15540 40460
rect 15484 40350 15486 40402
rect 15538 40350 15540 40402
rect 15484 40338 15540 40350
rect 15596 40962 15652 40974
rect 16044 40964 16100 40974
rect 15596 40910 15598 40962
rect 15650 40910 15652 40962
rect 15372 40226 15428 40236
rect 15596 40180 15652 40910
rect 15932 40962 16100 40964
rect 15932 40910 16046 40962
rect 16098 40910 16100 40962
rect 15932 40908 16100 40910
rect 15708 40628 15764 40638
rect 15708 40534 15764 40572
rect 15652 40124 15876 40180
rect 15596 40114 15652 40124
rect 15372 39844 15428 39854
rect 15372 39750 15428 39788
rect 15820 39842 15876 40124
rect 15820 39790 15822 39842
rect 15874 39790 15876 39842
rect 15820 39778 15876 39790
rect 15484 39620 15540 39630
rect 15932 39620 15988 40908
rect 16044 40898 16100 40908
rect 16156 40740 16212 41020
rect 16044 40684 16212 40740
rect 16268 40964 16324 41580
rect 16604 41298 16660 41916
rect 16828 41748 16884 44604
rect 17276 44548 17332 44558
rect 17052 44436 17108 44446
rect 17052 44342 17108 44380
rect 17276 44322 17332 44492
rect 17500 44546 17556 45836
rect 17724 45798 17780 45836
rect 17724 45218 17780 45230
rect 17724 45166 17726 45218
rect 17778 45166 17780 45218
rect 17500 44494 17502 44546
rect 17554 44494 17556 44546
rect 17500 44482 17556 44494
rect 17612 45108 17668 45118
rect 17276 44270 17278 44322
rect 17330 44270 17332 44322
rect 17276 43988 17332 44270
rect 17276 43932 17444 43988
rect 17388 43764 17444 43932
rect 17388 43698 17444 43708
rect 16940 43540 16996 43550
rect 16940 43446 16996 43484
rect 17164 43428 17220 43438
rect 17164 43092 17220 43372
rect 17500 43428 17556 43438
rect 17500 43334 17556 43372
rect 16940 43036 17220 43092
rect 17276 43316 17332 43326
rect 17612 43316 17668 45052
rect 17724 44660 17780 45166
rect 17724 44594 17780 44604
rect 17724 44210 17780 44222
rect 17724 44158 17726 44210
rect 17778 44158 17780 44210
rect 17724 43876 17780 44158
rect 17724 43810 17780 43820
rect 17724 43652 17780 43662
rect 17836 43652 17892 46172
rect 17948 45892 18004 46620
rect 18060 46116 18116 52332
rect 18284 52274 18340 52286
rect 18284 52222 18286 52274
rect 18338 52222 18340 52274
rect 18284 51716 18340 52222
rect 18956 52276 19012 52780
rect 19068 52388 19124 54462
rect 19180 53172 19236 54684
rect 19292 54738 19348 55020
rect 19292 54686 19294 54738
rect 19346 54686 19348 54738
rect 19292 54674 19348 54686
rect 19628 54628 19684 55132
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 20188 54738 20244 55244
rect 20412 55186 20468 57148
rect 20636 55972 20692 59200
rect 21196 56082 21252 56094
rect 21196 56030 21198 56082
rect 21250 56030 21252 56082
rect 20748 55972 20804 55982
rect 20636 55970 20804 55972
rect 20636 55918 20750 55970
rect 20802 55918 20804 55970
rect 20636 55916 20804 55918
rect 20748 55906 20804 55916
rect 20412 55134 20414 55186
rect 20466 55134 20468 55186
rect 20412 55122 20468 55134
rect 20188 54686 20190 54738
rect 20242 54686 20244 54738
rect 20188 54674 20244 54686
rect 19740 54628 19796 54638
rect 19628 54626 19796 54628
rect 19628 54574 19742 54626
rect 19794 54574 19796 54626
rect 19628 54572 19796 54574
rect 19740 54562 19796 54572
rect 19516 54516 19572 54526
rect 19516 54422 19572 54460
rect 20972 54404 21028 54414
rect 21196 54404 21252 56030
rect 20972 54402 21252 54404
rect 20972 54350 20974 54402
rect 21026 54350 21252 54402
rect 20972 54348 21252 54350
rect 20748 53842 20804 53854
rect 20748 53790 20750 53842
rect 20802 53790 20804 53842
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19404 53172 19460 53182
rect 19180 53170 19460 53172
rect 19180 53118 19406 53170
rect 19458 53118 19460 53170
rect 19180 53116 19460 53118
rect 19404 53106 19460 53116
rect 19180 52948 19236 52958
rect 19180 52854 19236 52892
rect 19852 52948 19908 52958
rect 19852 52854 19908 52892
rect 20076 52946 20132 52958
rect 20076 52894 20078 52946
rect 20130 52894 20132 52946
rect 19292 52836 19348 52846
rect 19292 52742 19348 52780
rect 19068 52332 19348 52388
rect 18732 52164 18788 52174
rect 18956 52164 19012 52220
rect 19180 52164 19236 52174
rect 18732 52070 18788 52108
rect 18844 52162 19236 52164
rect 18844 52110 19182 52162
rect 19234 52110 19236 52162
rect 18844 52108 19236 52110
rect 18172 51660 18284 51716
rect 18172 50428 18228 51660
rect 18284 51650 18340 51660
rect 18284 51492 18340 51502
rect 18284 51398 18340 51436
rect 18620 51492 18676 51502
rect 18508 51378 18564 51390
rect 18508 51326 18510 51378
rect 18562 51326 18564 51378
rect 18396 51156 18452 51166
rect 18396 50594 18452 51100
rect 18396 50542 18398 50594
rect 18450 50542 18452 50594
rect 18284 50484 18340 50494
rect 18172 50372 18340 50428
rect 18172 49812 18228 49822
rect 18172 47908 18228 49756
rect 18284 48468 18340 50372
rect 18396 49922 18452 50542
rect 18396 49870 18398 49922
rect 18450 49870 18452 49922
rect 18396 49858 18452 49870
rect 18508 50482 18564 51326
rect 18508 50430 18510 50482
rect 18562 50430 18564 50482
rect 18508 49140 18564 50430
rect 18620 50372 18676 51436
rect 18620 49810 18676 50316
rect 18732 50482 18788 50494
rect 18732 50430 18734 50482
rect 18786 50430 18788 50482
rect 18732 50036 18788 50430
rect 18732 49970 18788 49980
rect 18620 49758 18622 49810
rect 18674 49758 18676 49810
rect 18620 49746 18676 49758
rect 18396 48468 18452 48478
rect 18284 48466 18452 48468
rect 18284 48414 18398 48466
rect 18450 48414 18452 48466
rect 18284 48412 18452 48414
rect 18396 48402 18452 48412
rect 18508 48356 18564 49084
rect 18620 48356 18676 48366
rect 18508 48354 18676 48356
rect 18508 48302 18622 48354
rect 18674 48302 18676 48354
rect 18508 48300 18676 48302
rect 18620 48290 18676 48300
rect 18172 47842 18228 47852
rect 18396 48244 18452 48254
rect 18396 48130 18452 48188
rect 18396 48078 18398 48130
rect 18450 48078 18452 48130
rect 18396 47572 18452 48078
rect 18396 47506 18452 47516
rect 18508 47460 18564 47470
rect 18564 47404 18676 47460
rect 18508 47366 18564 47404
rect 18620 46674 18676 47404
rect 18620 46622 18622 46674
rect 18674 46622 18676 46674
rect 18620 46610 18676 46622
rect 18732 46562 18788 46574
rect 18732 46510 18734 46562
rect 18786 46510 18788 46562
rect 18732 46340 18788 46510
rect 18732 46274 18788 46284
rect 18844 46228 18900 52108
rect 19180 52098 19236 52108
rect 19068 51716 19124 51726
rect 19068 51490 19124 51660
rect 19068 51438 19070 51490
rect 19122 51438 19124 51490
rect 19068 51426 19124 51438
rect 18956 51156 19012 51166
rect 18956 51062 19012 51100
rect 18956 50932 19012 50942
rect 18956 50034 19012 50876
rect 19068 50594 19124 50606
rect 19068 50542 19070 50594
rect 19122 50542 19124 50594
rect 19068 50372 19124 50542
rect 19180 50484 19236 50522
rect 19180 50418 19236 50428
rect 19068 50306 19124 50316
rect 18956 49982 18958 50034
rect 19010 49982 19012 50034
rect 18956 49970 19012 49982
rect 19180 48242 19236 48254
rect 19180 48190 19182 48242
rect 19234 48190 19236 48242
rect 18956 47570 19012 47582
rect 18956 47518 18958 47570
rect 19010 47518 19012 47570
rect 18956 46676 19012 47518
rect 19180 47348 19236 48190
rect 19292 47908 19348 52332
rect 19740 52164 19796 52174
rect 19740 52070 19796 52108
rect 20076 52164 20132 52894
rect 20636 52948 20692 52958
rect 20636 52386 20692 52892
rect 20748 52500 20804 53790
rect 20972 53620 21028 54348
rect 21532 53732 21588 59200
rect 21644 55188 21700 55198
rect 21980 55188 22036 59200
rect 22092 56642 22148 56654
rect 22092 56590 22094 56642
rect 22146 56590 22148 56642
rect 22092 56194 22148 56590
rect 22876 56642 22932 59200
rect 22876 56590 22878 56642
rect 22930 56590 22932 56642
rect 22876 56578 22932 56590
rect 23324 56420 23380 59200
rect 22092 56142 22094 56194
rect 22146 56142 22148 56194
rect 22092 56130 22148 56142
rect 22204 56364 23380 56420
rect 23660 56642 23716 56654
rect 23660 56590 23662 56642
rect 23714 56590 23716 56642
rect 21644 55186 22036 55188
rect 21644 55134 21646 55186
rect 21698 55134 22036 55186
rect 21644 55132 22036 55134
rect 22092 55188 22148 55198
rect 22204 55188 22260 56364
rect 23660 56194 23716 56590
rect 24220 56642 24276 59200
rect 24220 56590 24222 56642
rect 24274 56590 24276 56642
rect 24220 56578 24276 56590
rect 24668 56306 24724 59200
rect 24668 56254 24670 56306
rect 24722 56254 24724 56306
rect 24668 56242 24724 56254
rect 23660 56142 23662 56194
rect 23714 56142 23716 56194
rect 23660 56130 23716 56142
rect 22764 56082 22820 56094
rect 22764 56030 22766 56082
rect 22818 56030 22820 56082
rect 22092 55186 22260 55188
rect 22092 55134 22094 55186
rect 22146 55134 22260 55186
rect 22092 55132 22260 55134
rect 22428 55412 22484 55422
rect 22764 55412 22820 56030
rect 25564 55970 25620 59200
rect 25564 55918 25566 55970
rect 25618 55918 25620 55970
rect 25564 55906 25620 55918
rect 22428 55410 22820 55412
rect 22428 55358 22430 55410
rect 22482 55358 22820 55410
rect 22428 55356 22820 55358
rect 21644 55122 21700 55132
rect 22092 55122 22148 55132
rect 21532 53666 21588 53676
rect 22204 53732 22260 53742
rect 22204 53638 22260 53676
rect 20972 53554 21028 53564
rect 22428 53060 22484 55356
rect 25228 55298 25284 55310
rect 25228 55246 25230 55298
rect 25282 55246 25284 55298
rect 24556 55186 24612 55198
rect 24556 55134 24558 55186
rect 24610 55134 24612 55186
rect 24444 54626 24500 54638
rect 24444 54574 24446 54626
rect 24498 54574 24500 54626
rect 23100 54516 23156 54526
rect 23100 54422 23156 54460
rect 23884 54514 23940 54526
rect 23884 54462 23886 54514
rect 23938 54462 23940 54514
rect 23884 54404 23940 54462
rect 24332 54516 24388 54526
rect 24332 54422 24388 54460
rect 23884 54338 23940 54348
rect 24220 54292 24276 54302
rect 23996 54290 24276 54292
rect 23996 54238 24222 54290
rect 24274 54238 24276 54290
rect 23996 54236 24276 54238
rect 23996 53956 24052 54236
rect 24220 54226 24276 54236
rect 23772 53900 24052 53956
rect 23772 53842 23828 53900
rect 23772 53790 23774 53842
rect 23826 53790 23828 53842
rect 23772 53778 23828 53790
rect 22428 52994 22484 53004
rect 22876 53730 22932 53742
rect 22876 53678 22878 53730
rect 22930 53678 22932 53730
rect 22204 52948 22260 52958
rect 20860 52836 20916 52846
rect 20860 52742 20916 52780
rect 20748 52434 20804 52444
rect 20636 52334 20638 52386
rect 20690 52334 20692 52386
rect 20636 52322 20692 52334
rect 20188 52276 20244 52286
rect 20188 52182 20244 52220
rect 20748 52276 20804 52286
rect 20076 52098 20132 52108
rect 20748 52162 20804 52220
rect 20748 52110 20750 52162
rect 20802 52110 20804 52162
rect 20748 52098 20804 52110
rect 20972 52164 21028 52174
rect 20636 52052 20692 52062
rect 20636 51958 20692 51996
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19852 51378 19908 51390
rect 19852 51326 19854 51378
rect 19906 51326 19908 51378
rect 19628 51044 19684 51054
rect 19516 50988 19628 51044
rect 19404 50820 19460 50830
rect 19404 50594 19460 50764
rect 19404 50542 19406 50594
rect 19458 50542 19460 50594
rect 19404 50484 19460 50542
rect 19404 50418 19460 50428
rect 19516 50428 19572 50988
rect 19628 50978 19684 50988
rect 19852 50932 19908 51326
rect 20188 51378 20244 51390
rect 20188 51326 20190 51378
rect 20242 51326 20244 51378
rect 20076 51268 20132 51278
rect 20076 51174 20132 51212
rect 19852 50866 19908 50876
rect 20188 51044 20244 51326
rect 19740 50594 19796 50606
rect 19740 50542 19742 50594
rect 19794 50542 19796 50594
rect 19740 50484 19796 50542
rect 20188 50594 20244 50988
rect 20524 51378 20580 51390
rect 20524 51326 20526 51378
rect 20578 51326 20580 51378
rect 20188 50542 20190 50594
rect 20242 50542 20244 50594
rect 20188 50530 20244 50542
rect 20412 50596 20468 50606
rect 20524 50596 20580 51326
rect 20412 50594 20580 50596
rect 20412 50542 20414 50594
rect 20466 50542 20580 50594
rect 20412 50540 20580 50542
rect 20412 50530 20468 50540
rect 19516 50372 19684 50428
rect 19740 50418 19796 50428
rect 19964 50484 20020 50522
rect 19964 50418 20020 50428
rect 19628 50036 19684 50372
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19404 49980 19684 50036
rect 19404 48468 19460 49980
rect 19628 49924 19684 49980
rect 19628 49868 19796 49924
rect 19516 49812 19572 49822
rect 19516 49718 19572 49756
rect 19740 49810 19796 49868
rect 19740 49758 19742 49810
rect 19794 49758 19796 49810
rect 19740 49746 19796 49758
rect 20076 49812 20132 49822
rect 20524 49812 20580 50540
rect 20076 49810 20580 49812
rect 20076 49758 20078 49810
rect 20130 49758 20526 49810
rect 20578 49758 20580 49810
rect 20076 49756 20580 49758
rect 20076 49746 20132 49756
rect 19628 49700 19684 49710
rect 19628 49606 19684 49644
rect 19964 49140 20020 49150
rect 19964 49046 20020 49084
rect 19628 48916 19684 48926
rect 19628 48468 19684 48860
rect 20188 48916 20244 48926
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19852 48468 19908 48478
rect 19628 48466 19908 48468
rect 19628 48414 19854 48466
rect 19906 48414 19908 48466
rect 19628 48412 19908 48414
rect 19404 48374 19460 48412
rect 19852 48402 19908 48412
rect 20076 48468 20132 48478
rect 20188 48468 20244 48860
rect 20300 48914 20356 49756
rect 20524 49746 20580 49756
rect 20748 49586 20804 49598
rect 20748 49534 20750 49586
rect 20802 49534 20804 49586
rect 20300 48862 20302 48914
rect 20354 48862 20356 48914
rect 20300 48850 20356 48862
rect 20524 49476 20580 49486
rect 20076 48466 20244 48468
rect 20076 48414 20078 48466
rect 20130 48414 20244 48466
rect 20076 48412 20244 48414
rect 20412 48468 20468 48478
rect 20076 48402 20132 48412
rect 20412 48354 20468 48412
rect 20524 48466 20580 49420
rect 20524 48414 20526 48466
rect 20578 48414 20580 48466
rect 20524 48402 20580 48414
rect 20636 49140 20692 49150
rect 20636 48914 20692 49084
rect 20636 48862 20638 48914
rect 20690 48862 20692 48914
rect 20412 48302 20414 48354
rect 20466 48302 20468 48354
rect 20412 48290 20468 48302
rect 19740 48242 19796 48254
rect 19740 48190 19742 48242
rect 19794 48190 19796 48242
rect 19292 47852 19684 47908
rect 19516 47684 19572 47694
rect 19404 47348 19460 47358
rect 18956 46610 19012 46620
rect 19068 47346 19460 47348
rect 19068 47294 19406 47346
rect 19458 47294 19460 47346
rect 19068 47292 19460 47294
rect 18844 46172 19012 46228
rect 18060 46050 18116 46060
rect 18956 46004 19012 46172
rect 19068 46116 19124 47292
rect 19404 47282 19460 47292
rect 19292 46900 19348 46910
rect 19516 46900 19572 47628
rect 19628 47460 19684 47852
rect 19628 47366 19684 47404
rect 19740 47236 19796 48190
rect 19292 46898 19572 46900
rect 19292 46846 19294 46898
rect 19346 46846 19572 46898
rect 19292 46844 19572 46846
rect 19628 47180 19796 47236
rect 20412 47460 20468 47470
rect 19628 46900 19684 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19740 46900 19796 46910
rect 19628 46844 19740 46900
rect 19292 46834 19348 46844
rect 19740 46806 19796 46844
rect 19068 46050 19124 46060
rect 19292 46676 19348 46686
rect 19292 46116 19348 46620
rect 19516 46676 19572 46686
rect 19516 46674 19684 46676
rect 19516 46622 19518 46674
rect 19570 46622 19684 46674
rect 19516 46620 19684 46622
rect 19516 46610 19572 46620
rect 19292 46050 19348 46060
rect 19404 46562 19460 46574
rect 19404 46510 19406 46562
rect 19458 46510 19460 46562
rect 18844 45948 19012 46004
rect 17948 45836 18116 45892
rect 17948 45666 18004 45678
rect 17948 45614 17950 45666
rect 18002 45614 18004 45666
rect 17948 45108 18004 45614
rect 17948 45042 18004 45052
rect 18060 45106 18116 45836
rect 18844 45890 18900 45948
rect 19404 45892 19460 46510
rect 18844 45838 18846 45890
rect 18898 45838 18900 45890
rect 18284 45780 18340 45790
rect 18284 45686 18340 45724
rect 18060 45054 18062 45106
rect 18114 45054 18116 45106
rect 18060 45042 18116 45054
rect 18396 45218 18452 45230
rect 18396 45166 18398 45218
rect 18450 45166 18452 45218
rect 17948 44884 18004 44894
rect 18284 44884 18340 44894
rect 17948 44790 18004 44828
rect 18172 44882 18340 44884
rect 18172 44830 18286 44882
rect 18338 44830 18340 44882
rect 18172 44828 18340 44830
rect 18172 44436 18228 44828
rect 18284 44818 18340 44828
rect 17948 44324 18004 44334
rect 17948 44230 18004 44268
rect 17724 43650 17892 43652
rect 17724 43598 17726 43650
rect 17778 43598 17892 43650
rect 17724 43596 17892 43598
rect 17724 43586 17780 43596
rect 18060 43540 18116 43550
rect 17612 43260 17892 43316
rect 16940 42754 16996 43036
rect 17052 42868 17108 42878
rect 17052 42774 17108 42812
rect 16940 42702 16942 42754
rect 16994 42702 16996 42754
rect 16940 42308 16996 42702
rect 17164 42644 17220 42654
rect 17164 42550 17220 42588
rect 16940 42242 16996 42252
rect 16940 41972 16996 41982
rect 17276 41972 17332 43260
rect 17724 42756 17780 42766
rect 17724 42662 17780 42700
rect 17500 42644 17556 42654
rect 17388 42530 17444 42542
rect 17388 42478 17390 42530
rect 17442 42478 17444 42530
rect 17388 42196 17444 42478
rect 17388 42130 17444 42140
rect 17388 41972 17444 41982
rect 17276 41970 17444 41972
rect 17276 41918 17390 41970
rect 17442 41918 17444 41970
rect 17276 41916 17444 41918
rect 16940 41878 16996 41916
rect 17388 41906 17444 41916
rect 16828 41692 17220 41748
rect 16604 41246 16606 41298
rect 16658 41246 16660 41298
rect 16604 41234 16660 41246
rect 16044 40514 16100 40684
rect 16044 40462 16046 40514
rect 16098 40462 16100 40514
rect 16044 40450 16100 40462
rect 16156 40516 16212 40526
rect 16268 40516 16324 40908
rect 17052 40962 17108 40974
rect 17052 40910 17054 40962
rect 17106 40910 17108 40962
rect 16828 40740 16884 40750
rect 16156 40514 16324 40516
rect 16156 40462 16158 40514
rect 16210 40462 16324 40514
rect 16156 40460 16324 40462
rect 16380 40626 16436 40638
rect 16380 40574 16382 40626
rect 16434 40574 16436 40626
rect 16156 40450 16212 40460
rect 15484 39526 15540 39564
rect 15596 39564 15988 39620
rect 16156 39730 16212 39742
rect 16156 39678 16158 39730
rect 16210 39678 16212 39730
rect 15372 39394 15428 39406
rect 15372 39342 15374 39394
rect 15426 39342 15428 39394
rect 15372 39284 15428 39342
rect 15372 39218 15428 39228
rect 15260 39106 15316 39116
rect 15148 39006 15150 39058
rect 15202 39006 15204 39058
rect 14476 38946 14532 39004
rect 14476 38894 14478 38946
rect 14530 38894 14532 38946
rect 14140 38836 14196 38846
rect 14028 37828 14084 37838
rect 14140 37828 14196 38780
rect 14252 38722 14308 38734
rect 14252 38670 14254 38722
rect 14306 38670 14308 38722
rect 14252 38668 14308 38670
rect 14252 38612 14420 38668
rect 14364 37938 14420 38612
rect 14364 37886 14366 37938
rect 14418 37886 14420 37938
rect 14028 37826 14308 37828
rect 14028 37774 14030 37826
rect 14082 37774 14308 37826
rect 14028 37772 14308 37774
rect 14028 37762 14084 37772
rect 13916 37102 13918 37154
rect 13970 37102 13972 37154
rect 13916 37090 13972 37102
rect 14028 37492 14084 37502
rect 14028 36932 14084 37436
rect 13804 36642 13860 36652
rect 13916 36876 14084 36932
rect 14140 37490 14196 37502
rect 14140 37438 14142 37490
rect 14194 37438 14196 37490
rect 13692 36430 13694 36482
rect 13746 36430 13748 36482
rect 13692 36418 13748 36430
rect 13804 36372 13860 36382
rect 13804 36278 13860 36316
rect 13916 35364 13972 36876
rect 14028 36484 14084 36494
rect 14028 36390 14084 36428
rect 14028 35364 14084 35374
rect 13916 35308 14028 35364
rect 14028 35298 14084 35308
rect 13580 35140 13636 35150
rect 13580 35026 13636 35084
rect 13804 35140 13860 35150
rect 14140 35140 14196 37438
rect 14252 36482 14308 37772
rect 14364 37492 14420 37886
rect 14364 37426 14420 37436
rect 14364 37268 14420 37278
rect 14364 37174 14420 37212
rect 14476 36708 14532 38894
rect 14588 38836 14644 38846
rect 14924 38836 14980 38846
rect 14588 38834 14980 38836
rect 14588 38782 14590 38834
rect 14642 38782 14926 38834
rect 14978 38782 14980 38834
rect 14588 38780 14980 38782
rect 14588 38770 14644 38780
rect 14924 38770 14980 38780
rect 15148 38836 15204 39006
rect 15372 38948 15428 38958
rect 15372 38854 15428 38892
rect 15148 38770 15204 38780
rect 15260 38834 15316 38846
rect 15260 38782 15262 38834
rect 15314 38782 15316 38834
rect 15260 38668 15316 38782
rect 15596 38834 15652 39564
rect 16044 39394 16100 39406
rect 16044 39342 16046 39394
rect 16098 39342 16100 39394
rect 15596 38782 15598 38834
rect 15650 38782 15652 38834
rect 15596 38770 15652 38782
rect 15708 39172 15764 39182
rect 15148 38612 15316 38668
rect 15036 38556 15204 38612
rect 14700 38276 14756 38286
rect 14700 38050 14756 38220
rect 14700 37998 14702 38050
rect 14754 37998 14756 38050
rect 14700 37986 14756 37998
rect 15036 38050 15092 38556
rect 15036 37998 15038 38050
rect 15090 37998 15092 38050
rect 15036 37986 15092 37998
rect 15596 38388 15652 38398
rect 14812 37940 14868 37950
rect 14812 37846 14868 37884
rect 15036 37380 15092 37390
rect 14700 37324 15036 37380
rect 14588 36708 14644 36718
rect 14476 36706 14644 36708
rect 14476 36654 14590 36706
rect 14642 36654 14644 36706
rect 14476 36652 14644 36654
rect 14588 36642 14644 36652
rect 14252 36430 14254 36482
rect 14306 36430 14308 36482
rect 14252 36418 14308 36430
rect 14476 36484 14532 36494
rect 14700 36484 14756 37324
rect 15036 37314 15092 37324
rect 15372 37380 15428 37390
rect 15372 37286 15428 37324
rect 15596 37266 15652 38332
rect 15596 37214 15598 37266
rect 15650 37214 15652 37266
rect 14476 36482 14756 36484
rect 14476 36430 14478 36482
rect 14530 36430 14756 36482
rect 14476 36428 14756 36430
rect 15036 37044 15092 37054
rect 14476 36418 14532 36428
rect 14924 36260 14980 36270
rect 13804 35138 14196 35140
rect 13804 35086 13806 35138
rect 13858 35086 14196 35138
rect 13804 35084 14196 35086
rect 14252 36258 14980 36260
rect 14252 36206 14926 36258
rect 14978 36206 14980 36258
rect 14252 36204 14980 36206
rect 13804 35074 13860 35084
rect 14252 35028 14308 36204
rect 14924 36194 14980 36204
rect 14924 35924 14980 35934
rect 15036 35924 15092 36988
rect 15596 36706 15652 37214
rect 15708 37156 15764 39116
rect 16044 38948 16100 39342
rect 16044 38882 16100 38892
rect 16156 38946 16212 39678
rect 16380 39396 16436 40574
rect 16716 40516 16772 40526
rect 16604 40514 16772 40516
rect 16604 40462 16718 40514
rect 16770 40462 16772 40514
rect 16604 40460 16772 40462
rect 16492 40402 16548 40414
rect 16492 40350 16494 40402
rect 16546 40350 16548 40402
rect 16492 39620 16548 40350
rect 16604 39620 16660 40460
rect 16716 40450 16772 40460
rect 16828 40514 16884 40684
rect 17052 40628 17108 40910
rect 17052 40562 17108 40572
rect 16828 40462 16830 40514
rect 16882 40462 16884 40514
rect 16828 40450 16884 40462
rect 16604 39564 16772 39620
rect 16492 39554 16548 39564
rect 16380 39340 16660 39396
rect 16492 39172 16548 39182
rect 16268 39060 16324 39070
rect 16268 38966 16324 39004
rect 16156 38894 16158 38946
rect 16210 38894 16212 38946
rect 16156 38882 16212 38894
rect 16492 38834 16548 39116
rect 16492 38782 16494 38834
rect 16546 38782 16548 38834
rect 16492 38770 16548 38782
rect 16380 38724 16436 38734
rect 15708 37090 15764 37100
rect 15820 38052 15876 38062
rect 15820 37044 15876 37996
rect 16044 37716 16100 37726
rect 16044 37268 16100 37660
rect 16380 37378 16436 38668
rect 16380 37326 16382 37378
rect 16434 37326 16436 37378
rect 16380 37314 16436 37326
rect 16492 38612 16548 38622
rect 15820 36978 15876 36988
rect 15932 37266 16100 37268
rect 15932 37214 16046 37266
rect 16098 37214 16100 37266
rect 15932 37212 16100 37214
rect 15932 36932 15988 37212
rect 16044 37202 16100 37212
rect 15932 36866 15988 36876
rect 15596 36654 15598 36706
rect 15650 36654 15652 36706
rect 15596 36642 15652 36654
rect 15820 36708 15876 36718
rect 15260 36484 15316 36494
rect 15316 36428 15540 36484
rect 15260 36390 15316 36428
rect 14924 35922 15092 35924
rect 14924 35870 14926 35922
rect 14978 35870 15092 35922
rect 14924 35868 15092 35870
rect 14924 35858 14980 35868
rect 15036 35252 15092 35262
rect 15036 35028 15092 35196
rect 15372 35028 15428 35038
rect 13580 34974 13582 35026
rect 13634 34974 13636 35026
rect 13580 34962 13636 34974
rect 13916 34972 14644 35028
rect 13916 34916 13972 34972
rect 13692 34860 13972 34916
rect 13580 34804 13636 34814
rect 13692 34804 13748 34860
rect 13580 34802 13748 34804
rect 13580 34750 13582 34802
rect 13634 34750 13748 34802
rect 13580 34748 13748 34750
rect 13580 34738 13636 34748
rect 14476 34132 14532 34142
rect 14364 34130 14532 34132
rect 14364 34078 14478 34130
rect 14530 34078 14532 34130
rect 14364 34076 14532 34078
rect 14364 34020 14420 34076
rect 14476 34066 14532 34076
rect 14140 33964 14420 34020
rect 14140 33796 14196 33964
rect 14476 33908 14532 33918
rect 13356 32610 13412 32620
rect 13580 33346 13636 33358
rect 13580 33294 13582 33346
rect 13634 33294 13636 33346
rect 12460 32564 12516 32574
rect 11564 30492 11844 30548
rect 12236 32508 12460 32564
rect 8988 30212 9044 30222
rect 8988 30210 9604 30212
rect 8988 30158 8990 30210
rect 9042 30158 9604 30210
rect 8988 30156 9604 30158
rect 8988 30146 9044 30156
rect 6412 29314 6804 29316
rect 6412 29262 6414 29314
rect 6466 29262 6804 29314
rect 6412 29260 6804 29262
rect 6412 29250 6468 29260
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 6748 28530 6804 29260
rect 8372 29260 8484 29316
rect 8540 29314 8596 29326
rect 8540 29262 8542 29314
rect 8594 29262 8596 29314
rect 7084 28644 7140 28654
rect 7532 28644 7588 28654
rect 7084 28642 7588 28644
rect 7084 28590 7086 28642
rect 7138 28590 7534 28642
rect 7586 28590 7588 28642
rect 7084 28588 7588 28590
rect 7084 28578 7140 28588
rect 7532 28578 7588 28588
rect 7868 28644 7924 28654
rect 7868 28550 7924 28588
rect 6748 28478 6750 28530
rect 6802 28478 6804 28530
rect 6748 28466 6804 28478
rect 8092 28530 8148 28542
rect 8092 28478 8094 28530
rect 8146 28478 8148 28530
rect 7644 27860 7700 27870
rect 4060 27858 4340 27860
rect 4060 27806 4062 27858
rect 4114 27806 4340 27858
rect 4060 27804 4340 27806
rect 4060 27794 4116 27804
rect 4284 24722 4340 27804
rect 7196 27858 7700 27860
rect 7196 27806 7646 27858
rect 7698 27806 7700 27858
rect 7196 27804 7700 27806
rect 4732 27748 4788 27758
rect 4732 27654 4788 27692
rect 5628 27748 5684 27758
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 5628 26962 5684 27692
rect 6860 27748 6916 27758
rect 7196 27748 7252 27804
rect 6860 27746 7252 27748
rect 6860 27694 6862 27746
rect 6914 27694 7252 27746
rect 6860 27692 7252 27694
rect 6860 27682 6916 27692
rect 5964 27636 6020 27646
rect 5964 27074 6020 27580
rect 7308 27636 7364 27646
rect 7308 27542 7364 27580
rect 5964 27022 5966 27074
rect 6018 27022 6020 27074
rect 5964 27010 6020 27022
rect 6972 27188 7028 27198
rect 5628 26910 5630 26962
rect 5682 26910 5684 26962
rect 5628 26898 5684 26910
rect 6972 26290 7028 27132
rect 7532 27186 7588 27804
rect 7644 27794 7700 27804
rect 8092 27858 8148 28478
rect 8092 27806 8094 27858
rect 8146 27806 8148 27858
rect 7532 27134 7534 27186
rect 7586 27134 7588 27186
rect 7532 27122 7588 27134
rect 6972 26238 6974 26290
rect 7026 26238 7028 26290
rect 6972 26226 7028 26238
rect 7084 26850 7140 26862
rect 7084 26798 7086 26850
rect 7138 26798 7140 26850
rect 7084 26628 7140 26798
rect 6636 26068 6692 26078
rect 5964 26066 6692 26068
rect 5964 26014 6638 26066
rect 6690 26014 6692 26066
rect 5964 26012 6692 26014
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 5964 25506 6020 26012
rect 6636 26002 6692 26012
rect 5964 25454 5966 25506
rect 6018 25454 6020 25506
rect 5964 25442 6020 25454
rect 7084 25508 7140 26572
rect 7644 26850 7700 26862
rect 7644 26798 7646 26850
rect 7698 26798 7700 26850
rect 7532 26402 7588 26414
rect 7532 26350 7534 26402
rect 7586 26350 7588 26402
rect 7420 26290 7476 26302
rect 7420 26238 7422 26290
rect 7474 26238 7476 26290
rect 7420 25732 7476 26238
rect 7420 25666 7476 25676
rect 7084 25506 7476 25508
rect 7084 25454 7086 25506
rect 7138 25454 7476 25506
rect 7084 25452 7476 25454
rect 7084 25442 7140 25452
rect 5628 25284 5684 25294
rect 4956 25282 5684 25284
rect 4956 25230 5630 25282
rect 5682 25230 5684 25282
rect 4956 25228 5684 25230
rect 4956 24834 5012 25228
rect 5628 25218 5684 25228
rect 4956 24782 4958 24834
rect 5010 24782 5012 24834
rect 4956 24770 5012 24782
rect 4284 24670 4286 24722
rect 4338 24670 4340 24722
rect 4284 24658 4340 24670
rect 7084 24610 7140 24622
rect 7084 24558 7086 24610
rect 7138 24558 7140 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 7084 24052 7140 24558
rect 7084 23986 7140 23996
rect 7420 24050 7476 25452
rect 7420 23998 7422 24050
rect 7474 23998 7476 24050
rect 7420 23986 7476 23998
rect 7532 24052 7588 26350
rect 7644 26292 7700 26798
rect 8092 26404 8148 27806
rect 8204 27970 8260 27982
rect 8204 27918 8206 27970
rect 8258 27918 8260 27970
rect 8204 27188 8260 27918
rect 8204 27122 8260 27132
rect 8316 26628 8372 29260
rect 8540 28644 8596 29262
rect 8988 29316 9044 29326
rect 8988 29222 9044 29260
rect 8540 27972 8596 28588
rect 8652 28532 8708 28542
rect 8652 28438 8708 28476
rect 8876 27972 8932 27982
rect 8540 27970 8932 27972
rect 8540 27918 8878 27970
rect 8930 27918 8932 27970
rect 8540 27916 8932 27918
rect 8876 27906 8932 27916
rect 9548 27860 9604 30156
rect 9660 30098 9716 30110
rect 9660 30046 9662 30098
rect 9714 30046 9716 30098
rect 9660 29652 9716 30046
rect 9772 29652 9828 29662
rect 9660 29650 9828 29652
rect 9660 29598 9774 29650
rect 9826 29598 9828 29650
rect 9660 29596 9828 29598
rect 9772 29586 9828 29596
rect 10108 29428 10164 29438
rect 10108 29426 10612 29428
rect 10108 29374 10110 29426
rect 10162 29374 10612 29426
rect 10108 29372 10612 29374
rect 10108 29362 10164 29372
rect 10556 28866 10612 29372
rect 10556 28814 10558 28866
rect 10610 28814 10612 28866
rect 10556 28802 10612 28814
rect 10892 28642 10948 28654
rect 10892 28590 10894 28642
rect 10946 28590 10948 28642
rect 10892 28532 10948 28590
rect 9548 27858 9716 27860
rect 9548 27806 9550 27858
rect 9602 27806 9716 27858
rect 9548 27804 9716 27806
rect 9548 27794 9604 27804
rect 8988 27634 9044 27646
rect 8988 27582 8990 27634
rect 9042 27582 9044 27634
rect 8988 26908 9044 27582
rect 8988 26852 9604 26908
rect 8316 26562 8372 26572
rect 8092 26348 8372 26404
rect 7644 26236 8260 26292
rect 7756 25394 7812 25406
rect 7756 25342 7758 25394
rect 7810 25342 7812 25394
rect 7756 24946 7812 25342
rect 7756 24894 7758 24946
rect 7810 24894 7812 24946
rect 7756 24882 7812 24894
rect 8092 25284 8148 25294
rect 8092 24834 8148 25228
rect 8092 24782 8094 24834
rect 8146 24782 8148 24834
rect 8092 24770 8148 24782
rect 7532 23986 7588 23996
rect 7308 23940 7364 23950
rect 7196 23884 7308 23940
rect 4620 23826 4676 23838
rect 4620 23774 4622 23826
rect 4674 23774 4676 23826
rect 4284 23716 4340 23726
rect 3948 23714 4340 23716
rect 3948 23662 4286 23714
rect 4338 23662 4340 23714
rect 3948 23660 4340 23662
rect 2380 23266 2436 23278
rect 2380 23214 2382 23266
rect 2434 23214 2436 23266
rect 2380 22484 2436 23214
rect 3948 23266 4004 23660
rect 4284 23650 4340 23660
rect 4620 23380 4676 23774
rect 4620 23314 4676 23324
rect 6412 23714 6468 23726
rect 6412 23662 6414 23714
rect 6466 23662 6468 23714
rect 3948 23214 3950 23266
rect 4002 23214 4004 23266
rect 3948 23202 4004 23214
rect 2716 23154 2772 23166
rect 2716 23102 2718 23154
rect 2770 23102 2772 23154
rect 2716 22596 2772 23102
rect 3276 23156 3332 23166
rect 3276 23062 3332 23100
rect 5068 23156 5124 23166
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 2716 22530 2772 22540
rect 2492 22484 2548 22494
rect 2380 22482 2548 22484
rect 2380 22430 2494 22482
rect 2546 22430 2548 22482
rect 2380 22428 2548 22430
rect 2492 22418 2548 22428
rect 4620 22482 4676 22494
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 1820 22370 1876 22382
rect 1820 22318 1822 22370
rect 1874 22318 1876 22370
rect 1820 21586 1876 22318
rect 4620 21924 4676 22430
rect 4620 21858 4676 21868
rect 5068 22146 5124 23100
rect 6412 23156 6468 23662
rect 6524 23380 6580 23390
rect 6524 23286 6580 23324
rect 6412 23090 6468 23100
rect 6076 23042 6132 23054
rect 6076 22990 6078 23042
rect 6130 22990 6132 23042
rect 5740 22596 5796 22606
rect 5740 22502 5796 22540
rect 6076 22596 6132 22990
rect 6076 22530 6132 22540
rect 6860 22930 6916 22942
rect 6860 22878 6862 22930
rect 6914 22878 6916 22930
rect 6860 22596 6916 22878
rect 6860 22530 6916 22540
rect 5068 22094 5070 22146
rect 5122 22094 5124 22146
rect 1820 21534 1822 21586
rect 1874 21534 1876 21586
rect 1820 17668 1876 21534
rect 2492 21474 2548 21486
rect 2492 21422 2494 21474
rect 2546 21422 2548 21474
rect 2380 20692 2436 20702
rect 2492 20692 2548 21422
rect 4620 21474 4676 21486
rect 4620 21422 4622 21474
rect 4674 21422 4676 21474
rect 4620 21364 4676 21422
rect 4172 21308 4620 21364
rect 4172 21026 4228 21308
rect 4620 21298 4676 21308
rect 5068 21474 5124 22094
rect 6076 22370 6132 22382
rect 6076 22318 6078 22370
rect 6130 22318 6132 22370
rect 6076 21924 6132 22318
rect 6860 22372 6916 22382
rect 6860 22278 6916 22316
rect 6076 21858 6132 21868
rect 6748 22258 6804 22270
rect 6748 22206 6750 22258
rect 6802 22206 6804 22258
rect 6748 22036 6804 22206
rect 6860 22036 6916 22046
rect 6748 21980 6860 22036
rect 5068 21422 5070 21474
rect 5122 21422 5124 21474
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4172 20974 4174 21026
rect 4226 20974 4228 21026
rect 4172 20962 4228 20974
rect 4956 20802 5012 20814
rect 4956 20750 4958 20802
rect 5010 20750 5012 20802
rect 2380 20690 2548 20692
rect 2380 20638 2382 20690
rect 2434 20638 2548 20690
rect 2380 20636 2548 20638
rect 2716 20692 2772 20702
rect 2380 20626 2436 20636
rect 2716 20598 2772 20636
rect 3836 20692 3892 20702
rect 3836 20598 3892 20636
rect 4732 20692 4788 20702
rect 4732 20598 4788 20636
rect 4956 20468 5012 20750
rect 4956 20402 5012 20412
rect 4844 20020 4900 20030
rect 5068 20020 5124 21422
rect 5964 20692 6020 20702
rect 6748 20692 6804 21980
rect 6860 21970 6916 21980
rect 5964 20690 6580 20692
rect 5964 20638 5966 20690
rect 6018 20638 6580 20690
rect 5964 20636 6580 20638
rect 5964 20626 6020 20636
rect 5628 20580 5684 20590
rect 5516 20578 5684 20580
rect 5516 20526 5630 20578
rect 5682 20526 5684 20578
rect 5516 20524 5684 20526
rect 5516 20130 5572 20524
rect 5628 20514 5684 20524
rect 5516 20078 5518 20130
rect 5570 20078 5572 20130
rect 5516 20066 5572 20078
rect 4844 20018 5124 20020
rect 4844 19966 4846 20018
rect 4898 19966 5124 20018
rect 4844 19964 5124 19966
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 2828 19122 2884 19134
rect 2828 19070 2830 19122
rect 2882 19070 2884 19122
rect 2492 19010 2548 19022
rect 2492 18958 2494 19010
rect 2546 18958 2548 19010
rect 2268 18450 2324 18462
rect 2268 18398 2270 18450
rect 2322 18398 2324 18450
rect 2268 17668 2324 18398
rect 2492 17778 2548 18958
rect 2828 18452 2884 19070
rect 3612 19122 3668 19134
rect 3612 19070 3614 19122
rect 3666 19070 3668 19122
rect 3276 19012 3332 19022
rect 3052 19010 3332 19012
rect 3052 18958 3278 19010
rect 3330 18958 3332 19010
rect 3052 18956 3332 18958
rect 3052 18562 3108 18956
rect 3276 18946 3332 18956
rect 3052 18510 3054 18562
rect 3106 18510 3108 18562
rect 3052 18498 3108 18510
rect 2828 18386 2884 18396
rect 3612 17892 3668 19070
rect 4844 19012 4900 19964
rect 6524 19458 6580 20636
rect 6748 20626 6804 20636
rect 6524 19406 6526 19458
rect 6578 19406 6580 19458
rect 6524 19394 6580 19406
rect 6860 19908 6916 19918
rect 6860 19458 6916 19852
rect 6860 19406 6862 19458
rect 6914 19406 6916 19458
rect 6860 19394 6916 19406
rect 5068 19012 5124 19022
rect 4844 18956 5068 19012
rect 4956 18340 5012 18350
rect 4844 18284 4956 18340
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 3612 17826 3668 17836
rect 2492 17726 2494 17778
rect 2546 17726 2548 17778
rect 2492 17714 2548 17726
rect 4620 17780 4676 17790
rect 4844 17780 4900 18284
rect 4956 18274 5012 18284
rect 4620 17778 4900 17780
rect 4620 17726 4622 17778
rect 4674 17726 4900 17778
rect 4620 17724 4900 17726
rect 4620 17714 4676 17724
rect 1820 17666 2324 17668
rect 1820 17614 1822 17666
rect 1874 17614 2324 17666
rect 1820 17612 2324 17614
rect 1820 17602 1876 17612
rect 1820 16100 1876 16110
rect 2268 16100 2324 17612
rect 5068 17442 5124 18956
rect 5740 19012 5796 19022
rect 5740 18918 5796 18956
rect 6860 18676 6916 18686
rect 6524 18564 6580 18574
rect 6748 18564 6804 18574
rect 6412 18562 6580 18564
rect 6412 18510 6526 18562
rect 6578 18510 6580 18562
rect 6412 18508 6580 18510
rect 5628 18452 5684 18462
rect 5628 18358 5684 18396
rect 5964 18452 6020 18462
rect 5964 18358 6020 18396
rect 5180 18338 5236 18350
rect 5180 18286 5182 18338
rect 5234 18286 5236 18338
rect 5180 17668 5236 18286
rect 5740 17892 5796 17902
rect 5740 17798 5796 17836
rect 6412 17780 6468 18508
rect 6524 18498 6580 18508
rect 6636 18508 6748 18564
rect 6636 18450 6692 18508
rect 6748 18498 6804 18508
rect 6636 18398 6638 18450
rect 6690 18398 6692 18450
rect 6636 18340 6692 18398
rect 6412 17714 6468 17724
rect 6524 18284 6692 18340
rect 6076 17668 6132 17678
rect 5180 17666 6132 17668
rect 5180 17614 6078 17666
rect 6130 17614 6132 17666
rect 5180 17612 6132 17614
rect 5068 17390 5070 17442
rect 5122 17390 5124 17442
rect 2380 16994 2436 17006
rect 2380 16942 2382 16994
rect 2434 16942 2436 16994
rect 2380 16212 2436 16942
rect 2716 16882 2772 16894
rect 2716 16830 2718 16882
rect 2770 16830 2772 16882
rect 2716 16660 2772 16830
rect 2716 16594 2772 16604
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4620 16324 4676 16334
rect 2492 16212 2548 16222
rect 2380 16210 2548 16212
rect 2380 16158 2494 16210
rect 2546 16158 2548 16210
rect 2380 16156 2548 16158
rect 2492 16146 2548 16156
rect 4620 16210 4676 16268
rect 4620 16158 4622 16210
rect 4674 16158 4676 16210
rect 4620 16146 4676 16158
rect 1820 16098 2324 16100
rect 1820 16046 1822 16098
rect 1874 16046 2324 16098
rect 1820 16044 2324 16046
rect 1820 16034 1876 16044
rect 2268 15316 2324 16044
rect 5068 15874 5124 17390
rect 5964 16772 6020 17612
rect 6076 17602 6132 17612
rect 6524 17666 6580 18284
rect 6860 17780 6916 18620
rect 7196 17890 7252 23884
rect 7308 23874 7364 23884
rect 7756 23940 7812 23950
rect 7756 23826 7812 23884
rect 7756 23774 7758 23826
rect 7810 23774 7812 23826
rect 7756 23762 7812 23774
rect 7980 23938 8036 23950
rect 7980 23886 7982 23938
rect 8034 23886 8036 23938
rect 7420 23266 7476 23278
rect 7420 23214 7422 23266
rect 7474 23214 7476 23266
rect 7420 21252 7476 23214
rect 7644 23154 7700 23166
rect 7644 23102 7646 23154
rect 7698 23102 7700 23154
rect 7644 22372 7700 23102
rect 7644 22278 7700 22316
rect 7980 22932 8036 23886
rect 7980 22370 8036 22876
rect 7980 22318 7982 22370
rect 8034 22318 8036 22370
rect 7980 22306 8036 22318
rect 7532 22148 7588 22158
rect 7868 22148 7924 22158
rect 7532 22146 8036 22148
rect 7532 22094 7534 22146
rect 7586 22094 7870 22146
rect 7922 22094 8036 22146
rect 7532 22092 8036 22094
rect 7532 22082 7588 22092
rect 7868 22082 7924 22092
rect 7532 21924 7588 21934
rect 7532 21698 7588 21868
rect 7532 21646 7534 21698
rect 7586 21646 7588 21698
rect 7532 21634 7588 21646
rect 7756 21698 7812 21710
rect 7756 21646 7758 21698
rect 7810 21646 7812 21698
rect 7196 17838 7198 17890
rect 7250 17838 7252 17890
rect 6524 17614 6526 17666
rect 6578 17614 6580 17666
rect 6524 17602 6580 17614
rect 6748 17724 6916 17780
rect 7084 17780 7140 17790
rect 6412 17556 6468 17566
rect 6412 17106 6468 17500
rect 6412 17054 6414 17106
rect 6466 17054 6468 17106
rect 6412 17042 6468 17054
rect 6748 17108 6804 17724
rect 6860 17556 6916 17566
rect 6860 17554 7028 17556
rect 6860 17502 6862 17554
rect 6914 17502 7028 17554
rect 6860 17500 7028 17502
rect 6860 17490 6916 17500
rect 6860 17108 6916 17118
rect 6748 17106 6916 17108
rect 6748 17054 6862 17106
rect 6914 17054 6916 17106
rect 6748 17052 6916 17054
rect 6860 17042 6916 17052
rect 6972 16996 7028 17500
rect 6076 16884 6132 16894
rect 6300 16884 6356 16894
rect 6748 16884 6804 16894
rect 6076 16790 6132 16828
rect 6188 16882 6356 16884
rect 6188 16830 6302 16882
rect 6354 16830 6356 16882
rect 6188 16828 6356 16830
rect 5964 16706 6020 16716
rect 5740 16660 5796 16670
rect 5740 16322 5796 16604
rect 5740 16270 5742 16322
rect 5794 16270 5796 16322
rect 5740 16258 5796 16270
rect 6076 16324 6132 16334
rect 6188 16324 6244 16828
rect 6300 16818 6356 16828
rect 6524 16882 6804 16884
rect 6524 16830 6750 16882
rect 6802 16830 6804 16882
rect 6524 16828 6804 16830
rect 6132 16268 6244 16324
rect 6076 16230 6132 16268
rect 5068 15822 5070 15874
rect 5122 15822 5124 15874
rect 2380 15316 2436 15326
rect 2268 15260 2380 15316
rect 2380 15250 2436 15260
rect 2940 15316 2996 15326
rect 2940 15222 2996 15260
rect 5068 15316 5124 15822
rect 3612 15202 3668 15214
rect 3612 15150 3614 15202
rect 3666 15150 3668 15202
rect 3612 15148 3668 15150
rect 3612 15092 3892 15148
rect 3836 14418 3892 15092
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 5068 14532 5124 15260
rect 5740 15204 5796 15214
rect 6524 15204 6580 16828
rect 6748 16818 6804 16828
rect 6972 16436 7028 16940
rect 5740 15202 6580 15204
rect 5740 15150 5742 15202
rect 5794 15150 6580 15202
rect 5740 15148 6580 15150
rect 5740 15138 5796 15148
rect 5068 14466 5124 14476
rect 5964 14532 6020 14542
rect 5964 14438 6020 14476
rect 3836 14366 3838 14418
rect 3890 14366 3892 14418
rect 3836 14354 3892 14366
rect 4172 14420 4228 14430
rect 4172 14326 4228 14364
rect 6188 14420 6244 14430
rect 6188 13970 6244 14364
rect 6188 13918 6190 13970
rect 6242 13918 6244 13970
rect 6188 13906 6244 13918
rect 2492 13860 2548 13870
rect 3052 13860 3108 13870
rect 2044 12964 2100 12974
rect 1820 12962 2100 12964
rect 1820 12910 2046 12962
rect 2098 12910 2100 12962
rect 1820 12908 2100 12910
rect 1820 12178 1876 12908
rect 2044 12898 2100 12908
rect 2492 12290 2548 13804
rect 2828 13858 3108 13860
rect 2828 13806 3054 13858
rect 3106 13806 3108 13858
rect 2828 13804 3108 13806
rect 2828 13074 2884 13804
rect 3052 13794 3108 13804
rect 3724 13860 3780 13870
rect 3724 13766 3780 13804
rect 3276 13746 3332 13758
rect 3276 13694 3278 13746
rect 3330 13694 3332 13746
rect 3276 13188 3332 13694
rect 3276 13122 3332 13132
rect 4060 13746 4116 13758
rect 4060 13694 4062 13746
rect 4114 13694 4116 13746
rect 2828 13022 2830 13074
rect 2882 13022 2884 13074
rect 2828 13010 2884 13022
rect 4060 12404 4116 13694
rect 6524 13746 6580 15148
rect 6524 13694 6526 13746
rect 6578 13694 6580 13746
rect 6524 13682 6580 13694
rect 6748 16380 7028 16436
rect 6748 15986 6804 16380
rect 6748 15934 6750 15986
rect 6802 15934 6804 15986
rect 5292 13636 5348 13646
rect 5292 13542 5348 13580
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 5740 13188 5796 13198
rect 5740 13094 5796 13132
rect 4956 13074 5012 13086
rect 4956 13022 4958 13074
rect 5010 13022 5012 13074
rect 4956 12964 5012 13022
rect 6412 13076 6468 13086
rect 4956 12898 5012 12908
rect 6076 12964 6132 12974
rect 6076 12870 6132 12908
rect 6412 12852 6468 13020
rect 6188 12850 6468 12852
rect 6188 12798 6414 12850
rect 6466 12798 6468 12850
rect 6188 12796 6468 12798
rect 6748 12852 6804 15934
rect 6860 16098 6916 16110
rect 6860 16046 6862 16098
rect 6914 16046 6916 16098
rect 6860 15988 6916 16046
rect 6860 15922 6916 15932
rect 6972 15316 7028 15326
rect 6972 15222 7028 15260
rect 7084 14756 7140 17724
rect 7196 16324 7252 17838
rect 7308 19124 7364 19134
rect 7308 16884 7364 19068
rect 7420 19122 7476 21196
rect 7644 21364 7700 21374
rect 7644 21026 7700 21308
rect 7644 20974 7646 21026
rect 7698 20974 7700 21026
rect 7644 20962 7700 20974
rect 7756 20804 7812 21646
rect 7868 21476 7924 21486
rect 7980 21476 8036 22092
rect 8204 21698 8260 26236
rect 8316 24050 8372 26348
rect 8876 25620 8932 25630
rect 8876 24834 8932 25564
rect 8876 24782 8878 24834
rect 8930 24782 8932 24834
rect 8876 24770 8932 24782
rect 8988 24498 9044 24510
rect 8988 24446 8990 24498
rect 9042 24446 9044 24498
rect 8316 23998 8318 24050
rect 8370 23998 8372 24050
rect 8316 23986 8372 23998
rect 8652 24052 8708 24062
rect 8652 23958 8708 23996
rect 8988 23828 9044 24446
rect 9212 24052 9268 24062
rect 9212 23958 9268 23996
rect 8988 23772 9268 23828
rect 8764 23716 8820 23726
rect 8764 23714 9156 23716
rect 8764 23662 8766 23714
rect 8818 23662 9156 23714
rect 8764 23660 9156 23662
rect 8764 23650 8820 23660
rect 8988 22820 9044 22830
rect 8652 22596 8708 22606
rect 8652 22502 8708 22540
rect 8988 22370 9044 22764
rect 8988 22318 8990 22370
rect 9042 22318 9044 22370
rect 8988 22306 9044 22318
rect 8764 22146 8820 22158
rect 8764 22094 8766 22146
rect 8818 22094 8820 22146
rect 8764 21812 8820 22094
rect 8764 21746 8820 21756
rect 8988 21810 9044 21822
rect 8988 21758 8990 21810
rect 9042 21758 9044 21810
rect 8204 21646 8206 21698
rect 8258 21646 8260 21698
rect 8204 21634 8260 21646
rect 8876 21700 8932 21710
rect 8540 21588 8596 21598
rect 7980 21420 8260 21476
rect 7868 21382 7924 21420
rect 7980 21028 8036 21066
rect 7980 20962 8036 20972
rect 7980 20804 8036 20814
rect 7756 20802 8036 20804
rect 7756 20750 7982 20802
rect 8034 20750 8036 20802
rect 7756 20748 8036 20750
rect 7756 20468 7812 20478
rect 7644 19908 7700 19918
rect 7644 19814 7700 19852
rect 7420 19070 7422 19122
rect 7474 19070 7476 19122
rect 7420 19058 7476 19070
rect 7532 19796 7588 19806
rect 7532 17108 7588 19740
rect 7644 19236 7700 19246
rect 7756 19236 7812 20412
rect 7980 19796 8036 20748
rect 7980 19730 8036 19740
rect 8092 19906 8148 19918
rect 8092 19854 8094 19906
rect 8146 19854 8148 19906
rect 7644 19234 7812 19236
rect 7644 19182 7646 19234
rect 7698 19182 7812 19234
rect 7644 19180 7812 19182
rect 7644 19170 7700 19180
rect 7980 19010 8036 19022
rect 7980 18958 7982 19010
rect 8034 18958 8036 19010
rect 7980 18564 8036 18958
rect 8092 19012 8148 19854
rect 8092 18946 8148 18956
rect 8204 19348 8260 21420
rect 8540 21252 8596 21532
rect 8876 21586 8932 21644
rect 8876 21534 8878 21586
rect 8930 21534 8932 21586
rect 8652 21476 8708 21486
rect 8652 21382 8708 21420
rect 8540 21196 8708 21252
rect 8540 21028 8596 21066
rect 8540 20962 8596 20972
rect 8204 19122 8260 19292
rect 8540 20804 8596 20814
rect 8204 19070 8206 19122
rect 8258 19070 8260 19122
rect 8204 18900 8260 19070
rect 8316 19124 8372 19134
rect 8316 19030 8372 19068
rect 8204 18844 8484 18900
rect 7980 18498 8036 18508
rect 8428 18450 8484 18844
rect 8540 18676 8596 20748
rect 8652 20692 8708 21196
rect 8876 20916 8932 21534
rect 8988 21028 9044 21758
rect 8988 20962 9044 20972
rect 8876 20850 8932 20860
rect 9100 20802 9156 23660
rect 9100 20750 9102 20802
rect 9154 20750 9156 20802
rect 9100 20738 9156 20750
rect 8876 20692 8932 20702
rect 8652 20690 8932 20692
rect 8652 20638 8878 20690
rect 8930 20638 8932 20690
rect 8652 20636 8932 20638
rect 8764 19908 8820 19918
rect 8652 19906 8820 19908
rect 8652 19854 8766 19906
rect 8818 19854 8820 19906
rect 8652 19852 8820 19854
rect 8652 19124 8708 19852
rect 8764 19842 8820 19852
rect 8876 19684 8932 20636
rect 8988 20578 9044 20590
rect 8988 20526 8990 20578
rect 9042 20526 9044 20578
rect 8988 20020 9044 20526
rect 8988 19954 9044 19964
rect 8652 19058 8708 19068
rect 8764 19628 8932 19684
rect 8652 18676 8708 18686
rect 8540 18674 8708 18676
rect 8540 18622 8654 18674
rect 8706 18622 8708 18674
rect 8540 18620 8708 18622
rect 8428 18398 8430 18450
rect 8482 18398 8484 18450
rect 8428 18386 8484 18398
rect 7644 17890 7700 17902
rect 7644 17838 7646 17890
rect 7698 17838 7700 17890
rect 7644 17778 7700 17838
rect 7644 17726 7646 17778
rect 7698 17726 7700 17778
rect 7644 17714 7700 17726
rect 8316 17668 8372 17678
rect 8204 17666 8372 17668
rect 8204 17614 8318 17666
rect 8370 17614 8372 17666
rect 8204 17612 8372 17614
rect 7868 17556 7924 17566
rect 7868 17462 7924 17500
rect 8092 17556 8148 17566
rect 8092 17462 8148 17500
rect 8204 17220 8260 17612
rect 8316 17602 8372 17612
rect 8652 17666 8708 18620
rect 8652 17614 8654 17666
rect 8706 17614 8708 17666
rect 8652 17602 8708 17614
rect 8764 17556 8820 19628
rect 8988 19124 9044 19134
rect 8876 19122 9044 19124
rect 8876 19070 8990 19122
rect 9042 19070 9044 19122
rect 8876 19068 9044 19070
rect 8876 18452 8932 19068
rect 8988 19058 9044 19068
rect 9100 19010 9156 19022
rect 9100 18958 9102 19010
rect 9154 18958 9156 19010
rect 8876 18386 8932 18396
rect 8988 18450 9044 18462
rect 8988 18398 8990 18450
rect 9042 18398 9044 18450
rect 8988 17892 9044 18398
rect 9100 18452 9156 18958
rect 9212 19012 9268 23772
rect 9324 22820 9380 22830
rect 9324 20132 9380 22764
rect 9548 21698 9604 26852
rect 9660 26292 9716 27804
rect 10332 27746 10388 27758
rect 10332 27694 10334 27746
rect 10386 27694 10388 27746
rect 9996 27076 10052 27086
rect 10220 27076 10276 27086
rect 9996 27074 10220 27076
rect 9996 27022 9998 27074
rect 10050 27022 10220 27074
rect 9996 27020 10220 27022
rect 9996 27010 10052 27020
rect 10220 27010 10276 27020
rect 10332 26962 10388 27694
rect 10780 27076 10836 27086
rect 10780 26982 10836 27020
rect 10332 26910 10334 26962
rect 10386 26910 10388 26962
rect 10332 26898 10388 26910
rect 10108 26628 10164 26638
rect 10108 26514 10164 26572
rect 10892 26516 10948 28476
rect 11564 28642 11620 30492
rect 11564 28590 11566 28642
rect 11618 28590 11620 28642
rect 10108 26462 10110 26514
rect 10162 26462 10164 26514
rect 10108 26450 10164 26462
rect 10668 26460 10948 26516
rect 11116 27188 11172 27198
rect 11116 26516 11172 27132
rect 11564 27074 11620 28590
rect 11788 30322 11844 30334
rect 11788 30270 11790 30322
rect 11842 30270 11844 30322
rect 11564 27022 11566 27074
rect 11618 27022 11620 27074
rect 11564 27010 11620 27022
rect 11676 28532 11732 28542
rect 11788 28532 11844 30270
rect 12236 30210 12292 32508
rect 12460 32470 12516 32508
rect 13580 32564 13636 33294
rect 13580 32498 13636 32508
rect 13132 32450 13188 32462
rect 13132 32398 13134 32450
rect 13186 32398 13188 32450
rect 13132 31892 13188 32398
rect 13132 31826 13188 31836
rect 13916 31892 13972 31902
rect 13916 31798 13972 31836
rect 13804 31780 13860 31790
rect 13468 31668 13524 31678
rect 13244 31220 13300 31230
rect 13244 31126 13300 31164
rect 13468 31106 13524 31612
rect 13468 31054 13470 31106
rect 13522 31054 13524 31106
rect 13468 31042 13524 31054
rect 13804 31106 13860 31724
rect 14140 31778 14196 33740
rect 14252 33906 14532 33908
rect 14252 33854 14478 33906
rect 14530 33854 14532 33906
rect 14252 33852 14532 33854
rect 14252 33458 14308 33852
rect 14476 33842 14532 33852
rect 14252 33406 14254 33458
rect 14306 33406 14308 33458
rect 14252 33394 14308 33406
rect 14140 31726 14142 31778
rect 14194 31726 14196 31778
rect 14140 31714 14196 31726
rect 14476 31890 14532 31902
rect 14476 31838 14478 31890
rect 14530 31838 14532 31890
rect 13804 31054 13806 31106
rect 13858 31054 13860 31106
rect 13804 31042 13860 31054
rect 14140 31220 14196 31230
rect 14140 30994 14196 31164
rect 14140 30942 14142 30994
rect 14194 30942 14196 30994
rect 14140 30930 14196 30942
rect 13132 30772 13188 30782
rect 12236 30158 12238 30210
rect 12290 30158 12292 30210
rect 12236 29428 12292 30158
rect 12908 30770 13188 30772
rect 12908 30718 13134 30770
rect 13186 30718 13188 30770
rect 12908 30716 13188 30718
rect 12908 29538 12964 30716
rect 13132 30706 13188 30716
rect 14140 30772 14196 30782
rect 14140 30770 14308 30772
rect 14140 30718 14142 30770
rect 14194 30718 14308 30770
rect 14140 30716 14308 30718
rect 14140 30706 14196 30716
rect 12908 29486 12910 29538
rect 12962 29486 12964 29538
rect 12908 29474 12964 29486
rect 12236 29334 12292 29372
rect 13468 29428 13524 29438
rect 11676 28530 11844 28532
rect 11676 28478 11678 28530
rect 11730 28478 11844 28530
rect 11676 28476 11844 28478
rect 12908 28644 12964 28654
rect 11676 26908 11732 28476
rect 12908 28082 12964 28588
rect 13468 28644 13524 29372
rect 14252 28754 14308 30716
rect 14252 28702 14254 28754
rect 14306 28702 14308 28754
rect 14252 28690 14308 28702
rect 13468 28550 13524 28588
rect 13804 28644 13860 28654
rect 12908 28030 12910 28082
rect 12962 28030 12964 28082
rect 12460 27746 12516 27758
rect 12460 27694 12462 27746
rect 12514 27694 12516 27746
rect 11900 26962 11956 26974
rect 11900 26910 11902 26962
rect 11954 26910 11956 26962
rect 11900 26908 11956 26910
rect 12460 26908 12516 27694
rect 11676 26852 11844 26908
rect 11900 26852 12516 26908
rect 9660 24722 9716 26236
rect 10556 26402 10612 26414
rect 10556 26350 10558 26402
rect 10610 26350 10612 26402
rect 9884 25620 9940 25630
rect 9884 25526 9940 25564
rect 10332 25284 10388 25294
rect 10332 25190 10388 25228
rect 10444 24836 10500 24846
rect 10556 24836 10612 26350
rect 10668 25730 10724 26460
rect 11116 26450 11172 26460
rect 10892 26292 10948 26302
rect 10892 26290 11172 26292
rect 10892 26238 10894 26290
rect 10946 26238 11172 26290
rect 10892 26236 11172 26238
rect 10892 26226 10948 26236
rect 10668 25678 10670 25730
rect 10722 25678 10724 25730
rect 10668 25396 10724 25678
rect 10668 25330 10724 25340
rect 10444 24834 10612 24836
rect 10444 24782 10446 24834
rect 10498 24782 10612 24834
rect 10444 24780 10612 24782
rect 10444 24770 10500 24780
rect 9660 24670 9662 24722
rect 9714 24670 9716 24722
rect 9660 24658 9716 24670
rect 11116 24164 11172 26236
rect 11452 25732 11508 25742
rect 11228 25620 11284 25630
rect 11228 25394 11284 25564
rect 11228 25342 11230 25394
rect 11282 25342 11284 25394
rect 11228 25330 11284 25342
rect 11452 25506 11508 25676
rect 11452 25454 11454 25506
rect 11506 25454 11508 25506
rect 11452 25284 11508 25454
rect 11452 25218 11508 25228
rect 11564 25396 11620 25406
rect 11228 24164 11284 24174
rect 11116 24162 11284 24164
rect 11116 24110 11230 24162
rect 11282 24110 11284 24162
rect 11116 24108 11284 24110
rect 11228 24098 11284 24108
rect 11564 24162 11620 25340
rect 11564 24110 11566 24162
rect 11618 24110 11620 24162
rect 11564 24098 11620 24110
rect 9660 23156 9716 23166
rect 9660 22370 9716 23100
rect 9660 22318 9662 22370
rect 9714 22318 9716 22370
rect 9660 22306 9716 22318
rect 10444 22260 10500 22270
rect 10444 22258 10948 22260
rect 10444 22206 10446 22258
rect 10498 22206 10948 22258
rect 10444 22204 10948 22206
rect 10444 22194 10500 22204
rect 9548 21646 9550 21698
rect 9602 21646 9604 21698
rect 9548 21634 9604 21646
rect 9884 21812 9940 21822
rect 9772 21588 9828 21598
rect 9884 21588 9940 21756
rect 10892 21810 10948 22204
rect 11788 21812 11844 26852
rect 11900 25396 11956 25406
rect 11900 25302 11956 25340
rect 10892 21758 10894 21810
rect 10946 21758 10948 21810
rect 10892 21746 10948 21758
rect 11676 21756 11844 21812
rect 10108 21700 10164 21710
rect 9996 21588 10052 21598
rect 9884 21586 10052 21588
rect 9884 21534 9998 21586
rect 10050 21534 10052 21586
rect 9884 21532 10052 21534
rect 9772 21494 9828 21532
rect 9996 21522 10052 21532
rect 10108 21586 10164 21644
rect 11228 21700 11284 21710
rect 11228 21606 11284 21644
rect 10108 21534 10110 21586
rect 10162 21534 10164 21586
rect 10108 21522 10164 21534
rect 11676 21588 11732 21756
rect 11900 21700 11956 21710
rect 11900 21606 11956 21644
rect 11676 21532 11844 21588
rect 9660 21476 9716 21486
rect 9660 21382 9716 21420
rect 11564 21364 11620 21374
rect 11228 20916 11284 20926
rect 11564 20916 11620 21308
rect 11788 21026 11844 21532
rect 11788 20974 11790 21026
rect 11842 20974 11844 21026
rect 11788 20962 11844 20974
rect 11228 20914 11620 20916
rect 11228 20862 11230 20914
rect 11282 20862 11620 20914
rect 11228 20860 11620 20862
rect 11228 20850 11284 20860
rect 11564 20690 11620 20860
rect 11564 20638 11566 20690
rect 11618 20638 11620 20690
rect 11564 20626 11620 20638
rect 11676 20578 11732 20590
rect 11676 20526 11678 20578
rect 11730 20526 11732 20578
rect 9772 20132 9828 20142
rect 9324 20130 9828 20132
rect 9324 20078 9774 20130
rect 9826 20078 9828 20130
rect 9324 20076 9828 20078
rect 9324 19234 9380 20076
rect 9772 20066 9828 20076
rect 9548 19908 9604 19918
rect 9548 19814 9604 19852
rect 9884 19796 9940 19806
rect 11564 19796 11620 19806
rect 9884 19794 10388 19796
rect 9884 19742 9886 19794
rect 9938 19742 10388 19794
rect 9884 19740 10388 19742
rect 9884 19730 9940 19740
rect 10332 19458 10388 19740
rect 11564 19702 11620 19740
rect 10332 19406 10334 19458
rect 10386 19406 10388 19458
rect 10332 19394 10388 19406
rect 10668 19292 11508 19348
rect 9324 19182 9326 19234
rect 9378 19182 9380 19234
rect 9324 19170 9380 19182
rect 10220 19234 10276 19246
rect 10668 19236 10724 19292
rect 10220 19182 10222 19234
rect 10274 19182 10276 19234
rect 9884 19122 9940 19134
rect 9884 19070 9886 19122
rect 9938 19070 9940 19122
rect 9884 19012 9940 19070
rect 9212 18956 9940 19012
rect 10108 19012 10164 19022
rect 10108 18918 10164 18956
rect 9548 18676 9604 18686
rect 9100 18386 9156 18396
rect 9436 18564 9492 18574
rect 8988 17836 9156 17892
rect 8988 17556 9044 17566
rect 8764 17500 8988 17556
rect 9100 17556 9156 17836
rect 9212 17556 9268 17566
rect 9100 17500 9212 17556
rect 8988 17462 9044 17500
rect 9212 17490 9268 17500
rect 8316 17444 8372 17454
rect 8316 17350 8372 17388
rect 9324 17442 9380 17454
rect 9324 17390 9326 17442
rect 9378 17390 9380 17442
rect 9212 17332 9268 17342
rect 7756 17164 8260 17220
rect 9100 17276 9212 17332
rect 7644 17108 7700 17118
rect 7532 17106 7700 17108
rect 7532 17054 7646 17106
rect 7698 17054 7700 17106
rect 7532 17052 7700 17054
rect 7644 17042 7700 17052
rect 7308 16818 7364 16828
rect 7644 16884 7700 16894
rect 7420 16772 7476 16782
rect 7420 16678 7476 16716
rect 7644 16436 7700 16828
rect 7756 16770 7812 17164
rect 8428 17108 8484 17118
rect 8988 17108 9044 17118
rect 9100 17108 9156 17276
rect 9212 17266 9268 17276
rect 8428 17106 9156 17108
rect 8428 17054 8430 17106
rect 8482 17054 8990 17106
rect 9042 17054 9156 17106
rect 8428 17052 9156 17054
rect 8428 17042 8484 17052
rect 8988 17042 9044 17052
rect 7868 16996 7924 17006
rect 8092 16996 8148 17006
rect 7924 16994 8148 16996
rect 7924 16942 8094 16994
rect 8146 16942 8148 16994
rect 7924 16940 8148 16942
rect 7868 16930 7924 16940
rect 8092 16930 8148 16940
rect 7756 16718 7758 16770
rect 7810 16718 7812 16770
rect 7756 16706 7812 16718
rect 9324 16548 9380 17390
rect 9324 16482 9380 16492
rect 7644 16380 7812 16436
rect 7196 16268 7700 16324
rect 7420 15988 7476 15998
rect 7420 15148 7476 15932
rect 7644 15986 7700 16268
rect 7644 15934 7646 15986
rect 7698 15934 7700 15986
rect 7644 15540 7700 15934
rect 7756 15988 7812 16380
rect 7756 15894 7812 15932
rect 8204 16098 8260 16110
rect 8204 16046 8206 16098
rect 8258 16046 8260 16098
rect 7644 15474 7700 15484
rect 7308 15092 7476 15148
rect 8204 15202 8260 16046
rect 8988 15986 9044 15998
rect 8988 15934 8990 15986
rect 9042 15934 9044 15986
rect 8204 15150 8206 15202
rect 8258 15150 8260 15202
rect 7084 14700 7252 14756
rect 7084 14532 7140 14542
rect 7084 14438 7140 14476
rect 7196 13858 7252 14700
rect 7196 13806 7198 13858
rect 7250 13806 7252 13858
rect 6860 12852 6916 12862
rect 6748 12850 6916 12852
rect 6748 12798 6862 12850
rect 6914 12798 6916 12850
rect 6748 12796 6916 12798
rect 4060 12338 4116 12348
rect 4620 12628 4676 12638
rect 2492 12238 2494 12290
rect 2546 12238 2548 12290
rect 2492 12226 2548 12238
rect 1820 12126 1822 12178
rect 1874 12126 1876 12178
rect 1820 11508 1876 12126
rect 4620 12066 4676 12572
rect 5404 12628 5460 12638
rect 5068 12404 5124 12414
rect 5068 12310 5124 12348
rect 5404 12178 5460 12572
rect 6076 12292 6132 12302
rect 6076 12198 6132 12236
rect 5404 12126 5406 12178
rect 5458 12126 5460 12178
rect 5404 12114 5460 12126
rect 6188 12178 6244 12796
rect 6412 12786 6468 12796
rect 6188 12126 6190 12178
rect 6242 12126 6244 12178
rect 6188 12114 6244 12126
rect 4620 12014 4622 12066
rect 4674 12014 4676 12066
rect 4620 12002 4676 12014
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 6860 11732 6916 12796
rect 7196 12292 7252 13806
rect 7308 13746 7364 15092
rect 8204 14532 8260 15150
rect 7756 14420 7812 14430
rect 7756 14418 8036 14420
rect 7756 14366 7758 14418
rect 7810 14366 8036 14418
rect 7756 14364 8036 14366
rect 7756 14354 7812 14364
rect 7980 13970 8036 14364
rect 7980 13918 7982 13970
rect 8034 13918 8036 13970
rect 7980 13906 8036 13918
rect 7308 13694 7310 13746
rect 7362 13694 7364 13746
rect 7308 13682 7364 13694
rect 8204 13636 8260 14476
rect 8316 15876 8372 15886
rect 8316 13858 8372 15820
rect 8316 13806 8318 13858
rect 8370 13806 8372 13858
rect 8316 13794 8372 13806
rect 8540 15316 8596 15326
rect 8204 13570 8260 13580
rect 8540 13412 8596 15260
rect 8988 14420 9044 15934
rect 8988 14354 9044 14364
rect 9100 13972 9156 13982
rect 9100 13878 9156 13916
rect 7196 12226 7252 12236
rect 8204 13300 8260 13310
rect 7308 11788 7588 11844
rect 7308 11732 7364 11788
rect 6860 11676 7364 11732
rect 7420 11620 7476 11630
rect 1820 11442 1876 11452
rect 4844 11508 4900 11518
rect 4844 11414 4900 11452
rect 5628 11508 5684 11518
rect 5628 11394 5684 11452
rect 5628 11342 5630 11394
rect 5682 11342 5684 11394
rect 5628 11330 5684 11342
rect 6076 11508 6132 11518
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 6076 9042 6132 11452
rect 6412 11282 6468 11294
rect 6412 11230 6414 11282
rect 6466 11230 6468 11282
rect 6300 10836 6356 10846
rect 6412 10836 6468 11230
rect 6300 10834 6468 10836
rect 6300 10782 6302 10834
rect 6354 10782 6468 10834
rect 6300 10780 6468 10782
rect 6300 10770 6356 10780
rect 6636 10612 6692 10622
rect 7084 10612 7140 10622
rect 6636 10610 7140 10612
rect 6636 10558 6638 10610
rect 6690 10558 7086 10610
rect 7138 10558 7140 10610
rect 6636 10556 7140 10558
rect 6636 10546 6692 10556
rect 7084 10546 7140 10556
rect 7420 10610 7476 11564
rect 7532 10724 7588 11788
rect 7980 10724 8036 10734
rect 7532 10722 8036 10724
rect 7532 10670 7982 10722
rect 8034 10670 8036 10722
rect 7532 10668 8036 10670
rect 7980 10658 8036 10668
rect 8204 10612 8260 13244
rect 8540 13074 8596 13356
rect 8540 13022 8542 13074
rect 8594 13022 8596 13074
rect 8540 13010 8596 13022
rect 8876 13636 8932 13646
rect 8876 12962 8932 13580
rect 8876 12910 8878 12962
rect 8930 12910 8932 12962
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 7420 10546 7476 10558
rect 8092 10610 8260 10612
rect 8092 10558 8206 10610
rect 8258 10558 8260 10610
rect 8092 10556 8260 10558
rect 6636 9826 6692 9838
rect 6636 9774 6638 9826
rect 6690 9774 6692 9826
rect 6636 9716 6692 9774
rect 7644 9826 7700 9838
rect 7644 9774 7646 9826
rect 7698 9774 7700 9826
rect 6636 9650 6692 9660
rect 7308 9716 7364 9726
rect 7308 9622 7364 9660
rect 6860 9602 6916 9614
rect 6860 9550 6862 9602
rect 6914 9550 6916 9602
rect 6860 9154 6916 9550
rect 6860 9102 6862 9154
rect 6914 9102 6916 9154
rect 6860 9090 6916 9102
rect 6076 8990 6078 9042
rect 6130 8990 6132 9042
rect 6076 8978 6132 8990
rect 7644 8932 7700 9774
rect 8092 9826 8148 10556
rect 8204 10546 8260 10556
rect 8316 12292 8372 12302
rect 8092 9774 8094 9826
rect 8146 9774 8148 9826
rect 8092 9762 8148 9774
rect 8316 9714 8372 12236
rect 8540 11620 8596 11630
rect 8540 11506 8596 11564
rect 8540 11454 8542 11506
rect 8594 11454 8596 11506
rect 8540 11284 8596 11454
rect 8876 11508 8932 12910
rect 9436 12628 9492 18508
rect 9548 18562 9604 18620
rect 9548 18510 9550 18562
rect 9602 18510 9604 18562
rect 9548 18498 9604 18510
rect 9884 18450 9940 18462
rect 9884 18398 9886 18450
rect 9938 18398 9940 18450
rect 9660 18338 9716 18350
rect 9660 18286 9662 18338
rect 9714 18286 9716 18338
rect 9660 18228 9716 18286
rect 9660 18162 9716 18172
rect 9884 18228 9940 18398
rect 9996 18452 10052 18462
rect 9996 18358 10052 18396
rect 10220 18452 10276 19182
rect 10220 18228 10276 18396
rect 9884 18172 10276 18228
rect 10332 19234 10724 19236
rect 10332 19182 10670 19234
rect 10722 19182 10724 19234
rect 10332 19180 10724 19182
rect 11452 19236 11508 19292
rect 11564 19236 11620 19246
rect 11452 19234 11620 19236
rect 11452 19182 11566 19234
rect 11618 19182 11620 19234
rect 11452 19180 11620 19182
rect 10332 18450 10388 19180
rect 10668 19170 10724 19180
rect 11116 19122 11172 19134
rect 11116 19070 11118 19122
rect 11170 19070 11172 19122
rect 11116 18564 11172 19070
rect 11340 19122 11396 19134
rect 11340 19070 11342 19122
rect 11394 19070 11396 19122
rect 11228 18564 11284 18574
rect 11116 18562 11284 18564
rect 11116 18510 11230 18562
rect 11282 18510 11284 18562
rect 11116 18508 11284 18510
rect 10332 18398 10334 18450
rect 10386 18398 10388 18450
rect 9548 17780 9604 17790
rect 9548 17106 9604 17724
rect 9548 17054 9550 17106
rect 9602 17054 9604 17106
rect 9548 17042 9604 17054
rect 9772 17666 9828 17678
rect 9772 17614 9774 17666
rect 9826 17614 9828 17666
rect 9772 16548 9828 17614
rect 9884 17556 9940 18172
rect 9996 17556 10052 17566
rect 9884 17554 10052 17556
rect 9884 17502 9998 17554
rect 10050 17502 10052 17554
rect 9884 17500 10052 17502
rect 9996 17490 10052 17500
rect 10332 17554 10388 18398
rect 11004 18450 11060 18462
rect 11004 18398 11006 18450
rect 11058 18398 11060 18450
rect 10332 17502 10334 17554
rect 10386 17502 10388 17554
rect 10332 17490 10388 17502
rect 10444 18116 10500 18126
rect 9884 17108 9940 17118
rect 10332 17108 10388 17118
rect 10444 17108 10500 18060
rect 10668 17556 10724 17566
rect 10668 17462 10724 17500
rect 9884 17106 10500 17108
rect 9884 17054 9886 17106
rect 9938 17054 10334 17106
rect 10386 17054 10500 17106
rect 9884 17052 10500 17054
rect 9884 17042 9940 17052
rect 10332 17042 10388 17052
rect 9772 16482 9828 16492
rect 10332 16884 10388 16894
rect 10332 15426 10388 16828
rect 10892 16770 10948 16782
rect 10892 16718 10894 16770
rect 10946 16718 10948 16770
rect 10332 15374 10334 15426
rect 10386 15374 10388 15426
rect 10332 15316 10388 15374
rect 10332 15250 10388 15260
rect 10444 15988 10500 15998
rect 10444 15314 10500 15932
rect 10892 15988 10948 16718
rect 10892 15922 10948 15932
rect 10444 15262 10446 15314
rect 10498 15262 10500 15314
rect 10444 15250 10500 15262
rect 9772 15202 9828 15214
rect 9772 15150 9774 15202
rect 9826 15150 9828 15202
rect 9772 13300 9828 15150
rect 11004 14754 11060 18398
rect 11116 18452 11172 18508
rect 11228 18498 11284 18508
rect 11116 18386 11172 18396
rect 11116 18004 11172 18014
rect 11116 17442 11172 17948
rect 11116 17390 11118 17442
rect 11170 17390 11172 17442
rect 11116 16884 11172 17390
rect 11340 17106 11396 19070
rect 11452 18674 11508 18686
rect 11452 18622 11454 18674
rect 11506 18622 11508 18674
rect 11452 18452 11508 18622
rect 11452 18386 11508 18396
rect 11564 18450 11620 19180
rect 11564 18398 11566 18450
rect 11618 18398 11620 18450
rect 11564 18386 11620 18398
rect 11564 18228 11620 18238
rect 11676 18228 11732 20526
rect 12012 20132 12068 26852
rect 12348 26292 12404 26302
rect 12908 26292 12964 28030
rect 13804 27858 13860 28588
rect 14476 27970 14532 31838
rect 14588 31666 14644 34972
rect 15036 35026 15372 35028
rect 15036 34974 15038 35026
rect 15090 34974 15372 35026
rect 15036 34972 15372 34974
rect 15036 34962 15092 34972
rect 15372 34914 15428 34972
rect 15372 34862 15374 34914
rect 15426 34862 15428 34914
rect 15372 34850 15428 34862
rect 15484 34356 15540 36428
rect 15820 35924 15876 36652
rect 16156 36708 16212 36718
rect 16156 36594 16212 36652
rect 16156 36542 16158 36594
rect 16210 36542 16212 36594
rect 16156 36530 16212 36542
rect 16492 36596 16548 38556
rect 16604 38276 16660 39340
rect 16604 38210 16660 38220
rect 16716 36596 16772 39564
rect 17052 39508 17108 39518
rect 17052 39414 17108 39452
rect 17164 38612 17220 41692
rect 17500 41300 17556 42588
rect 17388 41244 17556 41300
rect 17724 42532 17780 42542
rect 17388 41188 17444 41244
rect 17164 38546 17220 38556
rect 17276 41186 17444 41188
rect 17276 41134 17390 41186
rect 17442 41134 17444 41186
rect 17276 41132 17444 41134
rect 17276 38388 17332 41132
rect 17388 41122 17444 41132
rect 17724 41186 17780 42476
rect 17724 41134 17726 41186
rect 17778 41134 17780 41186
rect 17612 40962 17668 40974
rect 17612 40910 17614 40962
rect 17666 40910 17668 40962
rect 17500 40402 17556 40414
rect 17500 40350 17502 40402
rect 17554 40350 17556 40402
rect 17500 39508 17556 40350
rect 17612 40292 17668 40910
rect 17612 40226 17668 40236
rect 17724 39844 17780 41134
rect 17836 42082 17892 43260
rect 17948 42868 18004 42878
rect 17948 42642 18004 42812
rect 17948 42590 17950 42642
rect 18002 42590 18004 42642
rect 17948 42578 18004 42590
rect 18060 42642 18116 43484
rect 18172 43538 18228 44380
rect 18284 44324 18340 44334
rect 18284 44230 18340 44268
rect 18172 43486 18174 43538
rect 18226 43486 18228 43538
rect 18172 43474 18228 43486
rect 18284 43876 18340 43886
rect 18396 43876 18452 45166
rect 18844 45220 18900 45838
rect 18844 45154 18900 45164
rect 18956 45836 19460 45892
rect 19516 46340 19572 46350
rect 18620 45106 18676 45118
rect 18620 45054 18622 45106
rect 18674 45054 18676 45106
rect 18620 44996 18676 45054
rect 18620 44322 18676 44940
rect 18620 44270 18622 44322
rect 18674 44270 18676 44322
rect 18620 44258 18676 44270
rect 18956 45106 19012 45836
rect 19404 45668 19460 45678
rect 19180 45666 19460 45668
rect 19180 45614 19406 45666
rect 19458 45614 19460 45666
rect 19180 45612 19460 45614
rect 18956 45054 18958 45106
rect 19010 45054 19012 45106
rect 18956 44324 19012 45054
rect 18956 44258 19012 44268
rect 19068 45108 19124 45118
rect 19068 44772 19124 45052
rect 18844 44100 18900 44110
rect 18340 43820 18452 43876
rect 18732 44044 18844 44100
rect 18060 42590 18062 42642
rect 18114 42590 18116 42642
rect 18060 42420 18116 42590
rect 18060 42354 18116 42364
rect 17836 42030 17838 42082
rect 17890 42030 17892 42082
rect 17836 40628 17892 42030
rect 17948 42084 18004 42094
rect 17948 41972 18004 42028
rect 18172 41972 18228 41982
rect 17948 41970 18116 41972
rect 17948 41918 17950 41970
rect 18002 41918 18116 41970
rect 17948 41916 18116 41918
rect 17948 41906 18004 41916
rect 18060 41636 18116 41916
rect 18172 41878 18228 41916
rect 18284 41860 18340 43820
rect 18396 43652 18452 43662
rect 18396 43538 18452 43596
rect 18396 43486 18398 43538
rect 18450 43486 18452 43538
rect 18396 43474 18452 43486
rect 18620 43316 18676 43326
rect 18620 43222 18676 43260
rect 18508 42644 18564 42654
rect 18508 42550 18564 42588
rect 18732 42642 18788 44044
rect 18844 44034 18900 44044
rect 18844 43652 18900 43662
rect 19068 43652 19124 44716
rect 18844 43650 19124 43652
rect 18844 43598 18846 43650
rect 18898 43598 19124 43650
rect 18844 43596 19124 43598
rect 18844 43586 18900 43596
rect 19180 43540 19236 45612
rect 19404 45556 19460 45612
rect 19404 45490 19460 45500
rect 19292 44884 19348 44894
rect 19292 44210 19348 44828
rect 19292 44158 19294 44210
rect 19346 44158 19348 44210
rect 19292 43988 19348 44158
rect 19292 43922 19348 43932
rect 19404 44322 19460 44334
rect 19404 44270 19406 44322
rect 19458 44270 19460 44322
rect 19404 43876 19460 44270
rect 19404 43810 19460 43820
rect 19292 43764 19348 43774
rect 19516 43708 19572 46284
rect 19628 46004 19684 46620
rect 20412 46674 20468 47404
rect 20412 46622 20414 46674
rect 20466 46622 20468 46674
rect 20412 46610 20468 46622
rect 20524 47458 20580 47470
rect 20524 47406 20526 47458
rect 20578 47406 20580 47458
rect 20188 46562 20244 46574
rect 20188 46510 20190 46562
rect 20242 46510 20244 46562
rect 20188 46452 20244 46510
rect 20524 46452 20580 47406
rect 20636 46564 20692 48862
rect 20748 48244 20804 49534
rect 20748 48178 20804 48188
rect 20972 49028 21028 52108
rect 22204 51602 22260 52892
rect 22764 52052 22820 52062
rect 22204 51550 22206 51602
rect 22258 51550 22260 51602
rect 22204 51538 22260 51550
rect 22316 51604 22372 51614
rect 22092 51268 22148 51278
rect 22092 51174 22148 51212
rect 21980 50596 22036 50606
rect 21980 50034 22036 50540
rect 22316 50484 22372 51548
rect 22540 50484 22596 50494
rect 22316 50482 22596 50484
rect 22316 50430 22542 50482
rect 22594 50430 22596 50482
rect 22316 50428 22596 50430
rect 21980 49982 21982 50034
rect 22034 49982 22036 50034
rect 21980 49970 22036 49982
rect 22204 50372 22372 50428
rect 22540 50418 22596 50428
rect 22092 49924 22148 49934
rect 21084 49810 21140 49822
rect 21084 49758 21086 49810
rect 21138 49758 21140 49810
rect 21084 49476 21140 49758
rect 21196 49588 21252 49598
rect 21196 49494 21252 49532
rect 21308 49586 21364 49598
rect 21308 49534 21310 49586
rect 21362 49534 21364 49586
rect 21084 49410 21140 49420
rect 20972 48466 21028 48972
rect 21308 49026 21364 49534
rect 21868 49588 21924 49598
rect 21868 49494 21924 49532
rect 22092 49364 22148 49868
rect 22204 49812 22260 50372
rect 22428 49812 22484 49822
rect 22204 49810 22428 49812
rect 22204 49758 22206 49810
rect 22258 49758 22428 49810
rect 22204 49756 22428 49758
rect 22204 49746 22260 49756
rect 22428 49746 22484 49756
rect 22540 49810 22596 49822
rect 22540 49758 22542 49810
rect 22594 49758 22596 49810
rect 21868 49308 22148 49364
rect 21868 49250 21924 49308
rect 21868 49198 21870 49250
rect 21922 49198 21924 49250
rect 21868 49186 21924 49198
rect 22540 49252 22596 49758
rect 22652 49252 22708 49262
rect 22540 49250 22708 49252
rect 22540 49198 22654 49250
rect 22706 49198 22708 49250
rect 22540 49196 22708 49198
rect 22652 49186 22708 49196
rect 21420 49140 21476 49150
rect 21476 49084 21588 49140
rect 21420 49074 21476 49084
rect 21308 48974 21310 49026
rect 21362 48974 21364 49026
rect 21308 48916 21364 48974
rect 21532 49026 21588 49084
rect 22764 49028 22820 51996
rect 22876 51716 22932 53678
rect 24444 53732 24500 54574
rect 24556 53954 24612 55134
rect 25116 54964 25172 54974
rect 24556 53902 24558 53954
rect 24610 53902 24612 53954
rect 24556 53890 24612 53902
rect 24668 54404 24724 54414
rect 24556 53732 24612 53742
rect 24444 53730 24612 53732
rect 24444 53678 24558 53730
rect 24610 53678 24612 53730
rect 24444 53676 24612 53678
rect 23324 53620 23380 53630
rect 23212 53618 23380 53620
rect 23212 53566 23326 53618
rect 23378 53566 23380 53618
rect 23212 53564 23380 53566
rect 22988 52834 23044 52846
rect 22988 52782 22990 52834
rect 23042 52782 23044 52834
rect 22988 52164 23044 52782
rect 22988 52098 23044 52108
rect 23100 52162 23156 52174
rect 23100 52110 23102 52162
rect 23154 52110 23156 52162
rect 23100 52052 23156 52110
rect 23100 51986 23156 51996
rect 22876 51650 22932 51660
rect 23100 51492 23156 51502
rect 23100 51398 23156 51436
rect 22876 51378 22932 51390
rect 22876 51326 22878 51378
rect 22930 51326 22932 51378
rect 22876 50484 22932 51326
rect 22876 50418 22932 50428
rect 22988 50036 23044 50046
rect 23212 50036 23268 53564
rect 23324 53554 23380 53564
rect 23548 53620 23604 53630
rect 23884 53620 23940 53630
rect 24220 53620 24276 53630
rect 23548 53526 23604 53564
rect 23772 53618 23940 53620
rect 23772 53566 23886 53618
rect 23938 53566 23940 53618
rect 23772 53564 23940 53566
rect 23772 53172 23828 53564
rect 23884 53554 23940 53564
rect 23996 53618 24276 53620
rect 23996 53566 24222 53618
rect 24274 53566 24276 53618
rect 23996 53564 24276 53566
rect 23772 53106 23828 53116
rect 23884 53172 23940 53182
rect 23996 53172 24052 53564
rect 24220 53554 24276 53564
rect 23884 53170 24052 53172
rect 23884 53118 23886 53170
rect 23938 53118 24052 53170
rect 23884 53116 24052 53118
rect 24220 53172 24276 53182
rect 23884 53106 23940 53116
rect 23548 52948 23604 52958
rect 23548 52854 23604 52892
rect 23772 52948 23828 52958
rect 23996 52948 24052 52958
rect 23772 52946 23940 52948
rect 23772 52894 23774 52946
rect 23826 52894 23940 52946
rect 23772 52892 23940 52894
rect 23772 52882 23828 52892
rect 23884 52276 23940 52892
rect 23996 52854 24052 52892
rect 24220 52948 24276 53116
rect 24556 53060 24612 53676
rect 24668 53170 24724 54348
rect 24668 53118 24670 53170
rect 24722 53118 24724 53170
rect 24668 53106 24724 53118
rect 25004 53506 25060 53518
rect 25004 53454 25006 53506
rect 25058 53454 25060 53506
rect 24556 52994 24612 53004
rect 25004 53060 25060 53454
rect 25004 52994 25060 53004
rect 24220 52946 24388 52948
rect 24220 52894 24222 52946
rect 24274 52894 24388 52946
rect 24220 52892 24388 52894
rect 24220 52882 24276 52892
rect 23884 52220 24164 52276
rect 23548 52164 23604 52174
rect 23548 51268 23604 52108
rect 23996 52052 24052 52062
rect 23772 52050 24052 52052
rect 23772 51998 23998 52050
rect 24050 51998 24052 52050
rect 23772 51996 24052 51998
rect 23660 51604 23716 51614
rect 23660 51510 23716 51548
rect 23548 51212 23716 51268
rect 23436 51154 23492 51166
rect 23436 51102 23438 51154
rect 23490 51102 23492 51154
rect 23436 50820 23492 51102
rect 23436 50754 23492 50764
rect 23548 50596 23604 50606
rect 22988 50034 23268 50036
rect 22988 49982 22990 50034
rect 23042 49982 23268 50034
rect 22988 49980 23268 49982
rect 23324 50594 23604 50596
rect 23324 50542 23550 50594
rect 23602 50542 23604 50594
rect 23324 50540 23604 50542
rect 22988 49970 23044 49980
rect 22876 49924 22932 49934
rect 22876 49810 22932 49868
rect 22876 49758 22878 49810
rect 22930 49758 22932 49810
rect 22876 49746 22932 49758
rect 23100 49812 23156 49822
rect 23100 49718 23156 49756
rect 22988 49700 23044 49710
rect 22988 49606 23044 49644
rect 21532 48974 21534 49026
rect 21586 48974 21588 49026
rect 21532 48962 21588 48974
rect 21868 48972 22820 49028
rect 22988 49252 23044 49262
rect 22988 49026 23044 49196
rect 22988 48974 22990 49026
rect 23042 48974 23044 49026
rect 21308 48850 21364 48860
rect 20972 48414 20974 48466
rect 21026 48414 21028 48466
rect 20748 47234 20804 47246
rect 20748 47182 20750 47234
rect 20802 47182 20804 47234
rect 20748 47124 20804 47182
rect 20748 47058 20804 47068
rect 20748 46900 20804 46910
rect 20748 46806 20804 46844
rect 20860 46676 20916 46686
rect 20636 46508 20804 46564
rect 20188 46396 20580 46452
rect 19852 46004 19908 46014
rect 19628 46002 19908 46004
rect 19628 45950 19854 46002
rect 19906 45950 19908 46002
rect 19628 45948 19908 45950
rect 19628 44100 19684 45948
rect 19852 45938 19908 45948
rect 20300 45780 20356 45790
rect 20300 45686 20356 45724
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20300 44996 20356 45006
rect 20300 44902 20356 44940
rect 19852 44660 19908 44670
rect 19852 44322 19908 44604
rect 19852 44270 19854 44322
rect 19906 44270 19908 44322
rect 19852 44258 19908 44270
rect 20076 44324 20132 44334
rect 19740 44100 19796 44110
rect 19628 44044 19740 44100
rect 20076 44100 20132 44268
rect 20188 44100 20244 44110
rect 20076 44098 20244 44100
rect 20076 44046 20190 44098
rect 20242 44046 20244 44098
rect 20076 44044 20244 44046
rect 19740 44034 19796 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19292 43670 19348 43708
rect 19404 43652 19572 43708
rect 19964 43652 20020 43662
rect 19404 43540 19460 43652
rect 19180 43484 19348 43540
rect 19180 43316 19236 43326
rect 18956 43314 19236 43316
rect 18956 43262 19182 43314
rect 19234 43262 19236 43314
rect 18956 43260 19236 43262
rect 18844 42980 18900 42990
rect 18956 42980 19012 43260
rect 19180 43250 19236 43260
rect 18844 42978 19012 42980
rect 18844 42926 18846 42978
rect 18898 42926 19012 42978
rect 18844 42924 19012 42926
rect 18844 42914 18900 42924
rect 18732 42590 18734 42642
rect 18786 42590 18788 42642
rect 18732 42578 18788 42590
rect 19180 42420 19236 42430
rect 18844 42308 18900 42318
rect 18844 42196 18900 42252
rect 18620 42140 18900 42196
rect 18620 42138 18676 42140
rect 18508 42084 18564 42094
rect 18620 42086 18622 42138
rect 18674 42086 18676 42138
rect 18620 42074 18676 42086
rect 18508 41972 18564 42028
rect 18956 41972 19012 41982
rect 18508 41916 18788 41972
rect 18284 41804 18564 41860
rect 18508 41748 18564 41804
rect 18620 41748 18676 41758
rect 18508 41746 18676 41748
rect 18508 41694 18622 41746
rect 18674 41694 18676 41746
rect 18508 41692 18676 41694
rect 18060 41580 18340 41636
rect 18284 41410 18340 41580
rect 18284 41358 18286 41410
rect 18338 41358 18340 41410
rect 18284 41346 18340 41358
rect 17948 41188 18004 41198
rect 17948 41094 18004 41132
rect 18284 41186 18340 41198
rect 18284 41134 18286 41186
rect 18338 41134 18340 41186
rect 18284 40628 18340 41134
rect 18508 41188 18564 41692
rect 18620 41682 18676 41692
rect 18620 41412 18676 41422
rect 18732 41412 18788 41916
rect 18620 41410 18788 41412
rect 18620 41358 18622 41410
rect 18674 41358 18788 41410
rect 18620 41356 18788 41358
rect 18956 41748 19012 41916
rect 19068 41748 19124 41758
rect 18956 41746 19124 41748
rect 18956 41694 19070 41746
rect 19122 41694 19124 41746
rect 18956 41692 19124 41694
rect 18620 41346 18676 41356
rect 18508 41132 18676 41188
rect 17836 40572 18228 40628
rect 18060 40292 18116 40302
rect 17948 40290 18116 40292
rect 17948 40238 18062 40290
rect 18114 40238 18116 40290
rect 17948 40236 18116 40238
rect 17724 39778 17780 39788
rect 17836 40068 17892 40078
rect 17836 39618 17892 40012
rect 17836 39566 17838 39618
rect 17890 39566 17892 39618
rect 17836 39554 17892 39566
rect 17500 39442 17556 39452
rect 17724 39060 17780 39070
rect 17500 38836 17556 38846
rect 17276 38322 17332 38332
rect 17388 38610 17444 38622
rect 17388 38558 17390 38610
rect 17442 38558 17444 38610
rect 17388 38500 17444 38558
rect 17388 38164 17444 38444
rect 16492 36540 16660 36596
rect 15820 35810 15876 35868
rect 15820 35758 15822 35810
rect 15874 35758 15876 35810
rect 15820 35746 15876 35758
rect 15932 36482 15988 36494
rect 15932 36430 15934 36482
rect 15986 36430 15988 36482
rect 15932 36372 15988 36430
rect 15932 35812 15988 36316
rect 15932 35746 15988 35756
rect 16492 36372 16548 36382
rect 16044 35700 16100 35710
rect 16044 35606 16100 35644
rect 15596 35588 15652 35598
rect 15596 35586 15764 35588
rect 15596 35534 15598 35586
rect 15650 35534 15764 35586
rect 15596 35532 15764 35534
rect 15596 35522 15652 35532
rect 15596 34356 15652 34366
rect 15484 34354 15652 34356
rect 15484 34302 15598 34354
rect 15650 34302 15652 34354
rect 15484 34300 15652 34302
rect 15596 34290 15652 34300
rect 14812 33908 14868 33918
rect 14812 33814 14868 33852
rect 15708 33236 15764 35532
rect 16380 35476 16436 35486
rect 16492 35476 16548 36316
rect 16380 35474 16548 35476
rect 16380 35422 16382 35474
rect 16434 35422 16548 35474
rect 16380 35420 16548 35422
rect 16380 35410 16436 35420
rect 16044 34804 16100 34814
rect 16044 34802 16436 34804
rect 16044 34750 16046 34802
rect 16098 34750 16436 34802
rect 16044 34748 16436 34750
rect 16044 34738 16100 34748
rect 16380 34354 16436 34748
rect 16380 34302 16382 34354
rect 16434 34302 16436 34354
rect 16380 34290 16436 34302
rect 16268 34132 16324 34142
rect 16492 34132 16548 35420
rect 16604 35476 16660 36540
rect 16716 35700 16772 36540
rect 17052 38108 17444 38164
rect 16828 35812 16884 35822
rect 17052 35812 17108 38108
rect 17388 37828 17444 37838
rect 17388 37378 17444 37772
rect 17500 37490 17556 38780
rect 17724 38834 17780 39004
rect 17948 39060 18004 40236
rect 18060 40226 18116 40236
rect 17948 38994 18004 39004
rect 18060 39730 18116 39742
rect 18060 39678 18062 39730
rect 18114 39678 18116 39730
rect 17724 38782 17726 38834
rect 17778 38782 17780 38834
rect 17724 38770 17780 38782
rect 17948 38834 18004 38846
rect 17948 38782 17950 38834
rect 18002 38782 18004 38834
rect 17948 38668 18004 38782
rect 17836 38612 18004 38668
rect 17612 38164 17668 38174
rect 17612 38070 17668 38108
rect 17500 37438 17502 37490
rect 17554 37438 17556 37490
rect 17500 37426 17556 37438
rect 17388 37326 17390 37378
rect 17442 37326 17444 37378
rect 17388 37314 17444 37326
rect 17836 37380 17892 38556
rect 17836 37286 17892 37324
rect 17836 37044 17892 37054
rect 17276 36482 17332 36494
rect 17276 36430 17278 36482
rect 17330 36430 17332 36482
rect 16828 35810 17108 35812
rect 16828 35758 16830 35810
rect 16882 35758 17108 35810
rect 16828 35756 17108 35758
rect 17164 36258 17220 36270
rect 17164 36206 17166 36258
rect 17218 36206 17220 36258
rect 16828 35746 16884 35756
rect 16716 35634 16772 35644
rect 16604 35410 16660 35420
rect 16716 35474 16772 35486
rect 16716 35422 16718 35474
rect 16770 35422 16772 35474
rect 16604 34244 16660 34254
rect 16716 34244 16772 35422
rect 17164 35252 17220 36206
rect 17276 35700 17332 36430
rect 17388 35924 17444 35934
rect 17388 35830 17444 35868
rect 17724 35700 17780 35710
rect 17276 35698 17780 35700
rect 17276 35646 17726 35698
rect 17778 35646 17780 35698
rect 17276 35644 17780 35646
rect 17164 35186 17220 35196
rect 17276 35364 17332 35374
rect 16604 34242 16772 34244
rect 16604 34190 16606 34242
rect 16658 34190 16772 34242
rect 16604 34188 16772 34190
rect 16828 34244 16884 34254
rect 17276 34244 17332 35308
rect 16828 34242 17332 34244
rect 16828 34190 16830 34242
rect 16882 34190 17332 34242
rect 16828 34188 17332 34190
rect 16604 34178 16660 34188
rect 16828 34178 16884 34188
rect 16268 34130 16548 34132
rect 16268 34078 16270 34130
rect 16322 34078 16548 34130
rect 16268 34076 16548 34078
rect 16268 34066 16324 34076
rect 16380 33460 16436 33470
rect 16380 33458 16660 33460
rect 16380 33406 16382 33458
rect 16434 33406 16660 33458
rect 16380 33404 16660 33406
rect 16380 33394 16436 33404
rect 15820 33236 15876 33246
rect 15708 33180 15820 33236
rect 15708 32564 15764 33180
rect 15820 33170 15876 33180
rect 16380 33236 16436 33246
rect 16380 32786 16436 33180
rect 16380 32734 16382 32786
rect 16434 32734 16436 32786
rect 16380 32722 16436 32734
rect 15708 32498 15764 32508
rect 15260 32450 15316 32462
rect 15260 32398 15262 32450
rect 15314 32398 15316 32450
rect 15260 32340 15316 32398
rect 15820 32450 15876 32462
rect 15820 32398 15822 32450
rect 15874 32398 15876 32450
rect 15820 32340 15876 32398
rect 15260 32284 15876 32340
rect 15932 32338 15988 32350
rect 15932 32286 15934 32338
rect 15986 32286 15988 32338
rect 14812 31892 14868 31902
rect 14812 31798 14868 31836
rect 15596 31892 15652 31902
rect 15596 31798 15652 31836
rect 15708 31778 15764 32284
rect 15708 31726 15710 31778
rect 15762 31726 15764 31778
rect 15708 31714 15764 31726
rect 15932 31780 15988 32286
rect 16604 32004 16660 33404
rect 17276 33458 17332 34188
rect 17724 34132 17780 35644
rect 17836 34132 17892 36988
rect 18060 36370 18116 39678
rect 18172 38948 18228 40572
rect 18284 40562 18340 40572
rect 18508 40292 18564 40302
rect 18508 40198 18564 40236
rect 18284 40180 18340 40190
rect 18284 40086 18340 40124
rect 18284 39844 18340 39854
rect 18284 39506 18340 39788
rect 18620 39620 18676 41132
rect 18732 40628 18788 40638
rect 18732 40402 18788 40572
rect 18732 40350 18734 40402
rect 18786 40350 18788 40402
rect 18732 40338 18788 40350
rect 18620 39554 18676 39564
rect 18284 39454 18286 39506
rect 18338 39454 18340 39506
rect 18284 39442 18340 39454
rect 18956 39284 19012 41692
rect 19068 41682 19124 41692
rect 19180 41074 19236 42364
rect 19292 42308 19348 43484
rect 19404 42754 19460 43484
rect 19404 42702 19406 42754
rect 19458 42702 19460 42754
rect 19404 42532 19460 42702
rect 19516 43538 19572 43550
rect 19516 43486 19518 43538
rect 19570 43486 19572 43538
rect 19516 42756 19572 43486
rect 19852 42756 19908 42766
rect 19516 42700 19852 42756
rect 19852 42662 19908 42700
rect 19404 42466 19460 42476
rect 19964 42530 20020 43596
rect 19964 42478 19966 42530
rect 20018 42478 20020 42530
rect 19964 42466 20020 42478
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19292 42242 19348 42252
rect 19292 42084 19348 42094
rect 19740 42084 19796 42094
rect 19964 42084 20020 42094
rect 19292 41990 19348 42028
rect 19404 42082 19796 42084
rect 19404 42030 19742 42082
rect 19794 42030 19796 42082
rect 19404 42028 19796 42030
rect 19404 41858 19460 42028
rect 19740 42018 19796 42028
rect 19852 42082 20020 42084
rect 19852 42030 19966 42082
rect 20018 42030 20020 42082
rect 19852 42028 20020 42030
rect 19404 41806 19406 41858
rect 19458 41806 19460 41858
rect 19404 41794 19460 41806
rect 19628 41300 19684 41310
rect 19404 41298 19684 41300
rect 19404 41246 19630 41298
rect 19682 41246 19684 41298
rect 19404 41244 19684 41246
rect 19180 41022 19182 41074
rect 19234 41022 19236 41074
rect 19180 41010 19236 41022
rect 19292 41074 19348 41086
rect 19292 41022 19294 41074
rect 19346 41022 19348 41074
rect 19068 40964 19124 40974
rect 19068 40870 19124 40908
rect 19292 40404 19348 41022
rect 19404 40628 19460 41244
rect 19628 41234 19684 41244
rect 19740 41186 19796 41198
rect 19740 41134 19742 41186
rect 19794 41134 19796 41186
rect 19740 41076 19796 41134
rect 19404 40562 19460 40572
rect 19516 41020 19796 41076
rect 19516 40516 19572 41020
rect 19852 40964 19908 42028
rect 19964 42018 20020 42028
rect 20188 42084 20244 44044
rect 19964 41860 20020 41898
rect 19964 41794 20020 41804
rect 19964 41636 20020 41646
rect 19964 41410 20020 41580
rect 19964 41358 19966 41410
rect 20018 41358 20020 41410
rect 19964 41346 20020 41358
rect 20188 41412 20244 42028
rect 20300 41972 20356 41982
rect 20300 41878 20356 41916
rect 20300 41412 20356 41422
rect 20188 41410 20356 41412
rect 20188 41358 20302 41410
rect 20354 41358 20356 41410
rect 20188 41356 20356 41358
rect 20300 41346 20356 41356
rect 19516 40450 19572 40460
rect 19628 40908 19908 40964
rect 20188 41186 20244 41198
rect 20188 41134 20190 41186
rect 20242 41134 20244 41186
rect 18732 39228 19012 39284
rect 19068 40348 19348 40404
rect 19628 40402 19684 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19628 40350 19630 40402
rect 19682 40350 19684 40402
rect 18620 39172 18676 39182
rect 18396 38948 18452 38958
rect 18172 38946 18452 38948
rect 18172 38894 18398 38946
rect 18450 38894 18452 38946
rect 18172 38892 18452 38894
rect 18396 38882 18452 38892
rect 18284 38724 18340 38762
rect 18284 38658 18340 38668
rect 18508 38164 18564 38174
rect 18060 36318 18062 36370
rect 18114 36318 18116 36370
rect 18060 36306 18116 36318
rect 18172 38050 18228 38062
rect 18172 37998 18174 38050
rect 18226 37998 18228 38050
rect 18172 37490 18228 37998
rect 18172 37438 18174 37490
rect 18226 37438 18228 37490
rect 17948 35924 18004 35934
rect 17948 35698 18004 35868
rect 17948 35646 17950 35698
rect 18002 35646 18004 35698
rect 17948 35634 18004 35646
rect 18172 35026 18228 37438
rect 18396 37156 18452 37166
rect 18396 35922 18452 37100
rect 18508 36260 18564 38108
rect 18620 37266 18676 39116
rect 18732 37938 18788 39228
rect 18844 39058 18900 39070
rect 18844 39006 18846 39058
rect 18898 39006 18900 39058
rect 18844 38668 18900 39006
rect 19068 38668 19124 40348
rect 19628 40292 19684 40350
rect 19292 40236 19684 40292
rect 19740 40628 19796 40638
rect 19180 40180 19236 40190
rect 19180 40086 19236 40124
rect 19292 40068 19348 40236
rect 19740 40180 19796 40572
rect 19292 40002 19348 40012
rect 19404 40124 19796 40180
rect 19964 40402 20020 40414
rect 19964 40350 19966 40402
rect 20018 40350 20020 40402
rect 19292 39172 19348 39182
rect 19404 39172 19460 40124
rect 19348 39116 19460 39172
rect 19628 39618 19684 39630
rect 19628 39566 19630 39618
rect 19682 39566 19684 39618
rect 19292 39106 19348 39116
rect 18844 38612 19124 38668
rect 18732 37886 18734 37938
rect 18786 37886 18788 37938
rect 18732 37716 18788 37886
rect 19068 37828 19124 38612
rect 19628 37828 19684 39566
rect 19964 39508 20020 40350
rect 20188 40292 20244 41134
rect 20412 40404 20468 46396
rect 20636 46004 20692 46014
rect 20636 45892 20692 45948
rect 20524 45890 20692 45892
rect 20524 45838 20638 45890
rect 20690 45838 20692 45890
rect 20524 45836 20692 45838
rect 20524 44324 20580 45836
rect 20636 45826 20692 45836
rect 20524 44258 20580 44268
rect 20636 45106 20692 45118
rect 20636 45054 20638 45106
rect 20690 45054 20692 45106
rect 20636 44100 20692 45054
rect 20636 44034 20692 44044
rect 20636 43650 20692 43662
rect 20636 43598 20638 43650
rect 20690 43598 20692 43650
rect 20636 43540 20692 43598
rect 20636 43474 20692 43484
rect 20748 43316 20804 46508
rect 20860 43428 20916 46620
rect 20860 43362 20916 43372
rect 20636 43260 20804 43316
rect 20524 43204 20580 43214
rect 20524 42866 20580 43148
rect 20524 42814 20526 42866
rect 20578 42814 20580 42866
rect 20524 42802 20580 42814
rect 20636 42084 20692 43260
rect 20524 42028 20692 42084
rect 20524 41860 20580 42028
rect 20748 41972 20804 41982
rect 20524 41794 20580 41804
rect 20636 41970 20804 41972
rect 20636 41918 20750 41970
rect 20802 41918 20804 41970
rect 20636 41916 20804 41918
rect 20412 40402 20580 40404
rect 20412 40350 20414 40402
rect 20466 40350 20580 40402
rect 20412 40348 20580 40350
rect 20412 40338 20468 40348
rect 20188 40226 20244 40236
rect 20524 39732 20580 40348
rect 20636 40292 20692 41916
rect 20748 41906 20804 41916
rect 20748 41748 20804 41758
rect 20748 41654 20804 41692
rect 20972 41524 21028 48414
rect 21420 48132 21476 48142
rect 21476 48076 21588 48132
rect 21420 48038 21476 48076
rect 21308 47460 21364 47470
rect 21308 47366 21364 47404
rect 21420 47234 21476 47246
rect 21420 47182 21422 47234
rect 21474 47182 21476 47234
rect 21196 47124 21252 47134
rect 21420 47124 21476 47182
rect 21252 47068 21476 47124
rect 21196 47058 21252 47068
rect 21308 46676 21364 46686
rect 21420 46676 21476 47068
rect 21532 47124 21588 48076
rect 21756 47460 21812 47470
rect 21532 47058 21588 47068
rect 21644 47234 21700 47246
rect 21644 47182 21646 47234
rect 21698 47182 21700 47234
rect 21308 46674 21476 46676
rect 21308 46622 21310 46674
rect 21362 46622 21476 46674
rect 21308 46620 21476 46622
rect 21308 46610 21364 46620
rect 21308 45890 21364 45902
rect 21308 45838 21310 45890
rect 21362 45838 21364 45890
rect 21196 43764 21252 43774
rect 20636 40226 20692 40236
rect 20748 41468 21028 41524
rect 21084 42196 21140 42206
rect 21084 41746 21140 42140
rect 21084 41694 21086 41746
rect 21138 41694 21140 41746
rect 20524 39676 20692 39732
rect 19964 39442 20020 39452
rect 20524 39508 20580 39518
rect 20188 39394 20244 39406
rect 20188 39342 20190 39394
rect 20242 39342 20244 39394
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19740 39060 19796 39070
rect 19740 38946 19796 39004
rect 19740 38894 19742 38946
rect 19794 38894 19796 38946
rect 19740 38882 19796 38894
rect 20188 38668 20244 39342
rect 20524 38948 20580 39452
rect 20300 38836 20356 38874
rect 20300 38770 20356 38780
rect 20524 38834 20580 38892
rect 20524 38782 20526 38834
rect 20578 38782 20580 38834
rect 20524 38770 20580 38782
rect 20188 38612 20468 38668
rect 19964 38500 20020 38510
rect 19964 38162 20020 38444
rect 19964 38110 19966 38162
rect 20018 38110 20020 38162
rect 19964 38098 20020 38110
rect 19068 37772 19236 37828
rect 18732 37650 18788 37660
rect 18620 37214 18622 37266
rect 18674 37214 18676 37266
rect 18620 37202 18676 37214
rect 18732 37268 18788 37278
rect 18620 37044 18676 37054
rect 18732 37044 18788 37212
rect 19068 37268 19124 37278
rect 19068 37174 19124 37212
rect 18620 37042 18732 37044
rect 18620 36990 18622 37042
rect 18674 36990 18732 37042
rect 18620 36988 18732 36990
rect 18620 36978 18676 36988
rect 18732 36950 18788 36988
rect 19180 36820 19236 37772
rect 19628 37734 19684 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20076 37492 20132 37502
rect 19628 37266 19684 37278
rect 19628 37214 19630 37266
rect 19682 37214 19684 37266
rect 19628 37156 19684 37214
rect 20076 37266 20132 37436
rect 20076 37214 20078 37266
rect 20130 37214 20132 37266
rect 20076 37202 20132 37214
rect 20300 37380 20356 37390
rect 20300 37266 20356 37324
rect 20300 37214 20302 37266
rect 20354 37214 20356 37266
rect 20300 37202 20356 37214
rect 19628 37090 19684 37100
rect 19852 37156 19908 37166
rect 19852 37062 19908 37100
rect 19404 37044 19460 37054
rect 19180 36754 19236 36764
rect 19292 36932 19348 36942
rect 18956 36482 19012 36494
rect 18956 36430 18958 36482
rect 19010 36430 19012 36482
rect 18956 36260 19012 36430
rect 18508 36204 18788 36260
rect 18396 35870 18398 35922
rect 18450 35870 18452 35922
rect 18396 35858 18452 35870
rect 18620 35924 18676 35934
rect 18620 35830 18676 35868
rect 18508 35586 18564 35598
rect 18508 35534 18510 35586
rect 18562 35534 18564 35586
rect 18508 35140 18564 35534
rect 18508 35074 18564 35084
rect 18620 35476 18676 35486
rect 18172 34974 18174 35026
rect 18226 34974 18228 35026
rect 18172 34962 18228 34974
rect 18620 34804 18676 35420
rect 18732 35028 18788 36204
rect 18956 35922 19012 36204
rect 18956 35870 18958 35922
rect 19010 35870 19012 35922
rect 18956 35858 19012 35870
rect 19068 35812 19124 35822
rect 19068 35718 19124 35756
rect 19292 35588 19348 36876
rect 19404 36482 19460 36988
rect 20188 37044 20244 37054
rect 19404 36430 19406 36482
rect 19458 36430 19460 36482
rect 19404 36418 19460 36430
rect 19740 36484 19796 36494
rect 20076 36484 20132 36494
rect 19740 36482 20132 36484
rect 19740 36430 19742 36482
rect 19794 36430 20078 36482
rect 20130 36430 20132 36482
rect 19740 36428 20132 36430
rect 19740 36418 19796 36428
rect 20076 36418 20132 36428
rect 19516 36260 19572 36270
rect 19516 36166 19572 36204
rect 19836 36092 20100 36102
rect 19516 36036 19572 36046
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19404 35588 19460 35598
rect 19292 35586 19460 35588
rect 19292 35534 19406 35586
rect 19458 35534 19460 35586
rect 19292 35532 19460 35534
rect 19404 35522 19460 35532
rect 18956 35140 19012 35150
rect 18956 35046 19012 35084
rect 18732 34934 18788 34972
rect 18844 34916 18900 34926
rect 18620 34748 18788 34804
rect 17948 34132 18004 34142
rect 17836 34130 18004 34132
rect 17836 34078 17950 34130
rect 18002 34078 18004 34130
rect 17836 34076 18004 34078
rect 17724 34066 17780 34076
rect 17948 34020 18004 34076
rect 17948 33954 18004 33964
rect 18620 34132 18676 34142
rect 17276 33406 17278 33458
rect 17330 33406 17332 33458
rect 17276 33394 17332 33406
rect 17612 33908 17668 33918
rect 16828 33236 16884 33246
rect 16828 33142 16884 33180
rect 15932 31714 15988 31724
rect 16044 31948 16660 32004
rect 14588 31614 14590 31666
rect 14642 31614 14644 31666
rect 14588 31220 14644 31614
rect 15596 31556 15652 31566
rect 15596 31462 15652 31500
rect 15932 31554 15988 31566
rect 15932 31502 15934 31554
rect 15986 31502 15988 31554
rect 15932 31444 15988 31502
rect 15932 31378 15988 31388
rect 14588 31154 14644 31164
rect 15820 30996 15876 31006
rect 16044 30996 16100 31948
rect 16492 31778 16548 31790
rect 16492 31726 16494 31778
rect 16546 31726 16548 31778
rect 16156 31668 16212 31678
rect 16156 31666 16324 31668
rect 16156 31614 16158 31666
rect 16210 31614 16324 31666
rect 16156 31612 16324 31614
rect 16156 31602 16212 31612
rect 15820 30994 16100 30996
rect 15820 30942 15822 30994
rect 15874 30942 16100 30994
rect 15820 30940 16100 30942
rect 16156 30994 16212 31006
rect 16156 30942 16158 30994
rect 16210 30942 16212 30994
rect 15820 30930 15876 30940
rect 16156 30772 16212 30942
rect 16268 30884 16324 31612
rect 16492 31556 16548 31726
rect 16604 31668 16660 31948
rect 17500 31778 17556 31790
rect 17500 31726 17502 31778
rect 17554 31726 17556 31778
rect 16604 31666 16772 31668
rect 16604 31614 16606 31666
rect 16658 31614 16772 31666
rect 16604 31612 16772 31614
rect 16604 31602 16660 31612
rect 16492 31490 16548 31500
rect 16380 30884 16436 30894
rect 16268 30828 16380 30884
rect 16380 30818 16436 30828
rect 16156 30706 16212 30716
rect 16492 30772 16548 30782
rect 15708 30100 15764 30110
rect 15708 30006 15764 30044
rect 15932 29986 15988 29998
rect 15932 29934 15934 29986
rect 15986 29934 15988 29986
rect 15932 29540 15988 29934
rect 16044 29988 16100 29998
rect 16044 29894 16100 29932
rect 16156 29986 16212 29998
rect 16156 29934 16158 29986
rect 16210 29934 16212 29986
rect 16156 29876 16212 29934
rect 16492 29986 16548 30716
rect 16716 30210 16772 31612
rect 16828 30882 16884 30894
rect 16828 30830 16830 30882
rect 16882 30830 16884 30882
rect 16828 30660 16884 30830
rect 17388 30884 17444 30894
rect 17388 30790 17444 30828
rect 17500 30660 17556 31726
rect 17612 31554 17668 33852
rect 18060 33346 18116 33358
rect 18060 33294 18062 33346
rect 18114 33294 18116 33346
rect 17948 33124 18004 33134
rect 17948 33030 18004 33068
rect 17836 31780 17892 31790
rect 17612 31502 17614 31554
rect 17666 31502 17668 31554
rect 17612 31490 17668 31502
rect 17724 31554 17780 31566
rect 17724 31502 17726 31554
rect 17778 31502 17780 31554
rect 17724 31444 17780 31502
rect 17724 31378 17780 31388
rect 17836 31220 17892 31724
rect 17836 30994 17892 31164
rect 17836 30942 17838 30994
rect 17890 30942 17892 30994
rect 17836 30930 17892 30942
rect 16828 30604 17556 30660
rect 17948 30884 18004 30894
rect 16716 30158 16718 30210
rect 16770 30158 16772 30210
rect 16716 30146 16772 30158
rect 17164 30210 17220 30222
rect 17164 30158 17166 30210
rect 17218 30158 17220 30210
rect 16604 30100 16660 30110
rect 16604 30006 16660 30044
rect 16492 29934 16494 29986
rect 16546 29934 16548 29986
rect 16492 29922 16548 29934
rect 16156 29810 16212 29820
rect 15932 29474 15988 29484
rect 15036 29316 15092 29326
rect 15484 29316 15540 29326
rect 15036 29314 15428 29316
rect 15036 29262 15038 29314
rect 15090 29262 15428 29314
rect 15036 29260 15428 29262
rect 15036 29250 15092 29260
rect 14476 27918 14478 27970
rect 14530 27918 14532 27970
rect 14476 27906 14532 27918
rect 13804 27806 13806 27858
rect 13858 27806 13860 27858
rect 13804 27794 13860 27806
rect 13468 26962 13524 26974
rect 13468 26910 13470 26962
rect 13522 26910 13524 26962
rect 13468 26908 13524 26910
rect 13804 26962 13860 26974
rect 13804 26910 13806 26962
rect 13858 26910 13860 26962
rect 13804 26908 13860 26910
rect 13132 26852 13524 26908
rect 13580 26852 13860 26908
rect 13132 26402 13188 26852
rect 13132 26350 13134 26402
rect 13186 26350 13188 26402
rect 13132 26338 13188 26350
rect 12404 26236 13076 26292
rect 12348 26198 12404 26236
rect 12236 25732 12292 25742
rect 12236 25506 12292 25676
rect 12796 25732 12852 25742
rect 12796 25618 12852 25676
rect 12796 25566 12798 25618
rect 12850 25566 12852 25618
rect 12796 25554 12852 25566
rect 12236 25454 12238 25506
rect 12290 25454 12292 25506
rect 12236 25442 12292 25454
rect 12124 25396 12180 25406
rect 12124 23938 12180 25340
rect 12908 25396 12964 25406
rect 12572 24610 12628 24622
rect 12572 24558 12574 24610
rect 12626 24558 12628 24610
rect 12572 24052 12628 24558
rect 12124 23886 12126 23938
rect 12178 23886 12180 23938
rect 12124 23874 12180 23886
rect 12236 23996 12628 24052
rect 12236 23826 12292 23996
rect 12236 23774 12238 23826
rect 12290 23774 12292 23826
rect 12236 23268 12292 23774
rect 12908 23378 12964 25340
rect 13020 24946 13076 26236
rect 13580 25730 13636 26852
rect 13580 25678 13582 25730
rect 13634 25678 13636 25730
rect 13580 25666 13636 25678
rect 13916 26516 13972 26526
rect 13916 25730 13972 26460
rect 13916 25678 13918 25730
rect 13970 25678 13972 25730
rect 13916 25620 13972 25678
rect 13916 25554 13972 25564
rect 15260 26178 15316 26190
rect 15260 26126 15262 26178
rect 15314 26126 15316 26178
rect 14140 25396 14196 25406
rect 14140 25302 14196 25340
rect 14700 25396 14756 25406
rect 13020 24894 13022 24946
rect 13074 24894 13076 24946
rect 13020 24882 13076 24894
rect 14700 24164 14756 25340
rect 15260 25396 15316 26126
rect 15260 25330 15316 25340
rect 14924 24164 14980 24174
rect 14700 24162 14980 24164
rect 14700 24110 14926 24162
rect 14978 24110 14980 24162
rect 14700 24108 14980 24110
rect 14924 24098 14980 24108
rect 15372 24052 15428 29260
rect 15484 28644 15540 29260
rect 16828 29316 16884 29326
rect 16380 28756 16436 28766
rect 16380 28754 16548 28756
rect 16380 28702 16382 28754
rect 16434 28702 16548 28754
rect 16380 28700 16548 28702
rect 16380 28690 16436 28700
rect 15484 26908 15540 28588
rect 16380 27074 16436 27086
rect 16380 27022 16382 27074
rect 16434 27022 16436 27074
rect 16380 26908 16436 27022
rect 15484 26852 15764 26908
rect 15708 26514 15764 26852
rect 15708 26462 15710 26514
rect 15762 26462 15764 26514
rect 15708 26450 15764 26462
rect 16156 26852 16436 26908
rect 16492 26908 16548 28700
rect 16828 28754 16884 29260
rect 17164 29092 17220 30158
rect 17388 30210 17444 30604
rect 17388 30158 17390 30210
rect 17442 30158 17444 30210
rect 17388 30146 17444 30158
rect 17388 29988 17444 29998
rect 17388 29426 17444 29932
rect 17388 29374 17390 29426
rect 17442 29374 17444 29426
rect 17388 29362 17444 29374
rect 17948 29876 18004 30828
rect 17948 29426 18004 29820
rect 18060 29764 18116 33294
rect 18284 33124 18340 33134
rect 18284 32562 18340 33068
rect 18284 32510 18286 32562
rect 18338 32510 18340 32562
rect 18284 32498 18340 32510
rect 18396 31780 18452 31790
rect 18396 31444 18452 31724
rect 18396 31378 18452 31388
rect 18284 30884 18340 30894
rect 18284 30790 18340 30828
rect 18620 30434 18676 34076
rect 18732 33684 18788 34748
rect 18732 33234 18788 33628
rect 18844 33346 18900 34860
rect 19292 34916 19348 34926
rect 19516 34916 19572 35980
rect 20188 35924 20244 36988
rect 20300 36258 20356 36270
rect 20300 36206 20302 36258
rect 20354 36206 20356 36258
rect 20300 36148 20356 36206
rect 20300 36082 20356 36092
rect 20188 35858 20244 35868
rect 19292 34914 19572 34916
rect 19292 34862 19294 34914
rect 19346 34862 19572 34914
rect 19292 34860 19572 34862
rect 19628 35252 19684 35262
rect 19628 34914 19684 35196
rect 19628 34862 19630 34914
rect 19682 34862 19684 34914
rect 19068 34690 19124 34702
rect 19068 34638 19070 34690
rect 19122 34638 19124 34690
rect 18956 34244 19012 34254
rect 18956 33796 19012 34188
rect 19068 34132 19124 34638
rect 19068 34066 19124 34076
rect 19292 33796 19348 34860
rect 19012 33740 19124 33796
rect 18956 33730 19012 33740
rect 18844 33294 18846 33346
rect 18898 33294 18900 33346
rect 18844 33282 18900 33294
rect 18732 33182 18734 33234
rect 18786 33182 18788 33234
rect 18732 33170 18788 33182
rect 18956 32450 19012 32462
rect 18956 32398 18958 32450
rect 19010 32398 19012 32450
rect 18956 31890 19012 32398
rect 18956 31838 18958 31890
rect 19010 31838 19012 31890
rect 18956 31826 19012 31838
rect 19068 31778 19124 33740
rect 19292 33730 19348 33740
rect 19404 33684 19460 33694
rect 19404 33458 19460 33628
rect 19404 33406 19406 33458
rect 19458 33406 19460 33458
rect 19404 33394 19460 33406
rect 19068 31726 19070 31778
rect 19122 31726 19124 31778
rect 19068 31714 19124 31726
rect 18732 31668 18788 31678
rect 18732 31574 18788 31612
rect 18732 31220 18788 31230
rect 18732 30994 18788 31164
rect 18732 30942 18734 30994
rect 18786 30942 18788 30994
rect 18732 30930 18788 30942
rect 19068 30884 19124 30894
rect 19068 30790 19124 30828
rect 18732 30772 18788 30782
rect 18732 30678 18788 30716
rect 18620 30382 18622 30434
rect 18674 30382 18676 30434
rect 18620 30370 18676 30382
rect 18060 29698 18116 29708
rect 18396 30212 18452 30222
rect 18060 29540 18116 29550
rect 18116 29484 18340 29540
rect 18060 29446 18116 29484
rect 17948 29374 17950 29426
rect 18002 29374 18004 29426
rect 17948 29362 18004 29374
rect 17164 29026 17220 29036
rect 17836 29092 17892 29102
rect 16828 28702 16830 28754
rect 16882 28702 16884 28754
rect 16828 28084 16884 28702
rect 16828 28018 16884 28028
rect 17500 28084 17556 28094
rect 17500 27990 17556 28028
rect 16604 27748 16660 27758
rect 16604 27746 16772 27748
rect 16604 27694 16606 27746
rect 16658 27694 16772 27746
rect 16604 27692 16772 27694
rect 16604 27682 16660 27692
rect 16716 26908 16772 27692
rect 17164 27636 17220 27646
rect 17164 27186 17220 27580
rect 17164 27134 17166 27186
rect 17218 27134 17220 27186
rect 17164 27122 17220 27134
rect 16492 26852 16660 26908
rect 16716 26852 17220 26908
rect 15484 25620 15540 25630
rect 15484 24946 15540 25564
rect 15596 25508 15652 25518
rect 16156 25508 16212 26852
rect 15596 25506 16212 25508
rect 15596 25454 15598 25506
rect 15650 25454 16212 25506
rect 15596 25452 16212 25454
rect 15596 25442 15652 25452
rect 16156 25172 16212 25452
rect 16156 25106 16212 25116
rect 16268 25394 16324 25406
rect 16268 25342 16270 25394
rect 16322 25342 16324 25394
rect 15484 24894 15486 24946
rect 15538 24894 15540 24946
rect 15484 24882 15540 24894
rect 16268 24948 16324 25342
rect 16268 24882 16324 24892
rect 15820 24724 15876 24734
rect 15820 24630 15876 24668
rect 16268 24724 16324 24734
rect 16268 24630 16324 24668
rect 15372 23996 15652 24052
rect 15148 23826 15204 23838
rect 15148 23774 15150 23826
rect 15202 23774 15204 23826
rect 13804 23716 13860 23726
rect 12908 23326 12910 23378
rect 12962 23326 12964 23378
rect 12908 23314 12964 23326
rect 13468 23714 14084 23716
rect 13468 23662 13806 23714
rect 13858 23662 14084 23714
rect 13468 23660 14084 23662
rect 12348 23268 12404 23278
rect 13468 23268 13524 23660
rect 13804 23650 13860 23660
rect 12236 23212 12348 23268
rect 12348 23202 12404 23212
rect 13244 23212 13524 23268
rect 13692 23492 13748 23502
rect 13244 23154 13300 23212
rect 13244 23102 13246 23154
rect 13298 23102 13300 23154
rect 13244 23090 13300 23102
rect 12572 23044 12628 23054
rect 12460 22988 12572 23044
rect 12236 21588 12292 21598
rect 12236 21494 12292 21532
rect 12348 21476 12404 21486
rect 12348 21026 12404 21420
rect 12348 20974 12350 21026
rect 12402 20974 12404 21026
rect 12348 20962 12404 20974
rect 12348 20802 12404 20814
rect 12348 20750 12350 20802
rect 12402 20750 12404 20802
rect 12348 20692 12404 20750
rect 12348 20626 12404 20636
rect 11900 20076 12068 20132
rect 11900 20018 11956 20076
rect 11900 19966 11902 20018
rect 11954 19966 11956 20018
rect 11900 19954 11956 19966
rect 11900 19794 11956 19806
rect 12460 19796 12516 22988
rect 12572 22950 12628 22988
rect 13468 23042 13524 23054
rect 13468 22990 13470 23042
rect 13522 22990 13524 23042
rect 13468 22932 13524 22990
rect 13692 22932 13748 23436
rect 13916 23268 13972 23278
rect 13804 23154 13860 23166
rect 13804 23102 13806 23154
rect 13858 23102 13860 23154
rect 13804 23044 13860 23102
rect 13804 22978 13860 22988
rect 13524 22876 13748 22932
rect 13468 22866 13524 22876
rect 13580 22596 13636 22606
rect 13468 22594 13636 22596
rect 13468 22542 13582 22594
rect 13634 22542 13636 22594
rect 13468 22540 13636 22542
rect 12572 22482 12628 22494
rect 12572 22430 12574 22482
rect 12626 22430 12628 22482
rect 12572 21588 12628 22430
rect 12908 22260 12964 22270
rect 12572 21522 12628 21532
rect 12796 21698 12852 21710
rect 12796 21646 12798 21698
rect 12850 21646 12852 21698
rect 12796 21252 12852 21646
rect 12908 21586 12964 22204
rect 13468 22260 13524 22540
rect 13580 22530 13636 22540
rect 13692 22372 13748 22876
rect 13468 22194 13524 22204
rect 13580 22316 13748 22372
rect 13804 22596 13860 22606
rect 13580 22258 13636 22316
rect 13804 22260 13860 22540
rect 13580 22206 13582 22258
rect 13634 22206 13636 22258
rect 13580 22194 13636 22206
rect 13692 22204 13860 22260
rect 13692 22202 13748 22204
rect 12908 21534 12910 21586
rect 12962 21534 12964 21586
rect 12908 21522 12964 21534
rect 13692 22150 13694 22202
rect 13746 22150 13748 22202
rect 12796 21186 12852 21196
rect 13580 21362 13636 21374
rect 13580 21310 13582 21362
rect 13634 21310 13636 21362
rect 12908 20804 12964 20814
rect 12908 20710 12964 20748
rect 13580 20804 13636 21310
rect 13580 20738 13636 20748
rect 11900 19742 11902 19794
rect 11954 19742 11956 19794
rect 11900 19234 11956 19742
rect 11900 19182 11902 19234
rect 11954 19182 11956 19234
rect 11900 19170 11956 19182
rect 12012 19740 12516 19796
rect 12572 20692 12628 20702
rect 11564 18226 11732 18228
rect 11564 18174 11566 18226
rect 11618 18174 11732 18226
rect 11564 18172 11732 18174
rect 11900 19010 11956 19022
rect 11900 18958 11902 19010
rect 11954 18958 11956 19010
rect 11564 18162 11620 18172
rect 11900 17892 11956 18958
rect 11900 17826 11956 17836
rect 11340 17054 11342 17106
rect 11394 17054 11396 17106
rect 11340 17042 11396 17054
rect 11116 16818 11172 16828
rect 11788 16884 11844 16894
rect 12012 16884 12068 19740
rect 12572 19684 12628 20636
rect 12684 20690 12740 20702
rect 12684 20638 12686 20690
rect 12738 20638 12740 20690
rect 12684 20580 12740 20638
rect 12684 20514 12740 20524
rect 12796 20578 12852 20590
rect 12796 20526 12798 20578
rect 12850 20526 12852 20578
rect 12348 19628 12628 19684
rect 12348 18676 12404 19628
rect 12796 19460 12852 20526
rect 13692 20020 13748 22150
rect 13916 21586 13972 23212
rect 13916 21534 13918 21586
rect 13970 21534 13972 21586
rect 13916 21522 13972 21534
rect 12796 19394 12852 19404
rect 13468 19964 13748 20020
rect 12348 18620 12740 18676
rect 12348 18450 12404 18620
rect 12348 18398 12350 18450
rect 12402 18398 12404 18450
rect 12348 18386 12404 18398
rect 12460 18452 12516 18462
rect 12460 18226 12516 18396
rect 12460 18174 12462 18226
rect 12514 18174 12516 18226
rect 12460 18162 12516 18174
rect 12572 17892 12628 17902
rect 12572 17798 12628 17836
rect 12460 17666 12516 17678
rect 12460 17614 12462 17666
rect 12514 17614 12516 17666
rect 11788 16882 12068 16884
rect 11788 16830 11790 16882
rect 11842 16830 12068 16882
rect 11788 16828 12068 16830
rect 12124 17554 12180 17566
rect 12124 17502 12126 17554
rect 12178 17502 12180 17554
rect 11228 16770 11284 16782
rect 11228 16718 11230 16770
rect 11282 16718 11284 16770
rect 11116 16212 11172 16222
rect 11228 16212 11284 16718
rect 11116 16210 11284 16212
rect 11116 16158 11118 16210
rect 11170 16158 11284 16210
rect 11116 16156 11284 16158
rect 11676 16324 11732 16334
rect 11116 15316 11172 16156
rect 11564 15876 11620 15886
rect 11564 15782 11620 15820
rect 11452 15316 11508 15326
rect 11116 15314 11508 15316
rect 11116 15262 11454 15314
rect 11506 15262 11508 15314
rect 11116 15260 11508 15262
rect 11452 15250 11508 15260
rect 11004 14702 11006 14754
rect 11058 14702 11060 14754
rect 11004 14690 11060 14702
rect 11116 15090 11172 15102
rect 11116 15038 11118 15090
rect 11170 15038 11172 15090
rect 9884 14644 9940 14654
rect 9884 14550 9940 14588
rect 10892 14644 10948 14654
rect 10892 14550 10948 14588
rect 10220 14420 10276 14430
rect 10220 14326 10276 14364
rect 10556 14418 10612 14430
rect 10556 14366 10558 14418
rect 10610 14366 10612 14418
rect 10556 14196 10612 14366
rect 11116 14196 11172 15038
rect 11676 14754 11732 16268
rect 11676 14702 11678 14754
rect 11730 14702 11732 14754
rect 11676 14690 11732 14702
rect 10556 14140 11172 14196
rect 11228 14308 11284 14318
rect 9996 13746 10052 13758
rect 9996 13694 9998 13746
rect 10050 13694 10052 13746
rect 9996 13412 10052 13694
rect 10668 13636 10724 13646
rect 10668 13542 10724 13580
rect 9996 13346 10052 13356
rect 9772 13234 9828 13244
rect 11228 13076 11284 14252
rect 11788 13972 11844 16828
rect 12124 16324 12180 17502
rect 12460 17444 12516 17614
rect 12684 17666 12740 18620
rect 12908 18562 12964 18574
rect 12908 18510 12910 18562
rect 12962 18510 12964 18562
rect 12684 17614 12686 17666
rect 12738 17614 12740 17666
rect 12684 17602 12740 17614
rect 12796 18452 12852 18462
rect 12796 17444 12852 18396
rect 12908 18340 12964 18510
rect 13356 18564 13412 18574
rect 13020 18452 13076 18462
rect 13020 18450 13188 18452
rect 13020 18398 13022 18450
rect 13074 18398 13188 18450
rect 13020 18396 13188 18398
rect 13020 18386 13076 18396
rect 12908 18274 12964 18284
rect 12460 17388 12852 17444
rect 12908 17780 12964 17790
rect 12908 17442 12964 17724
rect 12908 17390 12910 17442
rect 12962 17390 12964 17442
rect 12460 16884 12516 17388
rect 12908 17378 12964 17390
rect 12460 16818 12516 16828
rect 12796 16882 12852 16894
rect 12796 16830 12798 16882
rect 12850 16830 12852 16882
rect 12124 16258 12180 16268
rect 11900 16100 11956 16110
rect 11900 16098 12068 16100
rect 11900 16046 11902 16098
rect 11954 16046 12068 16098
rect 11900 16044 12068 16046
rect 11900 16034 11956 16044
rect 12012 15652 12068 16044
rect 12236 15986 12292 15998
rect 12236 15934 12238 15986
rect 12290 15934 12292 15986
rect 12012 15596 12180 15652
rect 12012 15428 12068 15438
rect 12012 15334 12068 15372
rect 12124 15148 12180 15596
rect 12236 15540 12292 15934
rect 12460 15988 12516 15998
rect 12460 15894 12516 15932
rect 12796 15764 12852 16830
rect 13020 16884 13076 16894
rect 13020 16790 13076 16828
rect 12908 16770 12964 16782
rect 12908 16718 12910 16770
rect 12962 16718 12964 16770
rect 12908 16660 12964 16718
rect 12908 16594 12964 16604
rect 12684 15708 12852 15764
rect 12572 15540 12628 15550
rect 12236 15538 12628 15540
rect 12236 15486 12574 15538
rect 12626 15486 12628 15538
rect 12236 15484 12628 15486
rect 12236 15314 12292 15484
rect 12572 15474 12628 15484
rect 12236 15262 12238 15314
rect 12290 15262 12292 15314
rect 12236 15250 12292 15262
rect 11900 15092 12180 15148
rect 11900 14644 11956 15092
rect 11900 14578 11956 14588
rect 11788 13906 11844 13916
rect 12012 14530 12068 14542
rect 12012 14478 12014 14530
rect 12066 14478 12068 14530
rect 11228 13010 11284 13020
rect 11340 13524 11396 13534
rect 9548 12852 9604 12862
rect 9548 12850 9940 12852
rect 9548 12798 9550 12850
rect 9602 12798 9940 12850
rect 9548 12796 9940 12798
rect 9548 12786 9604 12796
rect 9436 12572 9828 12628
rect 8988 11508 9044 11518
rect 8932 11506 9044 11508
rect 8932 11454 8990 11506
rect 9042 11454 9044 11506
rect 8932 11452 9044 11454
rect 8876 11442 8932 11452
rect 8988 11442 9044 11452
rect 9548 11508 9604 11518
rect 8540 11218 8596 11228
rect 9548 11394 9604 11452
rect 9548 11342 9550 11394
rect 9602 11342 9604 11394
rect 8316 9662 8318 9714
rect 8370 9662 8372 9714
rect 8316 9650 8372 9662
rect 8988 9716 9044 9726
rect 7644 8866 7700 8876
rect 8988 8932 9044 9660
rect 8988 8838 9044 8876
rect 9548 9042 9604 11342
rect 9548 8990 9550 9042
rect 9602 8990 9604 9042
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 9548 8428 9604 8990
rect 9212 8372 9716 8428
rect 9212 8370 9268 8372
rect 9212 8318 9214 8370
rect 9266 8318 9268 8370
rect 9212 8306 9268 8318
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 9660 6804 9716 8372
rect 9772 8372 9828 12572
rect 9884 12402 9940 12796
rect 9884 12350 9886 12402
rect 9938 12350 9940 12402
rect 9884 12338 9940 12350
rect 10892 12740 10948 12750
rect 10556 12292 10612 12302
rect 10332 12290 10612 12292
rect 10332 12238 10558 12290
rect 10610 12238 10612 12290
rect 10332 12236 10612 12238
rect 10220 12180 10276 12190
rect 10220 12086 10276 12124
rect 10332 11506 10388 12236
rect 10556 12226 10612 12236
rect 10892 12290 10948 12684
rect 11340 12628 11396 13468
rect 11676 13188 11732 13198
rect 11676 13074 11732 13132
rect 11676 13022 11678 13074
rect 11730 13022 11732 13074
rect 11676 13010 11732 13022
rect 12012 12964 12068 14478
rect 12012 12898 12068 12908
rect 12236 14418 12292 14430
rect 12236 14366 12238 14418
rect 12290 14366 12292 14418
rect 12236 13860 12292 14366
rect 11340 12562 11396 12572
rect 10892 12238 10894 12290
rect 10946 12238 10948 12290
rect 10892 12226 10948 12238
rect 10332 11454 10334 11506
rect 10386 11454 10388 11506
rect 10332 11442 10388 11454
rect 11452 10386 11508 10398
rect 11452 10334 11454 10386
rect 11506 10334 11508 10386
rect 9772 8306 9828 8316
rect 10332 8930 10388 8942
rect 10332 8878 10334 8930
rect 10386 8878 10388 8930
rect 10332 8146 10388 8878
rect 11452 8428 11508 10334
rect 10668 8372 11508 8428
rect 11788 10386 11844 10398
rect 11788 10334 11790 10386
rect 11842 10334 11844 10386
rect 11788 8428 11844 10334
rect 11900 9716 11956 9726
rect 11900 9622 11956 9660
rect 12236 9714 12292 13804
rect 12572 14418 12628 14430
rect 12572 14366 12574 14418
rect 12626 14366 12628 14418
rect 12460 13412 12516 13422
rect 12460 13074 12516 13356
rect 12460 13022 12462 13074
rect 12514 13022 12516 13074
rect 12460 13010 12516 13022
rect 12572 13188 12628 14366
rect 12572 12404 12628 13132
rect 12460 12348 12628 12404
rect 12348 12180 12404 12190
rect 12348 12086 12404 12124
rect 12460 12068 12516 12348
rect 12684 12292 12740 15708
rect 12796 15540 12852 15550
rect 12796 15446 12852 15484
rect 12796 15316 12852 15326
rect 12796 14084 12852 15260
rect 12796 13970 12852 14028
rect 12796 13918 12798 13970
rect 12850 13918 12852 13970
rect 12796 13906 12852 13918
rect 12908 15314 12964 15326
rect 12908 15262 12910 15314
rect 12962 15262 12964 15314
rect 12908 14532 12964 15262
rect 12908 13858 12964 14476
rect 13132 13972 13188 18396
rect 13356 18450 13412 18508
rect 13356 18398 13358 18450
rect 13410 18398 13412 18450
rect 13356 18386 13412 18398
rect 13244 18228 13300 18238
rect 13244 16770 13300 18172
rect 13468 18004 13524 19964
rect 13692 19796 13748 19806
rect 13580 18564 13636 18574
rect 13580 18470 13636 18508
rect 13468 17938 13524 17948
rect 13244 16718 13246 16770
rect 13298 16718 13300 16770
rect 13244 16706 13300 16718
rect 13580 16882 13636 16894
rect 13580 16830 13582 16882
rect 13634 16830 13636 16882
rect 13132 13906 13188 13916
rect 13356 16212 13412 16222
rect 13356 15428 13412 16156
rect 13580 16100 13636 16830
rect 13692 16436 13748 19740
rect 13804 19012 13860 19022
rect 14028 19012 14084 23660
rect 14252 23714 14308 23726
rect 14252 23662 14254 23714
rect 14306 23662 14308 23714
rect 14252 22596 14308 23662
rect 14588 23716 14644 23726
rect 14588 23714 14980 23716
rect 14588 23662 14590 23714
rect 14642 23662 14980 23714
rect 14588 23660 14980 23662
rect 14588 23650 14644 23660
rect 14588 23044 14644 23054
rect 14252 22530 14308 22540
rect 14364 23042 14644 23044
rect 14364 22990 14590 23042
rect 14642 22990 14644 23042
rect 14364 22988 14644 22990
rect 14140 22370 14196 22382
rect 14140 22318 14142 22370
rect 14194 22318 14196 22370
rect 14140 22036 14196 22318
rect 14364 22258 14420 22988
rect 14588 22978 14644 22988
rect 14364 22206 14366 22258
rect 14418 22206 14420 22258
rect 14364 22194 14420 22206
rect 14812 22146 14868 22158
rect 14812 22094 14814 22146
rect 14866 22094 14868 22146
rect 14812 22036 14868 22094
rect 14140 21980 14868 22036
rect 14476 21698 14532 21710
rect 14476 21646 14478 21698
rect 14530 21646 14532 21698
rect 14476 21588 14532 21646
rect 14476 21522 14532 21532
rect 14700 21586 14756 21598
rect 14700 21534 14702 21586
rect 14754 21534 14756 21586
rect 14700 21476 14756 21534
rect 14700 21410 14756 21420
rect 14364 21028 14420 21038
rect 14364 20934 14420 20972
rect 14364 20804 14420 20814
rect 14364 20710 14420 20748
rect 14924 20802 14980 23660
rect 15148 22820 15204 23774
rect 15148 22754 15204 22764
rect 15484 23826 15540 23838
rect 15484 23774 15486 23826
rect 15538 23774 15540 23826
rect 15484 23044 15540 23774
rect 15148 22596 15204 22606
rect 15484 22596 15540 22988
rect 15148 22594 15540 22596
rect 15148 22542 15150 22594
rect 15202 22542 15540 22594
rect 15148 22540 15540 22542
rect 15148 22530 15204 22540
rect 15372 22260 15428 22270
rect 15372 22166 15428 22204
rect 15260 21476 15316 21486
rect 15316 21420 15428 21476
rect 15260 21382 15316 21420
rect 14924 20750 14926 20802
rect 14978 20750 14980 20802
rect 14924 20738 14980 20750
rect 15260 20804 15316 20814
rect 14700 20690 14756 20702
rect 14700 20638 14702 20690
rect 14754 20638 14756 20690
rect 14700 20580 14756 20638
rect 15260 20690 15316 20748
rect 15260 20638 15262 20690
rect 15314 20638 15316 20690
rect 15260 20626 15316 20638
rect 13804 18450 13860 18956
rect 13804 18398 13806 18450
rect 13858 18398 13860 18450
rect 13804 18386 13860 18398
rect 13916 18956 14084 19012
rect 14364 20018 14420 20030
rect 14364 19966 14366 20018
rect 14418 19966 14420 20018
rect 13916 17220 13972 18956
rect 14364 18900 14420 19966
rect 14588 20020 14644 20030
rect 14700 20020 14756 20524
rect 14812 20578 14868 20590
rect 14812 20526 14814 20578
rect 14866 20526 14868 20578
rect 14812 20244 14868 20526
rect 14812 20178 14868 20188
rect 14924 20020 14980 20030
rect 14700 20018 14980 20020
rect 14700 19966 14926 20018
rect 14978 19966 14980 20018
rect 14700 19964 14980 19966
rect 14588 19794 14644 19964
rect 14588 19742 14590 19794
rect 14642 19742 14644 19794
rect 14588 19730 14644 19742
rect 14476 19460 14532 19470
rect 14476 19234 14532 19404
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 14476 19170 14532 19182
rect 14700 19234 14756 19246
rect 14700 19182 14702 19234
rect 14754 19182 14756 19234
rect 14028 18844 14420 18900
rect 14028 18452 14084 18844
rect 14140 18676 14196 18686
rect 14700 18676 14756 19182
rect 14140 18674 14756 18676
rect 14140 18622 14142 18674
rect 14194 18622 14756 18674
rect 14140 18620 14756 18622
rect 14140 18610 14196 18620
rect 14812 18564 14868 19964
rect 14924 19954 14980 19964
rect 15036 20020 15092 20030
rect 15036 19926 15092 19964
rect 15148 20020 15204 20030
rect 15148 20018 15316 20020
rect 15148 19966 15150 20018
rect 15202 19966 15316 20018
rect 15148 19964 15316 19966
rect 15148 19954 15204 19964
rect 14924 19796 14980 19806
rect 14924 19458 14980 19740
rect 14924 19406 14926 19458
rect 14978 19406 14980 19458
rect 14924 19394 14980 19406
rect 15036 19236 15092 19246
rect 15036 19142 15092 19180
rect 14588 18508 14868 18564
rect 14140 18452 14196 18462
rect 14028 18450 14196 18452
rect 14028 18398 14142 18450
rect 14194 18398 14196 18450
rect 14028 18396 14196 18398
rect 13916 17154 13972 17164
rect 14140 17666 14196 18396
rect 14476 18340 14532 18350
rect 14140 17614 14142 17666
rect 14194 17614 14196 17666
rect 13916 16884 13972 16894
rect 13804 16436 13860 16446
rect 13692 16380 13804 16436
rect 13804 16370 13860 16380
rect 13580 16034 13636 16044
rect 13916 15986 13972 16828
rect 14140 16100 14196 17614
rect 14364 17666 14420 17678
rect 14364 17614 14366 17666
rect 14418 17614 14420 17666
rect 14364 17444 14420 17614
rect 14364 17378 14420 17388
rect 14140 16034 14196 16044
rect 14252 16884 14308 16894
rect 14252 16098 14308 16828
rect 14476 16882 14532 18284
rect 14476 16830 14478 16882
rect 14530 16830 14532 16882
rect 14476 16818 14532 16830
rect 14588 17554 14644 18508
rect 14700 17668 14756 17678
rect 14700 17574 14756 17612
rect 15148 17668 15204 17678
rect 15148 17574 15204 17612
rect 14588 17502 14590 17554
rect 14642 17502 14644 17554
rect 14588 16772 14644 17502
rect 14812 17556 14868 17566
rect 15260 17556 15316 19964
rect 15372 19796 15428 21420
rect 15596 20802 15652 23996
rect 16156 22820 16212 22830
rect 15932 22258 15988 22270
rect 15932 22206 15934 22258
rect 15986 22206 15988 22258
rect 15932 22036 15988 22206
rect 15932 21970 15988 21980
rect 16156 21586 16212 22764
rect 16156 21534 16158 21586
rect 16210 21534 16212 21586
rect 16156 21522 16212 21534
rect 15596 20750 15598 20802
rect 15650 20750 15652 20802
rect 15484 20132 15540 20142
rect 15484 20018 15540 20076
rect 15484 19966 15486 20018
rect 15538 19966 15540 20018
rect 15484 19954 15540 19966
rect 15372 19740 15540 19796
rect 15372 17780 15428 17790
rect 15372 17686 15428 17724
rect 14812 17554 15092 17556
rect 14812 17502 14814 17554
rect 14866 17502 15092 17554
rect 14812 17500 15092 17502
rect 15260 17500 15428 17556
rect 14812 17490 14868 17500
rect 14588 16706 14644 16716
rect 14700 17444 14756 17454
rect 14700 16770 14756 17388
rect 14924 17220 14980 17230
rect 14812 16996 14868 17006
rect 14812 16902 14868 16940
rect 14700 16718 14702 16770
rect 14754 16718 14756 16770
rect 14700 16706 14756 16718
rect 14364 16660 14420 16670
rect 14364 16566 14420 16604
rect 14252 16046 14254 16098
rect 14306 16046 14308 16098
rect 14252 16034 14308 16046
rect 14588 16436 14644 16446
rect 13916 15934 13918 15986
rect 13970 15934 13972 15986
rect 13916 15922 13972 15934
rect 14364 15988 14420 15998
rect 14364 15764 14420 15932
rect 14588 15986 14644 16380
rect 14588 15934 14590 15986
rect 14642 15934 14644 15986
rect 14588 15922 14644 15934
rect 14812 16100 14868 16110
rect 13468 15540 13524 15550
rect 13468 15446 13524 15484
rect 12908 13806 12910 13858
rect 12962 13806 12964 13858
rect 12908 13794 12964 13806
rect 12796 13524 12852 13534
rect 12796 13522 12964 13524
rect 12796 13470 12798 13522
rect 12850 13470 12964 13522
rect 12796 13468 12964 13470
rect 12796 13458 12852 13468
rect 12908 12852 12964 13468
rect 12460 12002 12516 12012
rect 12572 12236 12740 12292
rect 12796 12738 12852 12750
rect 12796 12686 12798 12738
rect 12850 12686 12852 12738
rect 12460 11844 12516 11854
rect 12460 11506 12516 11788
rect 12460 11454 12462 11506
rect 12514 11454 12516 11506
rect 12460 11442 12516 11454
rect 12572 11396 12628 12236
rect 12684 12068 12740 12078
rect 12684 11974 12740 12012
rect 12796 11508 12852 12686
rect 12908 12290 12964 12796
rect 12908 12238 12910 12290
rect 12962 12238 12964 12290
rect 12908 12226 12964 12238
rect 13356 12290 13412 15372
rect 13916 15202 13972 15214
rect 13916 15150 13918 15202
rect 13970 15150 13972 15202
rect 13804 14532 13860 14542
rect 13804 14438 13860 14476
rect 13580 14308 13636 14318
rect 13580 14214 13636 14252
rect 13468 14084 13524 14094
rect 13468 13970 13524 14028
rect 13468 13918 13470 13970
rect 13522 13918 13524 13970
rect 13468 13906 13524 13918
rect 13804 13972 13860 13982
rect 13804 13878 13860 13916
rect 13916 13860 13972 15150
rect 14140 14420 14196 14430
rect 14140 14326 14196 14364
rect 13916 13794 13972 13804
rect 14140 13524 14196 13534
rect 14140 13430 14196 13468
rect 13916 12964 13972 12974
rect 13580 12740 13636 12750
rect 13580 12646 13636 12684
rect 13356 12238 13358 12290
rect 13410 12238 13412 12290
rect 13356 12226 13412 12238
rect 13916 11844 13972 12908
rect 14140 12852 14196 12862
rect 14364 12852 14420 15708
rect 14476 15540 14532 15550
rect 14812 15540 14868 16044
rect 14476 15538 14868 15540
rect 14476 15486 14478 15538
rect 14530 15486 14868 15538
rect 14476 15484 14868 15486
rect 14924 15538 14980 17164
rect 14924 15486 14926 15538
rect 14978 15486 14980 15538
rect 14476 15474 14532 15484
rect 14924 14420 14980 15486
rect 14924 14354 14980 14364
rect 14812 14306 14868 14318
rect 14812 14254 14814 14306
rect 14866 14254 14868 14306
rect 14476 13860 14532 13870
rect 14476 13766 14532 13804
rect 14700 13858 14756 13870
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 12964 14756 13806
rect 14700 12898 14756 12908
rect 14476 12852 14532 12862
rect 14364 12850 14532 12852
rect 14364 12798 14478 12850
rect 14530 12798 14532 12850
rect 14364 12796 14532 12798
rect 14140 12758 14196 12796
rect 14476 12786 14532 12796
rect 13916 11778 13972 11788
rect 14812 11620 14868 14254
rect 15036 11620 15092 17500
rect 15148 16994 15204 17006
rect 15148 16942 15150 16994
rect 15202 16942 15204 16994
rect 15148 16772 15204 16942
rect 15148 16706 15204 16716
rect 15260 15988 15316 15998
rect 15260 15894 15316 15932
rect 15148 15876 15204 15886
rect 15148 15652 15204 15820
rect 15148 14754 15204 15596
rect 15372 15148 15428 17500
rect 15484 17500 15540 19740
rect 15596 18004 15652 20750
rect 16380 20130 16436 20142
rect 16380 20078 16382 20130
rect 16434 20078 16436 20130
rect 15708 20020 15764 20030
rect 15708 19926 15764 19964
rect 15932 19796 15988 19806
rect 15932 19702 15988 19740
rect 16044 19794 16100 19806
rect 16044 19742 16046 19794
rect 16098 19742 16100 19794
rect 16044 19460 16100 19742
rect 16380 19684 16436 20078
rect 16604 20020 16660 26852
rect 16828 23716 16884 23726
rect 16828 23714 17108 23716
rect 16828 23662 16830 23714
rect 16882 23662 17108 23714
rect 16828 23660 17108 23662
rect 16828 23650 16884 23660
rect 16716 23044 16772 23054
rect 16716 22950 16772 22988
rect 16716 21586 16772 21598
rect 16716 21534 16718 21586
rect 16770 21534 16772 21586
rect 16716 21476 16772 21534
rect 16716 21410 16772 21420
rect 16940 21476 16996 21486
rect 16604 19926 16660 19964
rect 16380 19628 16660 19684
rect 16492 19460 16548 19470
rect 15932 19404 16100 19460
rect 16380 19404 16492 19460
rect 15708 19236 15764 19246
rect 15708 19142 15764 19180
rect 15932 19012 15988 19404
rect 16156 19234 16212 19246
rect 16156 19182 16158 19234
rect 16210 19182 16212 19234
rect 15932 18956 16100 19012
rect 15932 18452 15988 18462
rect 15596 17938 15652 17948
rect 15820 18450 15988 18452
rect 15820 18398 15934 18450
rect 15986 18398 15988 18450
rect 15820 18396 15988 18398
rect 15708 17892 15764 17902
rect 15820 17892 15876 18396
rect 15932 18386 15988 18396
rect 16044 18338 16100 18956
rect 16044 18286 16046 18338
rect 16098 18286 16100 18338
rect 16044 18274 16100 18286
rect 16156 18450 16212 19182
rect 16380 18674 16436 19404
rect 16492 19394 16548 19404
rect 16380 18622 16382 18674
rect 16434 18622 16436 18674
rect 16380 18610 16436 18622
rect 16492 19234 16548 19246
rect 16492 19182 16494 19234
rect 16546 19182 16548 19234
rect 16156 18398 16158 18450
rect 16210 18398 16212 18450
rect 16156 18340 16212 18398
rect 16156 18274 16212 18284
rect 15708 17890 15876 17892
rect 15708 17838 15710 17890
rect 15762 17838 15876 17890
rect 15708 17836 15876 17838
rect 16044 18004 16100 18014
rect 15708 17826 15764 17836
rect 15596 17668 15652 17678
rect 15596 17574 15652 17612
rect 15484 17444 15652 17500
rect 15484 16884 15540 16894
rect 15484 16790 15540 16828
rect 15596 16660 15652 17444
rect 15484 16604 15652 16660
rect 15820 16994 15876 17006
rect 15820 16942 15822 16994
rect 15874 16942 15876 16994
rect 15484 15652 15540 16604
rect 15820 16212 15876 16942
rect 15820 16146 15876 16156
rect 16044 16324 16100 17948
rect 16156 17780 16212 17790
rect 16156 17332 16212 17724
rect 16156 17106 16212 17276
rect 16156 17054 16158 17106
rect 16210 17054 16212 17106
rect 16156 17042 16212 17054
rect 16492 17108 16548 19182
rect 16604 17668 16660 19628
rect 16716 19458 16772 19470
rect 16716 19406 16718 19458
rect 16770 19406 16772 19458
rect 16716 19236 16772 19406
rect 16716 19170 16772 19180
rect 16940 19012 16996 21420
rect 16604 17602 16660 17612
rect 16716 18956 16996 19012
rect 16492 17042 16548 17052
rect 16604 17444 16660 17454
rect 16716 17444 16772 18956
rect 16940 17892 16996 17902
rect 16940 17554 16996 17836
rect 16940 17502 16942 17554
rect 16994 17502 16996 17554
rect 16940 17490 16996 17502
rect 16604 17442 16772 17444
rect 16604 17390 16606 17442
rect 16658 17390 16772 17442
rect 16604 17388 16772 17390
rect 16604 16996 16660 17388
rect 16604 16882 16660 16940
rect 16604 16830 16606 16882
rect 16658 16830 16660 16882
rect 16604 16818 16660 16830
rect 16828 16994 16884 17006
rect 16828 16942 16830 16994
rect 16882 16942 16884 16994
rect 16828 16772 16884 16942
rect 16716 16660 16772 16670
rect 16044 16210 16100 16268
rect 16044 16158 16046 16210
rect 16098 16158 16100 16210
rect 16044 16146 16100 16158
rect 16380 16324 16436 16334
rect 16380 16098 16436 16268
rect 16380 16046 16382 16098
rect 16434 16046 16436 16098
rect 16380 16034 16436 16046
rect 15596 15986 15652 15998
rect 15596 15934 15598 15986
rect 15650 15934 15652 15986
rect 15596 15876 15652 15934
rect 16716 15986 16772 16604
rect 16828 16100 16884 16716
rect 16828 16034 16884 16044
rect 16716 15934 16718 15986
rect 16770 15934 16772 15986
rect 16716 15922 16772 15934
rect 15932 15876 15988 15886
rect 15596 15874 15988 15876
rect 15596 15822 15934 15874
rect 15986 15822 15988 15874
rect 15596 15820 15988 15822
rect 15484 15596 15764 15652
rect 15148 14702 15150 14754
rect 15202 14702 15204 14754
rect 15148 14690 15204 14702
rect 15260 15092 15428 15148
rect 15596 15204 15652 15242
rect 15148 11620 15204 11630
rect 15036 11618 15204 11620
rect 15036 11566 15150 11618
rect 15202 11566 15204 11618
rect 15036 11564 15204 11566
rect 14812 11554 14868 11564
rect 15148 11554 15204 11564
rect 12908 11508 12964 11518
rect 12796 11506 13188 11508
rect 12796 11454 12910 11506
rect 12962 11454 13188 11506
rect 12796 11452 13188 11454
rect 12908 11442 12964 11452
rect 12572 11340 12852 11396
rect 12236 9662 12238 9714
rect 12290 9662 12292 9714
rect 11788 8372 11956 8428
rect 10668 8258 10724 8372
rect 10668 8206 10670 8258
rect 10722 8206 10724 8258
rect 10668 8194 10724 8206
rect 11900 8260 11956 8372
rect 11900 8194 11956 8204
rect 10332 8094 10334 8146
rect 10386 8094 10388 8146
rect 10332 8082 10388 8094
rect 12236 8148 12292 9662
rect 12460 10722 12516 10734
rect 12460 10670 12462 10722
rect 12514 10670 12516 10722
rect 12460 10050 12516 10670
rect 12572 10724 12628 10734
rect 12572 10610 12628 10668
rect 12572 10558 12574 10610
rect 12626 10558 12628 10610
rect 12572 10546 12628 10558
rect 12460 9998 12462 10050
rect 12514 9998 12516 10050
rect 12460 8930 12516 9998
rect 12796 10050 12852 11340
rect 13132 10836 13188 11452
rect 14588 11396 14644 11406
rect 14028 11284 14084 11294
rect 14028 11190 14084 11228
rect 14588 11282 14644 11340
rect 14812 11396 14868 11406
rect 14812 11394 15092 11396
rect 14812 11342 14814 11394
rect 14866 11342 15092 11394
rect 14812 11340 15092 11342
rect 14812 11330 14868 11340
rect 14588 11230 14590 11282
rect 14642 11230 14644 11282
rect 14588 11218 14644 11230
rect 13132 10834 13412 10836
rect 13132 10782 13134 10834
rect 13186 10782 13412 10834
rect 13132 10780 13412 10782
rect 13132 10770 13188 10780
rect 12796 9998 12798 10050
rect 12850 9998 12852 10050
rect 12796 9986 12852 9998
rect 13356 9828 13412 10780
rect 14028 10724 14084 10734
rect 14028 10722 14308 10724
rect 14028 10670 14030 10722
rect 14082 10670 14308 10722
rect 14028 10668 14308 10670
rect 14028 10658 14084 10668
rect 14252 9938 14308 10668
rect 14252 9886 14254 9938
rect 14306 9886 14308 9938
rect 14252 9874 14308 9886
rect 14364 10610 14420 10622
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 13468 9828 13524 9838
rect 13356 9826 13524 9828
rect 13356 9774 13470 9826
rect 13522 9774 13524 9826
rect 13356 9772 13524 9774
rect 13132 9154 13188 9166
rect 13132 9102 13134 9154
rect 13186 9102 13188 9154
rect 12460 8878 12462 8930
rect 12514 8878 12516 8930
rect 12460 8866 12516 8878
rect 12908 9042 12964 9054
rect 12908 8990 12910 9042
rect 12962 8990 12964 9042
rect 12908 8708 12964 8990
rect 12908 8642 12964 8652
rect 12236 8082 12292 8092
rect 12572 8260 12628 8270
rect 12572 7474 12628 8204
rect 13132 8260 13188 9102
rect 13132 8194 13188 8204
rect 12572 7422 12574 7474
rect 12626 7422 12628 7474
rect 12572 7410 12628 7422
rect 12684 8036 12740 8046
rect 13468 8036 13524 9772
rect 14364 9266 14420 10558
rect 14364 9214 14366 9266
rect 14418 9214 14420 9266
rect 14364 9202 14420 9214
rect 15036 9940 15092 11340
rect 15036 9268 15092 9884
rect 15148 9380 15204 9390
rect 15148 9268 15204 9324
rect 15036 9212 15204 9268
rect 13692 8930 13748 8942
rect 13692 8878 13694 8930
rect 13746 8878 13748 8930
rect 13692 8708 13748 8878
rect 13692 8642 13748 8652
rect 14700 8820 14756 8830
rect 14700 8428 14756 8764
rect 13580 8372 13636 8382
rect 13580 8278 13636 8316
rect 14364 8372 14756 8428
rect 12684 8034 13524 8036
rect 12684 7982 12686 8034
rect 12738 7982 13524 8034
rect 12684 7980 13524 7982
rect 11452 7252 11508 7262
rect 9660 6748 10052 6804
rect 9996 6692 10052 6748
rect 10108 6692 10164 6702
rect 9996 6636 10108 6692
rect 10108 6598 10164 6636
rect 10780 6580 10836 6590
rect 10780 6578 11284 6580
rect 10780 6526 10782 6578
rect 10834 6526 11284 6578
rect 10780 6524 11284 6526
rect 10780 6514 10836 6524
rect 11228 6130 11284 6524
rect 11228 6078 11230 6130
rect 11282 6078 11284 6130
rect 11228 6066 11284 6078
rect 11452 5906 11508 7196
rect 12236 7252 12292 7262
rect 12236 7158 12292 7196
rect 11452 5854 11454 5906
rect 11506 5854 11508 5906
rect 11452 5842 11508 5854
rect 12236 6692 12292 6702
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 12236 4564 12292 6636
rect 12684 6692 12740 7980
rect 12908 7588 12964 7598
rect 12908 6802 12964 7532
rect 13356 7588 13412 7598
rect 13356 7494 13412 7532
rect 13244 7476 13300 7486
rect 13244 7382 13300 7420
rect 12908 6750 12910 6802
rect 12962 6750 12964 6802
rect 12908 6738 12964 6750
rect 13468 6692 13524 7980
rect 13916 8258 13972 8270
rect 13916 8206 13918 8258
rect 13970 8206 13972 8258
rect 13916 7588 13972 8206
rect 14140 8148 14196 8158
rect 14140 8054 14196 8092
rect 13916 7522 13972 7532
rect 14364 6914 14420 8372
rect 14700 8146 14756 8158
rect 14700 8094 14702 8146
rect 14754 8094 14756 8146
rect 14700 7588 14756 8094
rect 14700 7522 14756 7532
rect 14812 8148 14868 8158
rect 14364 6862 14366 6914
rect 14418 6862 14420 6914
rect 14364 6850 14420 6862
rect 14812 7476 14868 8092
rect 13580 6692 13636 6702
rect 13468 6690 13636 6692
rect 13468 6638 13582 6690
rect 13634 6638 13636 6690
rect 13468 6636 13636 6638
rect 12684 6626 12740 6636
rect 13580 6626 13636 6636
rect 14812 6690 14868 7420
rect 15260 6804 15316 15092
rect 15372 14644 15428 14654
rect 15596 14644 15652 15148
rect 15372 14642 15652 14644
rect 15372 14590 15374 14642
rect 15426 14590 15652 14642
rect 15372 14588 15652 14590
rect 15372 14578 15428 14588
rect 15708 14420 15764 15596
rect 15932 14756 15988 15820
rect 16492 15876 16548 15886
rect 16380 15652 16436 15662
rect 16380 15148 16436 15596
rect 15932 14690 15988 14700
rect 16268 15092 16436 15148
rect 15932 14420 15988 14430
rect 16268 14420 16324 15092
rect 16492 14530 16548 15820
rect 17052 15652 17108 23660
rect 17164 17668 17220 26852
rect 17836 24610 17892 29036
rect 18284 28866 18340 29484
rect 18396 29314 18452 30156
rect 18396 29262 18398 29314
rect 18450 29262 18452 29314
rect 18396 29250 18452 29262
rect 18620 30210 18676 30222
rect 18620 30158 18622 30210
rect 18674 30158 18676 30210
rect 18620 29092 18676 30158
rect 19516 30212 19572 30222
rect 19516 30118 19572 30156
rect 18620 29026 18676 29036
rect 18844 29764 18900 29774
rect 18844 29538 18900 29708
rect 19404 29652 19460 29662
rect 19628 29652 19684 34862
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19740 34018 19796 34030
rect 19740 33966 19742 34018
rect 19794 33966 19796 34018
rect 19740 33124 19796 33966
rect 20300 34018 20356 34030
rect 20300 33966 20302 34018
rect 20354 33966 20356 34018
rect 20076 33458 20132 33470
rect 20076 33406 20078 33458
rect 20130 33406 20132 33458
rect 20076 33124 20132 33406
rect 20076 33068 20244 33124
rect 19740 33058 19796 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32788 20244 33068
rect 20076 32732 20244 32788
rect 20076 31778 20132 32732
rect 20300 32004 20356 33966
rect 20412 34020 20468 38612
rect 20636 37156 20692 39676
rect 20748 39730 20804 41468
rect 20748 39678 20750 39730
rect 20802 39678 20804 39730
rect 20748 38836 20804 39678
rect 20748 38164 20804 38780
rect 20748 38098 20804 38108
rect 20860 39844 20916 39854
rect 20860 39060 20916 39788
rect 21084 39508 21140 41694
rect 21196 40402 21252 43708
rect 21308 43708 21364 45838
rect 21420 45892 21476 46620
rect 21532 45892 21588 45902
rect 21420 45890 21588 45892
rect 21420 45838 21534 45890
rect 21586 45838 21588 45890
rect 21420 45836 21588 45838
rect 21532 45106 21588 45836
rect 21644 45892 21700 47182
rect 21756 46676 21812 47404
rect 21756 46582 21812 46620
rect 21756 46004 21812 46014
rect 21756 45910 21812 45948
rect 21644 45826 21700 45836
rect 21532 45054 21534 45106
rect 21586 45054 21588 45106
rect 21532 45042 21588 45054
rect 21308 43652 21700 43708
rect 21532 43540 21588 43550
rect 21196 40350 21198 40402
rect 21250 40350 21252 40402
rect 21196 40338 21252 40350
rect 21308 43538 21588 43540
rect 21308 43486 21534 43538
rect 21586 43486 21588 43538
rect 21308 43484 21588 43486
rect 21308 42756 21364 43484
rect 21532 43474 21588 43484
rect 21308 41188 21364 42700
rect 21532 41972 21588 41982
rect 21532 41878 21588 41916
rect 21644 41636 21700 43652
rect 21868 43538 21924 48972
rect 22988 48962 23044 48974
rect 23212 48916 23268 48926
rect 23212 48822 23268 48860
rect 22764 48804 22820 48814
rect 22652 48802 22820 48804
rect 22652 48750 22766 48802
rect 22818 48750 22820 48802
rect 22652 48748 22820 48750
rect 22652 48356 22708 48748
rect 22764 48738 22820 48748
rect 23324 48466 23380 50540
rect 23548 50530 23604 50540
rect 23660 50428 23716 51212
rect 23772 51266 23828 51996
rect 23996 51986 24052 51996
rect 24108 51716 24164 52220
rect 23772 51214 23774 51266
rect 23826 51214 23828 51266
rect 23772 51202 23828 51214
rect 23996 51660 24164 51716
rect 24220 51938 24276 51950
rect 24220 51886 24222 51938
rect 24274 51886 24276 51938
rect 23884 50596 23940 50606
rect 23884 50482 23940 50540
rect 23884 50430 23886 50482
rect 23938 50430 23940 50482
rect 23660 50372 23828 50428
rect 23884 50418 23940 50430
rect 23660 49924 23716 49934
rect 23660 49810 23716 49868
rect 23660 49758 23662 49810
rect 23714 49758 23716 49810
rect 23660 48914 23716 49758
rect 23660 48862 23662 48914
rect 23714 48862 23716 48914
rect 23660 48850 23716 48862
rect 23772 48580 23828 50372
rect 23996 49138 24052 51660
rect 24108 50594 24164 50606
rect 24108 50542 24110 50594
rect 24162 50542 24164 50594
rect 24108 50484 24164 50542
rect 24108 50418 24164 50428
rect 24220 50034 24276 51886
rect 24332 51828 24388 52892
rect 24444 52444 24724 52500
rect 24444 52162 24500 52444
rect 24556 52276 24612 52286
rect 24668 52276 24724 52444
rect 25004 52276 25060 52286
rect 25116 52276 25172 54908
rect 25228 54404 25284 55246
rect 25788 55298 25844 55310
rect 25788 55246 25790 55298
rect 25842 55246 25844 55298
rect 25228 54338 25284 54348
rect 25340 54402 25396 54414
rect 25340 54350 25342 54402
rect 25394 54350 25396 54402
rect 25340 53060 25396 54350
rect 25788 54404 25844 55246
rect 26012 54740 26068 59200
rect 26908 56308 26964 59200
rect 27356 56642 27412 59200
rect 27356 56590 27358 56642
rect 27410 56590 27412 56642
rect 27356 56578 27412 56590
rect 27020 56308 27076 56318
rect 26908 56306 27076 56308
rect 26908 56254 27022 56306
rect 27074 56254 27076 56306
rect 26908 56252 27076 56254
rect 27020 56242 27076 56252
rect 26124 56082 26180 56094
rect 26124 56030 26126 56082
rect 26178 56030 26180 56082
rect 26124 54964 26180 56030
rect 27804 56082 27860 56094
rect 27804 56030 27806 56082
rect 27858 56030 27860 56082
rect 27804 55972 27860 56030
rect 27804 55906 27860 55916
rect 26124 54898 26180 54908
rect 26460 55186 26516 55198
rect 26460 55134 26462 55186
rect 26514 55134 26516 55186
rect 26236 54740 26292 54750
rect 26012 54738 26292 54740
rect 26012 54686 26238 54738
rect 26290 54686 26292 54738
rect 26012 54684 26292 54686
rect 26236 54674 26292 54684
rect 25788 54310 25844 54348
rect 26460 54068 26516 55134
rect 28252 54740 28308 59200
rect 28364 56642 28420 56654
rect 28364 56590 28366 56642
rect 28418 56590 28420 56642
rect 28364 56306 28420 56590
rect 28364 56254 28366 56306
rect 28418 56254 28420 56306
rect 28364 56242 28420 56254
rect 28700 56308 28756 59200
rect 29484 56642 29540 56654
rect 29484 56590 29486 56642
rect 29538 56590 29540 56642
rect 28924 56308 28980 56318
rect 28700 56306 28980 56308
rect 28700 56254 28926 56306
rect 28978 56254 28980 56306
rect 28700 56252 28980 56254
rect 28924 56242 28980 56252
rect 29484 56306 29540 56590
rect 29484 56254 29486 56306
rect 29538 56254 29540 56306
rect 29484 56242 29540 56254
rect 29596 56308 29652 59200
rect 30044 56642 30100 59200
rect 30044 56590 30046 56642
rect 30098 56590 30100 56642
rect 30044 56578 30100 56590
rect 29596 56242 29652 56252
rect 30716 56308 30772 56318
rect 30268 56082 30324 56094
rect 30268 56030 30270 56082
rect 30322 56030 30324 56082
rect 29932 55972 29988 55982
rect 29988 55916 30212 55972
rect 29932 55878 29988 55916
rect 28252 54674 28308 54684
rect 28588 55410 28644 55422
rect 28588 55358 28590 55410
rect 28642 55358 28644 55410
rect 28588 54514 28644 55358
rect 28588 54462 28590 54514
rect 28642 54462 28644 54514
rect 28588 54450 28644 54462
rect 29148 55298 29204 55310
rect 29148 55246 29150 55298
rect 29202 55246 29204 55298
rect 29148 54404 29204 55246
rect 29932 55188 29988 55198
rect 29932 55186 30100 55188
rect 29932 55134 29934 55186
rect 29986 55134 30100 55186
rect 29932 55132 30100 55134
rect 29932 55122 29988 55132
rect 29260 54740 29316 54750
rect 29260 54646 29316 54684
rect 30044 54738 30100 55132
rect 30044 54686 30046 54738
rect 30098 54686 30100 54738
rect 30044 54674 30100 54686
rect 29148 54338 29204 54348
rect 29708 54404 29764 54414
rect 29708 54310 29764 54348
rect 26460 54002 26516 54012
rect 28252 53956 28308 53966
rect 25452 53060 25508 53070
rect 26012 53060 26068 53070
rect 25396 53058 26068 53060
rect 25396 53006 25454 53058
rect 25506 53006 26014 53058
rect 26066 53006 26068 53058
rect 25396 53004 26068 53006
rect 24668 52274 25172 52276
rect 24668 52222 25006 52274
rect 25058 52222 25172 52274
rect 24668 52220 25172 52222
rect 25228 52722 25284 52734
rect 25228 52670 25230 52722
rect 25282 52670 25284 52722
rect 25228 52276 25284 52670
rect 24556 52182 24612 52220
rect 25004 52210 25060 52220
rect 25228 52210 25284 52220
rect 24444 52110 24446 52162
rect 24498 52110 24500 52162
rect 24444 52098 24500 52110
rect 24556 51938 24612 51950
rect 24556 51886 24558 51938
rect 24610 51886 24612 51938
rect 24556 51828 24612 51886
rect 24332 51772 24612 51828
rect 24332 51492 24388 51772
rect 24332 50706 24388 51436
rect 25228 51716 25284 51726
rect 24332 50654 24334 50706
rect 24386 50654 24388 50706
rect 24332 50642 24388 50654
rect 24444 51268 24500 51278
rect 25228 51268 25284 51660
rect 24444 50370 24500 51212
rect 25004 51266 25284 51268
rect 25004 51214 25230 51266
rect 25282 51214 25284 51266
rect 25004 51212 25284 51214
rect 25004 50706 25060 51212
rect 25228 51202 25284 51212
rect 25004 50654 25006 50706
rect 25058 50654 25060 50706
rect 25004 50642 25060 50654
rect 24556 50484 24612 50494
rect 24892 50484 24948 50494
rect 24556 50482 24948 50484
rect 24556 50430 24558 50482
rect 24610 50430 24894 50482
rect 24946 50430 24948 50482
rect 24556 50428 24948 50430
rect 25340 50428 25396 53004
rect 25452 52994 25508 53004
rect 26012 52994 26068 53004
rect 28252 53058 28308 53900
rect 28252 53006 28254 53058
rect 28306 53006 28308 53058
rect 28252 52994 28308 53006
rect 27580 52946 27636 52958
rect 27580 52894 27582 52946
rect 27634 52894 27636 52946
rect 25564 52724 25620 52734
rect 25564 52630 25620 52668
rect 27132 52724 27188 52734
rect 25564 52500 25620 52510
rect 24556 50418 24612 50428
rect 24892 50418 24948 50428
rect 24444 50318 24446 50370
rect 24498 50318 24500 50370
rect 24444 50306 24500 50318
rect 25228 50372 25396 50428
rect 25452 50484 25508 50522
rect 25452 50418 25508 50428
rect 24220 49982 24222 50034
rect 24274 49982 24276 50034
rect 24220 49970 24276 49982
rect 24108 49810 24164 49822
rect 24332 49812 24388 49822
rect 24108 49758 24110 49810
rect 24162 49758 24164 49810
rect 24108 49252 24164 49758
rect 24108 49186 24164 49196
rect 24220 49810 24388 49812
rect 24220 49758 24334 49810
rect 24386 49758 24388 49810
rect 24220 49756 24388 49758
rect 23996 49086 23998 49138
rect 24050 49086 24052 49138
rect 23996 49074 24052 49086
rect 24108 49028 24164 49038
rect 24220 49028 24276 49756
rect 24332 49746 24388 49756
rect 24108 49026 24276 49028
rect 24108 48974 24110 49026
rect 24162 48974 24276 49026
rect 24108 48972 24276 48974
rect 23884 48916 23940 48926
rect 23884 48822 23940 48860
rect 23772 48524 23940 48580
rect 23324 48414 23326 48466
rect 23378 48414 23380 48466
rect 23324 48402 23380 48414
rect 22540 47348 22596 47358
rect 22540 47254 22596 47292
rect 22652 47068 22708 48300
rect 23772 48356 23828 48366
rect 23772 48262 23828 48300
rect 23100 48244 23156 48254
rect 22764 48132 22820 48142
rect 22764 48038 22820 48076
rect 22988 48020 23044 48030
rect 22988 47926 23044 47964
rect 22764 47796 22820 47806
rect 22764 47458 22820 47740
rect 22764 47406 22766 47458
rect 22818 47406 22820 47458
rect 22764 47394 22820 47406
rect 23100 47458 23156 48188
rect 23660 48242 23716 48254
rect 23660 48190 23662 48242
rect 23714 48190 23716 48242
rect 23100 47406 23102 47458
rect 23154 47406 23156 47458
rect 23100 47394 23156 47406
rect 23548 48132 23604 48142
rect 22764 47236 22820 47246
rect 22764 47234 23380 47236
rect 22764 47182 22766 47234
rect 22818 47182 23380 47234
rect 22764 47180 23380 47182
rect 22764 47170 22820 47180
rect 22652 47012 22820 47068
rect 22092 46676 22148 46686
rect 21980 46674 22148 46676
rect 21980 46622 22094 46674
rect 22146 46622 22148 46674
rect 21980 46620 22148 46622
rect 21980 46116 22036 46620
rect 22092 46610 22148 46620
rect 22316 46674 22372 46686
rect 22316 46622 22318 46674
rect 22370 46622 22372 46674
rect 22316 46564 22372 46622
rect 22316 46116 22372 46508
rect 21980 46050 22036 46060
rect 22092 46060 22372 46116
rect 22092 44996 22148 46060
rect 22540 45890 22596 45902
rect 22540 45838 22542 45890
rect 22594 45838 22596 45890
rect 22204 45668 22260 45678
rect 22204 45666 22372 45668
rect 22204 45614 22206 45666
rect 22258 45614 22372 45666
rect 22204 45612 22372 45614
rect 22204 45602 22260 45612
rect 22092 44930 22148 44940
rect 22316 44322 22372 45612
rect 22540 45556 22596 45838
rect 22316 44270 22318 44322
rect 22370 44270 22372 44322
rect 22316 44258 22372 44270
rect 22428 45500 22596 45556
rect 22204 44210 22260 44222
rect 22204 44158 22206 44210
rect 22258 44158 22260 44210
rect 22204 43764 22260 44158
rect 22428 43988 22484 45500
rect 22204 43698 22260 43708
rect 22316 43932 22484 43988
rect 21868 43486 21870 43538
rect 21922 43486 21924 43538
rect 21868 43428 21924 43486
rect 21868 43362 21924 43372
rect 21868 43092 21924 43102
rect 21924 43036 22036 43092
rect 21868 43026 21924 43036
rect 21980 42084 22036 43036
rect 22316 42980 22372 43932
rect 22428 43764 22484 43774
rect 22428 43670 22484 43708
rect 22204 42924 22372 42980
rect 22652 42980 22708 42990
rect 22764 42980 22820 47012
rect 23100 46900 23156 46910
rect 22652 42978 22820 42980
rect 22652 42926 22654 42978
rect 22706 42926 22820 42978
rect 22652 42924 22820 42926
rect 22876 46786 22932 46798
rect 22876 46734 22878 46786
rect 22930 46734 22932 46786
rect 21644 41570 21700 41580
rect 21868 41972 21924 41982
rect 21308 40180 21364 41132
rect 21420 41186 21476 41198
rect 21420 41134 21422 41186
rect 21474 41134 21476 41186
rect 21420 40292 21476 41134
rect 21756 41076 21812 41086
rect 21644 40964 21700 40974
rect 21644 40870 21700 40908
rect 21420 40226 21476 40236
rect 21644 40402 21700 40414
rect 21644 40350 21646 40402
rect 21698 40350 21700 40402
rect 21084 39442 21140 39452
rect 21196 40124 21364 40180
rect 20860 37378 20916 39004
rect 20860 37326 20862 37378
rect 20914 37326 20916 37378
rect 20860 37314 20916 37326
rect 21196 37266 21252 40124
rect 21308 39732 21364 39742
rect 21644 39732 21700 40350
rect 21756 40290 21812 41020
rect 21868 40628 21924 41916
rect 21980 41970 22036 42028
rect 21980 41918 21982 41970
rect 22034 41918 22036 41970
rect 21980 41906 22036 41918
rect 22092 42642 22148 42654
rect 22092 42590 22094 42642
rect 22146 42590 22148 42642
rect 22092 42532 22148 42590
rect 21980 41188 22036 41198
rect 21980 40740 22036 41132
rect 22092 40964 22148 42476
rect 22204 42420 22260 42924
rect 22652 42914 22708 42924
rect 22204 41524 22260 42364
rect 22316 42754 22372 42766
rect 22316 42702 22318 42754
rect 22370 42702 22372 42754
rect 22316 42196 22372 42702
rect 22316 42130 22372 42140
rect 22876 42084 22932 46734
rect 23100 46786 23156 46844
rect 23100 46734 23102 46786
rect 23154 46734 23156 46786
rect 23100 46722 23156 46734
rect 23212 46228 23268 46238
rect 22988 45892 23044 45902
rect 22988 45556 23044 45836
rect 22988 45490 23044 45500
rect 23212 45106 23268 46172
rect 23324 46116 23380 47180
rect 23436 47124 23492 47134
rect 23436 46674 23492 47068
rect 23548 46788 23604 48076
rect 23660 48020 23716 48190
rect 23660 46900 23716 47964
rect 23884 47460 23940 48524
rect 23996 48468 24052 48478
rect 24108 48468 24164 48972
rect 25004 48916 25060 48926
rect 23996 48466 24164 48468
rect 23996 48414 23998 48466
rect 24050 48414 24164 48466
rect 23996 48412 24164 48414
rect 24668 48468 24724 48478
rect 23996 48402 24052 48412
rect 24668 48354 24724 48412
rect 24668 48302 24670 48354
rect 24722 48302 24724 48354
rect 24668 48290 24724 48302
rect 24332 48244 24388 48254
rect 24332 48150 24388 48188
rect 24332 48018 24388 48030
rect 24332 47966 24334 48018
rect 24386 47966 24388 48018
rect 24332 47684 24388 47966
rect 24332 47618 24388 47628
rect 23884 47404 24948 47460
rect 24108 47236 24164 47246
rect 24108 47142 24164 47180
rect 24556 47236 24612 47246
rect 24556 47142 24612 47180
rect 24108 46900 24164 46910
rect 23660 46844 23828 46900
rect 23548 46732 23716 46788
rect 23436 46622 23438 46674
rect 23490 46622 23492 46674
rect 23436 46564 23492 46622
rect 23436 46508 23604 46564
rect 23436 46116 23492 46126
rect 23324 46114 23492 46116
rect 23324 46062 23438 46114
rect 23490 46062 23492 46114
rect 23324 46060 23492 46062
rect 23436 46050 23492 46060
rect 23548 45892 23604 46508
rect 23660 46114 23716 46732
rect 23660 46062 23662 46114
rect 23714 46062 23716 46114
rect 23660 46050 23716 46062
rect 23212 45054 23214 45106
rect 23266 45054 23268 45106
rect 23212 45042 23268 45054
rect 23436 45836 23604 45892
rect 23436 45108 23492 45836
rect 23436 45042 23492 45052
rect 23548 44994 23604 45006
rect 23548 44942 23550 44994
rect 23602 44942 23604 44994
rect 23324 44324 23380 44334
rect 23548 44324 23604 44942
rect 23324 44322 23604 44324
rect 23324 44270 23326 44322
rect 23378 44270 23604 44322
rect 23324 44268 23604 44270
rect 23324 44258 23380 44268
rect 23212 44210 23268 44222
rect 23212 44158 23214 44210
rect 23266 44158 23268 44210
rect 22988 44100 23044 44110
rect 22988 42754 23044 44044
rect 23212 43708 23268 44158
rect 23660 43764 23716 43774
rect 23772 43764 23828 46844
rect 24108 46806 24164 46844
rect 24668 46562 24724 46574
rect 24668 46510 24670 46562
rect 24722 46510 24724 46562
rect 24220 46004 24276 46014
rect 24220 45910 24276 45948
rect 23884 45890 23940 45902
rect 23884 45838 23886 45890
rect 23938 45838 23940 45890
rect 23884 45556 23940 45838
rect 23884 45490 23940 45500
rect 24108 45666 24164 45678
rect 24108 45614 24110 45666
rect 24162 45614 24164 45666
rect 23996 45220 24052 45230
rect 23884 45108 23940 45118
rect 23884 45014 23940 45052
rect 23660 43762 23828 43764
rect 23660 43710 23662 43762
rect 23714 43710 23828 43762
rect 23660 43708 23828 43710
rect 23212 43652 23380 43708
rect 23660 43698 23716 43708
rect 23212 43540 23268 43550
rect 23212 43446 23268 43484
rect 22988 42702 22990 42754
rect 23042 42702 23044 42754
rect 22988 42690 23044 42702
rect 23212 42644 23268 42654
rect 23212 42550 23268 42588
rect 22428 42082 22932 42084
rect 22428 42030 22878 42082
rect 22930 42030 22932 42082
rect 22428 42028 22932 42030
rect 22204 41468 22372 41524
rect 22204 41300 22260 41310
rect 22204 41186 22260 41244
rect 22204 41134 22206 41186
rect 22258 41134 22260 41186
rect 22204 41122 22260 41134
rect 22316 40964 22372 41468
rect 22428 41074 22484 42028
rect 22876 42018 22932 42028
rect 22988 41970 23044 41982
rect 22988 41918 22990 41970
rect 23042 41918 23044 41970
rect 22540 41524 22596 41534
rect 22540 41410 22596 41468
rect 22540 41358 22542 41410
rect 22594 41358 22596 41410
rect 22540 41346 22596 41358
rect 22652 41412 22708 41422
rect 22652 41186 22708 41356
rect 22988 41300 23044 41918
rect 23100 41972 23156 41982
rect 23324 41972 23380 43652
rect 23548 43540 23604 43550
rect 23548 43538 23716 43540
rect 23548 43486 23550 43538
rect 23602 43486 23716 43538
rect 23548 43484 23716 43486
rect 23548 43474 23604 43484
rect 23548 42980 23604 42990
rect 23548 42866 23604 42924
rect 23548 42814 23550 42866
rect 23602 42814 23604 42866
rect 23548 42802 23604 42814
rect 23100 41970 23268 41972
rect 23100 41918 23102 41970
rect 23154 41918 23268 41970
rect 23100 41916 23268 41918
rect 23100 41906 23156 41916
rect 23100 41300 23156 41310
rect 22988 41244 23100 41300
rect 23100 41234 23156 41244
rect 22652 41134 22654 41186
rect 22706 41134 22708 41186
rect 22652 41122 22708 41134
rect 22876 41188 22932 41198
rect 22932 41132 23044 41188
rect 22876 41122 22932 41132
rect 22428 41022 22430 41074
rect 22482 41022 22484 41074
rect 22428 41010 22484 41022
rect 22988 41076 23044 41132
rect 23212 41076 23268 41916
rect 23324 41906 23380 41916
rect 23660 42644 23716 43484
rect 23772 43538 23828 43550
rect 23772 43486 23774 43538
rect 23826 43486 23828 43538
rect 23772 42868 23828 43486
rect 23772 42802 23828 42812
rect 23548 41748 23604 41758
rect 23548 41654 23604 41692
rect 23660 41636 23716 42588
rect 23660 41570 23716 41580
rect 23324 41300 23380 41310
rect 23324 41206 23380 41244
rect 22988 41074 23268 41076
rect 22988 41022 22990 41074
rect 23042 41022 23268 41074
rect 22988 41020 23268 41022
rect 23436 41076 23492 41086
rect 23996 41076 24052 45164
rect 24108 42980 24164 45614
rect 24332 45666 24388 45678
rect 24332 45614 24334 45666
rect 24386 45614 24388 45666
rect 24332 45332 24388 45614
rect 24668 45444 24724 46510
rect 24668 45378 24724 45388
rect 24388 45276 24612 45332
rect 24332 45266 24388 45276
rect 24220 44324 24276 44334
rect 24220 43652 24276 44268
rect 24556 43652 24612 45276
rect 24668 43652 24724 43662
rect 24556 43650 24724 43652
rect 24556 43598 24670 43650
rect 24722 43598 24724 43650
rect 24556 43596 24724 43598
rect 24220 43558 24276 43596
rect 24444 43538 24500 43550
rect 24444 43486 24446 43538
rect 24498 43486 24500 43538
rect 24220 43428 24276 43438
rect 24444 43428 24500 43486
rect 24276 43372 24500 43428
rect 24220 43362 24276 43372
rect 24108 41300 24164 42924
rect 24444 42644 24500 43372
rect 24556 43428 24612 43438
rect 24556 43334 24612 43372
rect 24668 43092 24724 43596
rect 24668 43026 24724 43036
rect 24892 42756 24948 47404
rect 25004 46676 25060 48860
rect 25116 48804 25172 48814
rect 25116 47570 25172 48748
rect 25116 47518 25118 47570
rect 25170 47518 25172 47570
rect 25116 46900 25172 47518
rect 25116 46834 25172 46844
rect 25004 46620 25172 46676
rect 25004 46452 25060 46462
rect 25004 45890 25060 46396
rect 25004 45838 25006 45890
rect 25058 45838 25060 45890
rect 25004 45826 25060 45838
rect 25004 44436 25060 44446
rect 25004 44342 25060 44380
rect 25116 43204 25172 46620
rect 25116 43138 25172 43148
rect 24444 42578 24500 42588
rect 24556 42754 24948 42756
rect 24556 42702 24894 42754
rect 24946 42702 24948 42754
rect 24556 42700 24948 42702
rect 24164 41244 24276 41300
rect 24108 41234 24164 41244
rect 23996 41020 24164 41076
rect 22988 41010 23044 41020
rect 23436 40982 23492 41020
rect 22092 40898 22148 40908
rect 22204 40908 22372 40964
rect 22876 40962 22932 40974
rect 22876 40910 22878 40962
rect 22930 40910 22932 40962
rect 21980 40684 22148 40740
rect 21868 40572 22036 40628
rect 21756 40238 21758 40290
rect 21810 40238 21812 40290
rect 21756 40226 21812 40238
rect 21868 40402 21924 40414
rect 21868 40350 21870 40402
rect 21922 40350 21924 40402
rect 21868 39844 21924 40350
rect 21868 39778 21924 39788
rect 21364 39676 21700 39732
rect 21308 39618 21364 39676
rect 21308 39566 21310 39618
rect 21362 39566 21364 39618
rect 21308 39554 21364 39566
rect 21868 39618 21924 39630
rect 21868 39566 21870 39618
rect 21922 39566 21924 39618
rect 21868 39508 21924 39566
rect 21868 39442 21924 39452
rect 21756 38836 21812 38846
rect 21756 38742 21812 38780
rect 21980 38668 22036 40572
rect 22092 40626 22148 40684
rect 22092 40574 22094 40626
rect 22146 40574 22148 40626
rect 22092 40562 22148 40574
rect 21756 38612 21812 38622
rect 21756 38164 21812 38556
rect 21756 38070 21812 38108
rect 21868 38612 22036 38668
rect 22092 40292 22148 40302
rect 21420 37938 21476 37950
rect 21420 37886 21422 37938
rect 21474 37886 21476 37938
rect 21196 37214 21198 37266
rect 21250 37214 21252 37266
rect 21196 37202 21252 37214
rect 21308 37826 21364 37838
rect 21308 37774 21310 37826
rect 21362 37774 21364 37826
rect 21308 37268 21364 37774
rect 21420 37380 21476 37886
rect 21420 37314 21476 37324
rect 21868 37826 21924 38612
rect 21868 37774 21870 37826
rect 21922 37774 21924 37826
rect 21308 37202 21364 37212
rect 21644 37268 21700 37278
rect 21644 37174 21700 37212
rect 20636 37090 20692 37100
rect 20636 36820 20692 36830
rect 20524 36484 20580 36494
rect 20524 36390 20580 36428
rect 20636 35140 20692 36764
rect 21756 36484 21812 36494
rect 20748 36370 20804 36382
rect 20748 36318 20750 36370
rect 20802 36318 20804 36370
rect 20748 35924 20804 36318
rect 21308 36148 21364 36158
rect 21364 36092 21588 36148
rect 21308 36082 21364 36092
rect 20748 35364 20804 35868
rect 21532 35810 21588 36092
rect 21532 35758 21534 35810
rect 21586 35758 21588 35810
rect 21532 35746 21588 35758
rect 20748 35298 20804 35308
rect 20636 35084 21476 35140
rect 20412 33954 20468 33964
rect 20524 35026 20580 35038
rect 20524 34974 20526 35026
rect 20578 34974 20580 35026
rect 20412 33796 20468 33806
rect 20412 33124 20468 33740
rect 20524 33684 20580 34974
rect 20636 34914 20692 35084
rect 20636 34862 20638 34914
rect 20690 34862 20692 34914
rect 20636 34850 20692 34862
rect 21308 34916 21364 34926
rect 21308 34822 21364 34860
rect 21420 34914 21476 35084
rect 21420 34862 21422 34914
rect 21474 34862 21476 34914
rect 21420 34850 21476 34862
rect 20748 34804 20804 34814
rect 20748 34710 20804 34748
rect 21756 34692 21812 36428
rect 21868 34804 21924 37774
rect 22092 37378 22148 40236
rect 22092 37326 22094 37378
rect 22146 37326 22148 37378
rect 22092 36594 22148 37326
rect 22092 36542 22094 36594
rect 22146 36542 22148 36594
rect 22092 36530 22148 36542
rect 21980 36482 22036 36494
rect 21980 36430 21982 36482
rect 22034 36430 22036 36482
rect 21980 36036 22036 36430
rect 22204 36484 22260 40908
rect 22428 40628 22484 40638
rect 22316 40516 22372 40526
rect 22316 40422 22372 40460
rect 22428 40514 22484 40572
rect 22428 40462 22430 40514
rect 22482 40462 22484 40514
rect 22428 40450 22484 40462
rect 22876 40404 22932 40910
rect 22428 39620 22484 39630
rect 22428 39526 22484 39564
rect 22540 39394 22596 39406
rect 22764 39396 22820 39406
rect 22540 39342 22542 39394
rect 22594 39342 22596 39394
rect 22540 39284 22596 39342
rect 22540 39218 22596 39228
rect 22652 39394 22820 39396
rect 22652 39342 22766 39394
rect 22818 39342 22820 39394
rect 22652 39340 22820 39342
rect 22540 38948 22596 38958
rect 22652 38948 22708 39340
rect 22764 39330 22820 39340
rect 22540 38946 22708 38948
rect 22540 38894 22542 38946
rect 22594 38894 22708 38946
rect 22540 38892 22708 38894
rect 22540 38882 22596 38892
rect 22540 37828 22596 37838
rect 22540 37826 22708 37828
rect 22540 37774 22542 37826
rect 22594 37774 22708 37826
rect 22540 37772 22708 37774
rect 22540 37762 22596 37772
rect 22428 37268 22484 37278
rect 22428 37174 22484 37212
rect 22652 37042 22708 37772
rect 22652 36990 22654 37042
rect 22706 36990 22708 37042
rect 22652 36978 22708 36990
rect 22540 36596 22596 36606
rect 22540 36594 22820 36596
rect 22540 36542 22542 36594
rect 22594 36542 22820 36594
rect 22540 36540 22820 36542
rect 22540 36530 22596 36540
rect 22204 36418 22260 36428
rect 22428 36482 22484 36494
rect 22428 36430 22430 36482
rect 22482 36430 22484 36482
rect 22428 36372 22484 36430
rect 22428 36306 22484 36316
rect 22204 36036 22260 36046
rect 21980 35980 22204 36036
rect 22204 35970 22260 35980
rect 22316 35698 22372 35710
rect 22316 35646 22318 35698
rect 22370 35646 22372 35698
rect 21980 34804 22036 34814
rect 21868 34748 21980 34804
rect 21980 34710 22036 34748
rect 21756 34636 21924 34692
rect 21868 34354 21924 34636
rect 21868 34302 21870 34354
rect 21922 34302 21924 34354
rect 21868 34290 21924 34302
rect 20860 34132 20916 34142
rect 20860 34038 20916 34076
rect 21308 34020 21364 34030
rect 21308 33926 21364 33964
rect 20524 33618 20580 33628
rect 21756 33684 21812 33694
rect 20524 33124 20580 33134
rect 20412 33068 20524 33124
rect 20524 33030 20580 33068
rect 21420 33122 21476 33134
rect 21420 33070 21422 33122
rect 21474 33070 21476 33122
rect 21420 33012 21476 33070
rect 21420 32946 21476 32956
rect 21084 32450 21140 32462
rect 21084 32398 21086 32450
rect 21138 32398 21140 32450
rect 20300 31948 20580 32004
rect 20076 31726 20078 31778
rect 20130 31726 20132 31778
rect 20076 31556 20132 31726
rect 20524 31780 20580 31948
rect 20524 31686 20580 31724
rect 20412 31668 20468 31678
rect 20412 31574 20468 31612
rect 20748 31668 20804 31678
rect 20748 31574 20804 31612
rect 20076 31490 20132 31500
rect 20300 31554 20356 31566
rect 20300 31502 20302 31554
rect 20354 31502 20356 31554
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20300 31220 20356 31502
rect 21084 31220 21140 32398
rect 21532 32450 21588 32462
rect 21532 32398 21534 32450
rect 21586 32398 21588 32450
rect 21308 31778 21364 31790
rect 21308 31726 21310 31778
rect 21362 31726 21364 31778
rect 21308 31556 21364 31726
rect 21308 31490 21364 31500
rect 21532 31666 21588 32398
rect 21532 31614 21534 31666
rect 21586 31614 21588 31666
rect 20300 31164 21476 31220
rect 21420 30994 21476 31164
rect 21420 30942 21422 30994
rect 21474 30942 21476 30994
rect 21308 30884 21364 30894
rect 21308 30434 21364 30828
rect 21308 30382 21310 30434
rect 21362 30382 21364 30434
rect 21308 30370 21364 30382
rect 20076 30098 20132 30110
rect 20076 30046 20078 30098
rect 20130 30046 20132 30098
rect 20076 29988 20132 30046
rect 21420 30098 21476 30942
rect 21532 30212 21588 31614
rect 21644 30212 21700 30222
rect 21532 30156 21644 30212
rect 21644 30118 21700 30156
rect 21420 30046 21422 30098
rect 21474 30046 21476 30098
rect 21420 30034 21476 30046
rect 20076 29922 20132 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 21756 29652 21812 33628
rect 22316 33348 22372 35646
rect 22428 35476 22484 35486
rect 22764 35476 22820 36540
rect 22876 36036 22932 40348
rect 23884 40180 23940 40190
rect 23548 39732 23604 39742
rect 23548 39638 23604 39676
rect 22988 39396 23044 39406
rect 22988 38724 23044 39340
rect 23100 39394 23156 39406
rect 23100 39342 23102 39394
rect 23154 39342 23156 39394
rect 23100 39284 23156 39342
rect 23100 39218 23156 39228
rect 22988 38658 23044 38668
rect 22988 38388 23044 38398
rect 22988 38164 23044 38332
rect 22988 38070 23044 38108
rect 22988 37492 23044 37502
rect 23044 37436 23268 37492
rect 22988 37398 23044 37436
rect 22876 35970 22932 35980
rect 22988 37042 23044 37054
rect 22988 36990 22990 37042
rect 23042 36990 23044 37042
rect 22988 35924 23044 36990
rect 23212 36484 23268 37436
rect 23324 37266 23380 37278
rect 23884 37268 23940 40124
rect 23996 39394 24052 39406
rect 23996 39342 23998 39394
rect 24050 39342 24052 39394
rect 23996 38500 24052 39342
rect 23996 38434 24052 38444
rect 23996 37940 24052 37950
rect 23996 37846 24052 37884
rect 24108 37492 24164 41020
rect 24108 37426 24164 37436
rect 23324 37214 23326 37266
rect 23378 37214 23380 37266
rect 23324 37044 23380 37214
rect 23548 37266 23940 37268
rect 23548 37214 23886 37266
rect 23938 37214 23940 37266
rect 23548 37212 23940 37214
rect 23548 37156 23604 37212
rect 23884 37202 23940 37212
rect 23324 36978 23380 36988
rect 23436 37100 23604 37156
rect 23324 36484 23380 36494
rect 23212 36482 23380 36484
rect 23212 36430 23326 36482
rect 23378 36430 23380 36482
rect 23212 36428 23380 36430
rect 23324 36418 23380 36428
rect 23100 36260 23156 36270
rect 23100 36258 23380 36260
rect 23100 36206 23102 36258
rect 23154 36206 23380 36258
rect 23100 36204 23380 36206
rect 23100 36194 23156 36204
rect 22988 35858 23044 35868
rect 23212 36036 23268 36046
rect 23212 35698 23268 35980
rect 23212 35646 23214 35698
rect 23266 35646 23268 35698
rect 23212 35634 23268 35646
rect 23324 35700 23380 36204
rect 23324 35634 23380 35644
rect 23436 35586 23492 37100
rect 23996 36484 24052 36494
rect 24220 36484 24276 41244
rect 24556 40514 24612 42700
rect 24892 42690 24948 42700
rect 25004 40964 25060 40974
rect 24668 40628 24724 40638
rect 24668 40534 24724 40572
rect 24556 40462 24558 40514
rect 24610 40462 24612 40514
rect 24556 39284 24612 40462
rect 25004 39618 25060 40908
rect 25228 40740 25284 50372
rect 25340 48802 25396 48814
rect 25340 48750 25342 48802
rect 25394 48750 25396 48802
rect 25340 47684 25396 48750
rect 25340 47618 25396 47628
rect 25452 48018 25508 48030
rect 25452 47966 25454 48018
rect 25506 47966 25508 48018
rect 25340 47346 25396 47358
rect 25340 47294 25342 47346
rect 25394 47294 25396 47346
rect 25340 46676 25396 47294
rect 25452 47124 25508 47966
rect 25452 47058 25508 47068
rect 25340 45890 25396 46620
rect 25564 46116 25620 52444
rect 27132 52274 27188 52668
rect 27132 52222 27134 52274
rect 27186 52222 27188 52274
rect 27132 52210 27188 52222
rect 27580 52164 27636 52894
rect 27916 52164 27972 52174
rect 27580 52162 27972 52164
rect 27580 52110 27918 52162
rect 27970 52110 27972 52162
rect 27580 52108 27972 52110
rect 27356 51268 27412 51278
rect 27356 51174 27412 51212
rect 26908 50484 26964 50494
rect 25676 48802 25732 48814
rect 25676 48750 25678 48802
rect 25730 48750 25732 48802
rect 25676 48580 25732 48750
rect 26796 48802 26852 48814
rect 26796 48750 26798 48802
rect 26850 48750 26852 48802
rect 26796 48692 26852 48750
rect 26796 48626 26852 48636
rect 25676 48514 25732 48524
rect 25788 48468 25844 48478
rect 25788 48242 25844 48412
rect 26460 48468 26516 48478
rect 25788 48190 25790 48242
rect 25842 48190 25844 48242
rect 25788 48178 25844 48190
rect 26012 48244 26068 48254
rect 26012 48150 26068 48188
rect 26460 48242 26516 48412
rect 26460 48190 26462 48242
rect 26514 48190 26516 48242
rect 26460 48178 26516 48190
rect 26684 48354 26740 48366
rect 26684 48302 26686 48354
rect 26738 48302 26740 48354
rect 26684 48132 26740 48302
rect 26684 48066 26740 48076
rect 25676 47684 25732 47722
rect 25676 47618 25732 47628
rect 26684 47684 26740 47694
rect 25676 47458 25732 47470
rect 25676 47406 25678 47458
rect 25730 47406 25732 47458
rect 25676 47236 25732 47406
rect 25676 46674 25732 47180
rect 25676 46622 25678 46674
rect 25730 46622 25732 46674
rect 25676 46610 25732 46622
rect 26012 47348 26068 47358
rect 25340 45838 25342 45890
rect 25394 45838 25396 45890
rect 25340 45826 25396 45838
rect 25452 46060 25620 46116
rect 25452 44436 25508 46060
rect 25900 45778 25956 45790
rect 25900 45726 25902 45778
rect 25954 45726 25956 45778
rect 25564 45666 25620 45678
rect 25564 45614 25566 45666
rect 25618 45614 25620 45666
rect 25564 45556 25620 45614
rect 25676 45668 25732 45678
rect 25900 45668 25956 45726
rect 25676 45666 25844 45668
rect 25676 45614 25678 45666
rect 25730 45614 25844 45666
rect 25676 45612 25844 45614
rect 25676 45602 25732 45612
rect 25564 45490 25620 45500
rect 25340 44380 25508 44436
rect 25676 45444 25732 45454
rect 25676 45330 25732 45388
rect 25676 45278 25678 45330
rect 25730 45278 25732 45330
rect 25340 43650 25396 44380
rect 25676 44324 25732 45278
rect 25788 45220 25844 45612
rect 25900 45602 25956 45612
rect 26012 45666 26068 47292
rect 26236 47234 26292 47246
rect 26236 47182 26238 47234
rect 26290 47182 26292 47234
rect 26236 47124 26292 47182
rect 26236 47058 26292 47068
rect 26572 47234 26628 47246
rect 26572 47182 26574 47234
rect 26626 47182 26628 47234
rect 26236 46564 26292 46574
rect 26236 46562 26404 46564
rect 26236 46510 26238 46562
rect 26290 46510 26404 46562
rect 26236 46508 26404 46510
rect 26236 46498 26292 46508
rect 26236 45668 26292 45678
rect 26012 45614 26014 45666
rect 26066 45614 26068 45666
rect 26012 45556 26068 45614
rect 25900 45220 25956 45230
rect 25788 45218 25956 45220
rect 25788 45166 25902 45218
rect 25954 45166 25956 45218
rect 25788 45164 25956 45166
rect 25900 45154 25956 45164
rect 26012 44996 26068 45500
rect 25900 44940 26068 44996
rect 26124 45666 26292 45668
rect 26124 45614 26238 45666
rect 26290 45614 26292 45666
rect 26124 45612 26292 45614
rect 25340 43598 25342 43650
rect 25394 43598 25396 43650
rect 25340 43316 25396 43598
rect 25452 44322 25732 44324
rect 25452 44270 25678 44322
rect 25730 44270 25732 44322
rect 25452 44268 25732 44270
rect 25452 43652 25508 44268
rect 25676 44258 25732 44268
rect 25788 44434 25844 44446
rect 25788 44382 25790 44434
rect 25842 44382 25844 44434
rect 25788 43876 25844 44382
rect 25900 44100 25956 44940
rect 26012 44212 26068 44222
rect 26124 44212 26180 45612
rect 26236 45602 26292 45612
rect 26348 45332 26404 46508
rect 26572 46116 26628 47182
rect 26572 46050 26628 46060
rect 26684 46786 26740 47628
rect 26684 46734 26686 46786
rect 26738 46734 26740 46786
rect 26684 45892 26740 46734
rect 26796 46452 26852 46462
rect 26796 46358 26852 46396
rect 26908 46340 26964 50428
rect 27692 49810 27748 52108
rect 27916 51604 27972 52108
rect 28364 51938 28420 51950
rect 28364 51886 28366 51938
rect 28418 51886 28420 51938
rect 28364 51604 28420 51886
rect 28588 51604 28644 51614
rect 27916 51548 28588 51604
rect 28140 51378 28196 51548
rect 28140 51326 28142 51378
rect 28194 51326 28196 51378
rect 28140 51314 28196 51326
rect 28364 50706 28420 51548
rect 28588 51378 28644 51548
rect 28588 51326 28590 51378
rect 28642 51326 28644 51378
rect 28588 51314 28644 51326
rect 28364 50654 28366 50706
rect 28418 50654 28420 50706
rect 28364 50642 28420 50654
rect 29260 51266 29316 51278
rect 29260 51214 29262 51266
rect 29314 51214 29316 51266
rect 29260 50428 29316 51214
rect 29260 50372 29652 50428
rect 27692 49758 27694 49810
rect 27746 49758 27748 49810
rect 27692 49746 27748 49758
rect 28364 49700 28420 49710
rect 28140 49698 28420 49700
rect 28140 49646 28366 49698
rect 28418 49646 28420 49698
rect 28140 49644 28420 49646
rect 27580 49140 27636 49150
rect 27468 48914 27524 48926
rect 27468 48862 27470 48914
rect 27522 48862 27524 48914
rect 27244 48802 27300 48814
rect 27244 48750 27246 48802
rect 27298 48750 27300 48802
rect 27244 47796 27300 48750
rect 27244 47730 27300 47740
rect 27356 48692 27412 48702
rect 27356 48242 27412 48636
rect 27356 48190 27358 48242
rect 27410 48190 27412 48242
rect 27244 47572 27300 47582
rect 27356 47572 27412 48190
rect 27300 47516 27412 47572
rect 27244 47478 27300 47516
rect 27468 47348 27524 48862
rect 27580 48914 27636 49084
rect 28140 49138 28196 49644
rect 28364 49634 28420 49644
rect 28140 49086 28142 49138
rect 28194 49086 28196 49138
rect 28140 49074 28196 49086
rect 28476 49140 28532 49150
rect 27804 49028 27860 49038
rect 27804 48934 27860 48972
rect 27580 48862 27582 48914
rect 27634 48862 27636 48914
rect 27580 48850 27636 48862
rect 28028 48802 28084 48814
rect 28028 48750 28030 48802
rect 28082 48750 28084 48802
rect 27580 48580 27636 48590
rect 27580 48466 27636 48524
rect 27580 48414 27582 48466
rect 27634 48414 27636 48466
rect 27580 48402 27636 48414
rect 27692 48468 27748 48478
rect 28028 48468 28084 48750
rect 28252 48804 28308 48814
rect 28252 48710 28308 48748
rect 27692 48466 28084 48468
rect 27692 48414 27694 48466
rect 27746 48414 28084 48466
rect 27692 48412 28084 48414
rect 27692 48402 27748 48412
rect 27804 48242 27860 48254
rect 27804 48190 27806 48242
rect 27858 48190 27860 48242
rect 27804 47684 27860 48190
rect 27916 48242 27972 48254
rect 27916 48190 27918 48242
rect 27970 48190 27972 48242
rect 27916 48132 27972 48190
rect 28364 48132 28420 48142
rect 27916 48066 27972 48076
rect 28252 48076 28364 48132
rect 27804 47628 28084 47684
rect 27692 47460 27748 47470
rect 27916 47460 27972 47470
rect 27692 47366 27748 47404
rect 27804 47458 27972 47460
rect 27804 47406 27918 47458
rect 27970 47406 27972 47458
rect 27804 47404 27972 47406
rect 27580 47348 27636 47358
rect 27468 47346 27636 47348
rect 27468 47294 27582 47346
rect 27634 47294 27636 47346
rect 27468 47292 27636 47294
rect 27580 47236 27636 47292
rect 27692 47236 27748 47246
rect 27580 47180 27692 47236
rect 27692 47170 27748 47180
rect 27804 47012 27860 47404
rect 27916 47394 27972 47404
rect 28028 47348 28084 47628
rect 28028 47282 28084 47292
rect 28140 47234 28196 47246
rect 28140 47182 28142 47234
rect 28194 47182 28196 47234
rect 28140 47012 28196 47182
rect 27356 46956 27860 47012
rect 27916 46956 28196 47012
rect 27132 46900 27188 46910
rect 27132 46674 27188 46844
rect 27356 46898 27412 46956
rect 27356 46846 27358 46898
rect 27410 46846 27412 46898
rect 27356 46834 27412 46846
rect 27132 46622 27134 46674
rect 27186 46622 27188 46674
rect 27132 46610 27188 46622
rect 27468 46450 27524 46462
rect 27468 46398 27470 46450
rect 27522 46398 27524 46450
rect 26908 46284 27188 46340
rect 27020 46116 27076 46126
rect 26796 45892 26852 45902
rect 26348 45266 26404 45276
rect 26572 45890 26852 45892
rect 26572 45838 26798 45890
rect 26850 45838 26852 45890
rect 26572 45836 26852 45838
rect 26348 44996 26404 45006
rect 26012 44210 26180 44212
rect 26012 44158 26014 44210
rect 26066 44158 26180 44210
rect 26012 44156 26180 44158
rect 26236 44994 26404 44996
rect 26236 44942 26350 44994
rect 26402 44942 26404 44994
rect 26236 44940 26404 44942
rect 26012 44146 26068 44156
rect 25900 44034 25956 44044
rect 26236 43988 26292 44940
rect 26348 44930 26404 44940
rect 26460 44324 26516 44334
rect 26236 43922 26292 43932
rect 26348 44322 26516 44324
rect 26348 44270 26462 44322
rect 26514 44270 26516 44322
rect 26348 44268 26516 44270
rect 25788 43810 25844 43820
rect 26348 43708 26404 44268
rect 26460 44258 26516 44268
rect 26572 44100 26628 45836
rect 26796 45826 26852 45836
rect 26908 45666 26964 45678
rect 26908 45614 26910 45666
rect 26962 45614 26964 45666
rect 26796 45220 26852 45230
rect 26684 45108 26740 45118
rect 26684 45014 26740 45052
rect 26684 44212 26740 44222
rect 26796 44212 26852 45164
rect 26908 44660 26964 45614
rect 27020 45666 27076 46060
rect 27132 45892 27188 46284
rect 27468 46116 27524 46398
rect 27468 46050 27524 46060
rect 27580 46452 27636 46462
rect 27132 45836 27524 45892
rect 27020 45614 27022 45666
rect 27074 45614 27076 45666
rect 27020 45444 27076 45614
rect 27244 45668 27300 45678
rect 27468 45668 27524 45836
rect 27580 45890 27636 46396
rect 27580 45838 27582 45890
rect 27634 45838 27636 45890
rect 27580 45826 27636 45838
rect 27692 45780 27748 45790
rect 27468 45612 27636 45668
rect 27244 45574 27300 45612
rect 27020 45378 27076 45388
rect 27244 45106 27300 45118
rect 27244 45054 27246 45106
rect 27298 45054 27300 45106
rect 27244 44884 27300 45054
rect 27244 44818 27300 44828
rect 27468 45106 27524 45118
rect 27468 45054 27470 45106
rect 27522 45054 27524 45106
rect 26908 44594 26964 44604
rect 27356 44324 27412 44334
rect 27356 44230 27412 44268
rect 26684 44210 26852 44212
rect 26684 44158 26686 44210
rect 26738 44158 26852 44210
rect 26684 44156 26852 44158
rect 26684 44146 26740 44156
rect 25452 43586 25508 43596
rect 25564 43652 26404 43708
rect 26460 44044 26628 44100
rect 25340 43250 25396 43260
rect 25564 42866 25620 43652
rect 25676 43540 25732 43550
rect 25676 43538 26068 43540
rect 25676 43486 25678 43538
rect 25730 43486 26068 43538
rect 25676 43484 26068 43486
rect 25676 43474 25732 43484
rect 25788 43316 25844 43326
rect 25844 43260 25956 43316
rect 25788 43250 25844 43260
rect 25564 42814 25566 42866
rect 25618 42814 25620 42866
rect 25452 42756 25508 42766
rect 25452 42662 25508 42700
rect 25340 41970 25396 41982
rect 25340 41918 25342 41970
rect 25394 41918 25396 41970
rect 25340 41410 25396 41918
rect 25340 41358 25342 41410
rect 25394 41358 25396 41410
rect 25340 41346 25396 41358
rect 25452 41188 25508 41198
rect 25564 41188 25620 42814
rect 25452 41186 25620 41188
rect 25452 41134 25454 41186
rect 25506 41134 25620 41186
rect 25452 41132 25620 41134
rect 25676 43204 25732 43214
rect 25452 41122 25508 41132
rect 25340 40964 25396 40974
rect 25340 40870 25396 40908
rect 25228 40684 25620 40740
rect 25228 40404 25284 40414
rect 25116 40402 25284 40404
rect 25116 40350 25230 40402
rect 25282 40350 25284 40402
rect 25116 40348 25284 40350
rect 25116 39730 25172 40348
rect 25228 40338 25284 40348
rect 25116 39678 25118 39730
rect 25170 39678 25172 39730
rect 25116 39666 25172 39678
rect 25340 39620 25396 39630
rect 25004 39566 25006 39618
rect 25058 39566 25060 39618
rect 24556 39228 24836 39284
rect 24668 38722 24724 38734
rect 24668 38670 24670 38722
rect 24722 38670 24724 38722
rect 24668 38500 24724 38670
rect 24668 38434 24724 38444
rect 24780 38050 24836 39228
rect 24780 37998 24782 38050
rect 24834 37998 24836 38050
rect 24780 37986 24836 37998
rect 24332 37938 24388 37950
rect 24332 37886 24334 37938
rect 24386 37886 24388 37938
rect 24332 37378 24388 37886
rect 25004 37492 25060 39566
rect 25228 39564 25340 39620
rect 25228 39058 25284 39564
rect 25340 39526 25396 39564
rect 25228 39006 25230 39058
rect 25282 39006 25284 39058
rect 25228 38994 25284 39006
rect 25452 38834 25508 38846
rect 25452 38782 25454 38834
rect 25506 38782 25508 38834
rect 25452 38668 25508 38782
rect 25340 38612 25508 38668
rect 25228 38052 25284 38062
rect 25340 38052 25396 38612
rect 25452 38546 25508 38556
rect 25228 38050 25396 38052
rect 25228 37998 25230 38050
rect 25282 37998 25396 38050
rect 25228 37996 25396 37998
rect 25228 37986 25284 37996
rect 24332 37326 24334 37378
rect 24386 37326 24388 37378
rect 24332 37314 24388 37326
rect 24556 37436 25060 37492
rect 23996 36482 24276 36484
rect 23996 36430 23998 36482
rect 24050 36430 24276 36482
rect 23996 36428 24276 36430
rect 24444 37154 24500 37166
rect 24444 37102 24446 37154
rect 24498 37102 24500 37154
rect 23996 36418 24052 36428
rect 23436 35534 23438 35586
rect 23490 35534 23492 35586
rect 23436 35522 23492 35534
rect 23772 36258 23828 36270
rect 23772 36206 23774 36258
rect 23826 36206 23828 36258
rect 22764 35420 23156 35476
rect 22428 35026 22484 35420
rect 22428 34974 22430 35026
rect 22482 34974 22484 35026
rect 22428 34962 22484 34974
rect 22764 35252 22820 35262
rect 22764 34356 22820 35196
rect 22540 34354 22820 34356
rect 22540 34302 22766 34354
rect 22818 34302 22820 34354
rect 22540 34300 22820 34302
rect 22316 33292 22484 33348
rect 22204 33234 22260 33246
rect 22204 33182 22206 33234
rect 22258 33182 22260 33234
rect 21868 33122 21924 33134
rect 21868 33070 21870 33122
rect 21922 33070 21924 33122
rect 21868 33012 21924 33070
rect 21868 32946 21924 32956
rect 21868 31892 21924 31902
rect 22204 31892 22260 33182
rect 22316 33122 22372 33134
rect 22316 33070 22318 33122
rect 22370 33070 22372 33122
rect 22316 32564 22372 33070
rect 22428 33012 22484 33292
rect 22540 33346 22596 34300
rect 22764 34290 22820 34300
rect 22540 33294 22542 33346
rect 22594 33294 22596 33346
rect 22540 33282 22596 33294
rect 22428 32946 22484 32956
rect 22316 32498 22372 32508
rect 21924 31836 22260 31892
rect 21868 31798 21924 31836
rect 22540 31780 22596 31790
rect 21980 31668 22036 31678
rect 21980 30770 22036 31612
rect 22540 31666 22596 31724
rect 22540 31614 22542 31666
rect 22594 31614 22596 31666
rect 22540 31602 22596 31614
rect 22652 31778 22708 31790
rect 22652 31726 22654 31778
rect 22706 31726 22708 31778
rect 21980 30718 21982 30770
rect 22034 30718 22036 30770
rect 21868 30436 21924 30446
rect 21868 30210 21924 30380
rect 21868 30158 21870 30210
rect 21922 30158 21924 30210
rect 21868 30146 21924 30158
rect 19404 29650 20132 29652
rect 19404 29598 19406 29650
rect 19458 29598 20132 29650
rect 19404 29596 20132 29598
rect 19404 29586 19460 29596
rect 18844 29486 18846 29538
rect 18898 29486 18900 29538
rect 18284 28814 18286 28866
rect 18338 28814 18340 28866
rect 18284 28802 18340 28814
rect 18396 28532 18452 28542
rect 18396 28438 18452 28476
rect 18620 27748 18676 27758
rect 18620 26180 18676 27692
rect 18508 26178 18676 26180
rect 18508 26126 18622 26178
rect 18674 26126 18676 26178
rect 18508 26124 18676 26126
rect 18396 25620 18452 25630
rect 18284 25618 18452 25620
rect 18284 25566 18398 25618
rect 18450 25566 18452 25618
rect 18284 25564 18452 25566
rect 17836 24558 17838 24610
rect 17890 24558 17892 24610
rect 17276 23938 17332 23950
rect 17276 23886 17278 23938
rect 17330 23886 17332 23938
rect 17276 23828 17332 23886
rect 17276 23762 17332 23772
rect 17500 23938 17556 23950
rect 17500 23886 17502 23938
rect 17554 23886 17556 23938
rect 17500 23380 17556 23886
rect 17500 23314 17556 23324
rect 17612 23826 17668 23838
rect 17612 23774 17614 23826
rect 17666 23774 17668 23826
rect 17612 22372 17668 23774
rect 17724 23828 17780 23838
rect 17724 23378 17780 23772
rect 17724 23326 17726 23378
rect 17778 23326 17780 23378
rect 17724 23314 17780 23326
rect 17836 23826 17892 24558
rect 18172 25284 18228 25294
rect 18284 25284 18340 25564
rect 18396 25554 18452 25564
rect 18228 25228 18340 25284
rect 18172 24722 18228 25228
rect 18396 25172 18452 25182
rect 18508 25172 18564 26124
rect 18620 26114 18676 26124
rect 18732 25284 18788 25294
rect 18732 25190 18788 25228
rect 18452 25116 18564 25172
rect 18396 25106 18452 25116
rect 18844 24948 18900 29486
rect 19180 28532 19236 28542
rect 19068 28420 19124 28430
rect 19068 28082 19124 28364
rect 19068 28030 19070 28082
rect 19122 28030 19124 28082
rect 19068 28018 19124 28030
rect 18956 27636 19012 27646
rect 18956 27542 19012 27580
rect 19180 27188 19236 28476
rect 19628 28418 19684 28430
rect 19628 28366 19630 28418
rect 19682 28366 19684 28418
rect 19628 27860 19684 28366
rect 20076 28420 20132 29596
rect 21756 29586 21812 29596
rect 21868 29764 21924 29774
rect 21308 28868 21364 28878
rect 20412 28866 21364 28868
rect 20412 28814 21310 28866
rect 21362 28814 21364 28866
rect 20412 28812 21364 28814
rect 20076 28364 20244 28420
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19740 27860 19796 27870
rect 19628 27858 19796 27860
rect 19628 27806 19742 27858
rect 19794 27806 19796 27858
rect 19628 27804 19796 27806
rect 19740 27748 19796 27804
rect 19740 27682 19796 27692
rect 19292 27636 19348 27646
rect 19292 27634 19684 27636
rect 19292 27582 19294 27634
rect 19346 27582 19684 27634
rect 19292 27580 19684 27582
rect 19292 27570 19348 27580
rect 19292 27188 19348 27198
rect 19180 27186 19348 27188
rect 19180 27134 19294 27186
rect 19346 27134 19348 27186
rect 19180 27132 19348 27134
rect 19180 26908 19236 27132
rect 19292 27122 19348 27132
rect 19628 27186 19684 27580
rect 19628 27134 19630 27186
rect 19682 27134 19684 27186
rect 19628 27122 19684 27134
rect 18620 24892 18900 24948
rect 18956 26852 19236 26908
rect 20076 27074 20132 27086
rect 20076 27022 20078 27074
rect 20130 27022 20132 27074
rect 20076 26852 20132 27022
rect 20188 26908 20244 28364
rect 20412 27970 20468 28812
rect 21308 28802 21364 28812
rect 21644 28644 21700 28654
rect 21868 28644 21924 29708
rect 21980 29314 22036 30718
rect 22092 30882 22148 30894
rect 22092 30830 22094 30882
rect 22146 30830 22148 30882
rect 22092 30210 22148 30830
rect 22428 30436 22484 30446
rect 22652 30436 22708 31726
rect 22988 30994 23044 31006
rect 22988 30942 22990 30994
rect 23042 30942 23044 30994
rect 22764 30436 22820 30446
rect 22652 30434 22820 30436
rect 22652 30382 22766 30434
rect 22818 30382 22820 30434
rect 22652 30380 22820 30382
rect 22092 30158 22094 30210
rect 22146 30158 22148 30210
rect 22092 30146 22148 30158
rect 22316 30212 22372 30222
rect 22316 30098 22372 30156
rect 22428 30210 22484 30380
rect 22764 30370 22820 30380
rect 22428 30158 22430 30210
rect 22482 30158 22484 30210
rect 22428 30146 22484 30158
rect 22988 30212 23044 30942
rect 22988 30146 23044 30156
rect 22316 30046 22318 30098
rect 22370 30046 22372 30098
rect 22316 30034 22372 30046
rect 22876 30100 22932 30110
rect 22876 30006 22932 30044
rect 21980 29262 21982 29314
rect 22034 29262 22036 29314
rect 21980 29250 22036 29262
rect 22092 29426 22148 29438
rect 22092 29374 22094 29426
rect 22146 29374 22148 29426
rect 20412 27918 20414 27970
rect 20466 27918 20468 27970
rect 20412 27906 20468 27918
rect 21308 28642 21700 28644
rect 21308 28590 21646 28642
rect 21698 28590 21700 28642
rect 21308 28588 21700 28590
rect 21308 27186 21364 28588
rect 21644 28578 21700 28588
rect 21756 28588 21924 28644
rect 21420 28420 21476 28430
rect 21420 28326 21476 28364
rect 21756 28420 21812 28588
rect 21308 27134 21310 27186
rect 21362 27134 21364 27186
rect 21308 27122 21364 27134
rect 21532 27524 21588 27534
rect 20524 27076 20580 27086
rect 20524 26982 20580 27020
rect 20188 26852 20356 26908
rect 18956 26290 19012 26852
rect 20076 26786 20132 26796
rect 18956 26238 18958 26290
rect 19010 26238 19012 26290
rect 18508 24836 18564 24846
rect 18508 24742 18564 24780
rect 18172 24670 18174 24722
rect 18226 24670 18228 24722
rect 17836 23774 17838 23826
rect 17890 23774 17892 23826
rect 17724 22372 17780 22382
rect 17612 22316 17724 22372
rect 17724 22306 17780 22316
rect 17836 22260 17892 23774
rect 17948 24500 18004 24510
rect 17948 23378 18004 24444
rect 18172 23940 18228 24670
rect 18172 23884 18452 23940
rect 18284 23714 18340 23726
rect 18284 23662 18286 23714
rect 18338 23662 18340 23714
rect 18284 23492 18340 23662
rect 18284 23426 18340 23436
rect 17948 23326 17950 23378
rect 18002 23326 18004 23378
rect 17948 23314 18004 23326
rect 18172 23380 18228 23390
rect 18060 23156 18116 23166
rect 18060 23062 18116 23100
rect 17948 22260 18004 22270
rect 17836 22204 17948 22260
rect 17948 22194 18004 22204
rect 18172 22258 18228 23324
rect 18172 22206 18174 22258
rect 18226 22206 18228 22258
rect 18172 22194 18228 22206
rect 18284 22036 18340 22046
rect 17500 21476 17556 21486
rect 17500 21382 17556 21420
rect 17612 21252 17668 21262
rect 17388 21028 17444 21038
rect 17388 20802 17444 20972
rect 17388 20750 17390 20802
rect 17442 20750 17444 20802
rect 17388 20738 17444 20750
rect 17612 20578 17668 21196
rect 18060 21252 18116 21262
rect 17612 20526 17614 20578
rect 17666 20526 17668 20578
rect 17612 20244 17668 20526
rect 17612 20178 17668 20188
rect 17836 21028 17892 21038
rect 17836 20242 17892 20972
rect 17836 20190 17838 20242
rect 17890 20190 17892 20242
rect 17836 20178 17892 20190
rect 18060 20802 18116 21196
rect 18060 20750 18062 20802
rect 18114 20750 18116 20802
rect 17388 20020 17444 20030
rect 17388 18450 17444 19964
rect 17612 19796 17668 19806
rect 17388 18398 17390 18450
rect 17442 18398 17444 18450
rect 17388 18386 17444 18398
rect 17500 19234 17556 19246
rect 17500 19182 17502 19234
rect 17554 19182 17556 19234
rect 17500 18452 17556 19182
rect 17500 18386 17556 18396
rect 17500 18226 17556 18238
rect 17500 18174 17502 18226
rect 17554 18174 17556 18226
rect 17500 17892 17556 18174
rect 17612 17892 17668 19740
rect 17948 18340 18004 18350
rect 17948 18246 18004 18284
rect 17500 17836 17780 17892
rect 17612 17668 17668 17678
rect 17164 17666 17668 17668
rect 17164 17614 17166 17666
rect 17218 17614 17614 17666
rect 17666 17614 17668 17666
rect 17164 17612 17668 17614
rect 17164 17602 17220 17612
rect 17612 17602 17668 17612
rect 17388 16994 17444 17006
rect 17388 16942 17390 16994
rect 17442 16942 17444 16994
rect 17388 16548 17444 16942
rect 17388 16482 17444 16492
rect 17500 16996 17556 17006
rect 17724 16996 17780 17836
rect 18060 17780 18116 20750
rect 18060 17714 18116 17724
rect 18172 21028 18228 21038
rect 18172 18116 18228 20972
rect 18284 20578 18340 21980
rect 18396 21700 18452 23884
rect 18620 23380 18676 24892
rect 18956 24500 19012 26238
rect 19516 26740 19572 26750
rect 19516 26290 19572 26684
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19516 26238 19518 26290
rect 19570 26238 19572 26290
rect 19516 26180 19572 26238
rect 19292 25394 19348 25406
rect 19292 25342 19294 25394
rect 19346 25342 19348 25394
rect 19068 25172 19124 25182
rect 19068 24722 19124 25116
rect 19068 24670 19070 24722
rect 19122 24670 19124 24722
rect 19068 24658 19124 24670
rect 18956 24434 19012 24444
rect 19180 24610 19236 24622
rect 19180 24558 19182 24610
rect 19234 24558 19236 24610
rect 18732 23828 18788 23838
rect 18732 23734 18788 23772
rect 18620 23154 18676 23324
rect 18620 23102 18622 23154
rect 18674 23102 18676 23154
rect 18620 23090 18676 23102
rect 18508 22932 18564 22942
rect 18508 22930 18676 22932
rect 18508 22878 18510 22930
rect 18562 22878 18676 22930
rect 18508 22876 18676 22878
rect 18508 22866 18564 22876
rect 18396 21634 18452 21644
rect 18508 21474 18564 21486
rect 18508 21422 18510 21474
rect 18562 21422 18564 21474
rect 18508 21252 18564 21422
rect 18508 21186 18564 21196
rect 18620 20804 18676 22876
rect 19180 22482 19236 24558
rect 19292 23716 19348 25342
rect 19292 23650 19348 23660
rect 19516 23380 19572 26124
rect 20300 25506 20356 26852
rect 20636 26516 20692 26526
rect 20300 25454 20302 25506
rect 20354 25454 20356 25506
rect 19852 25394 19908 25406
rect 19852 25342 19854 25394
rect 19906 25342 19908 25394
rect 19852 25284 19908 25342
rect 20300 25396 20356 25454
rect 20300 25330 20356 25340
rect 20412 26290 20468 26302
rect 20412 26238 20414 26290
rect 20466 26238 20468 26290
rect 19964 25284 20020 25294
rect 19852 25228 19964 25284
rect 19964 25218 20020 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19628 24722 19684 24734
rect 19628 24670 19630 24722
rect 19682 24670 19684 24722
rect 19628 24500 19684 24670
rect 19628 24434 19684 24444
rect 20076 24610 20132 24622
rect 20076 24558 20078 24610
rect 20130 24558 20132 24610
rect 19516 23314 19572 23324
rect 19628 23938 19684 23950
rect 19628 23886 19630 23938
rect 19682 23886 19684 23938
rect 19628 23828 19684 23886
rect 19180 22430 19182 22482
rect 19234 22430 19236 22482
rect 18732 22372 18788 22382
rect 18732 22278 18788 22316
rect 19068 22260 19124 22270
rect 19068 22166 19124 22204
rect 18956 21140 19012 21150
rect 18956 21026 19012 21084
rect 18956 20974 18958 21026
rect 19010 20974 19012 21026
rect 18956 20962 19012 20974
rect 18284 20526 18286 20578
rect 18338 20526 18340 20578
rect 18284 20468 18340 20526
rect 18284 20402 18340 20412
rect 18508 20748 18676 20804
rect 18284 20130 18340 20142
rect 18284 20078 18286 20130
rect 18338 20078 18340 20130
rect 18284 19346 18340 20078
rect 18284 19294 18286 19346
rect 18338 19294 18340 19346
rect 18284 19282 18340 19294
rect 17948 17498 18004 17510
rect 17948 17446 17950 17498
rect 18002 17446 18004 17498
rect 17836 16996 17892 17006
rect 17724 16940 17836 16996
rect 17500 16100 17556 16940
rect 17836 16930 17892 16940
rect 17612 16882 17668 16894
rect 17612 16830 17614 16882
rect 17666 16830 17668 16882
rect 17612 16772 17668 16830
rect 17948 16884 18004 17446
rect 17948 16818 18004 16828
rect 17612 16706 17668 16716
rect 18172 16772 18228 18060
rect 18284 18452 18340 18462
rect 18284 16882 18340 18396
rect 18396 18340 18452 18350
rect 18396 18246 18452 18284
rect 18284 16830 18286 16882
rect 18338 16830 18340 16882
rect 18284 16818 18340 16830
rect 18172 16706 18228 16716
rect 18284 16324 18340 16334
rect 18060 16100 18116 16110
rect 17500 16098 17892 16100
rect 17500 16046 17502 16098
rect 17554 16046 17892 16098
rect 17500 16044 17892 16046
rect 17500 16034 17556 16044
rect 17164 15876 17220 15886
rect 17164 15782 17220 15820
rect 17052 15586 17108 15596
rect 17836 15538 17892 16044
rect 18060 16006 18116 16044
rect 18284 15986 18340 16268
rect 18284 15934 18286 15986
rect 18338 15934 18340 15986
rect 18284 15922 18340 15934
rect 17836 15486 17838 15538
rect 17890 15486 17892 15538
rect 17836 15474 17892 15486
rect 16492 14478 16494 14530
rect 16546 14478 16548 14530
rect 16492 14466 16548 14478
rect 16828 14756 16884 14766
rect 16828 14530 16884 14700
rect 16828 14478 16830 14530
rect 16882 14478 16884 14530
rect 16828 14466 16884 14478
rect 18508 14532 18564 20748
rect 19180 20690 19236 22430
rect 19516 23156 19572 23166
rect 19516 21812 19572 23100
rect 19628 22930 19684 23772
rect 19964 23938 20020 23950
rect 19964 23886 19966 23938
rect 20018 23886 20020 23938
rect 19964 23716 20020 23886
rect 20076 23716 20132 24558
rect 20300 23716 20356 23726
rect 20412 23716 20468 26238
rect 20636 24946 20692 26460
rect 21084 26404 21140 26414
rect 20748 26402 21140 26404
rect 20748 26350 21086 26402
rect 21138 26350 21140 26402
rect 20748 26348 21140 26350
rect 20748 26290 20804 26348
rect 21084 26338 21140 26348
rect 20748 26238 20750 26290
rect 20802 26238 20804 26290
rect 20748 26226 20804 26238
rect 21196 26290 21252 26302
rect 21196 26238 21198 26290
rect 21250 26238 21252 26290
rect 20860 26178 20916 26190
rect 20860 26126 20862 26178
rect 20914 26126 20916 26178
rect 20748 25394 20804 25406
rect 20748 25342 20750 25394
rect 20802 25342 20804 25394
rect 20748 25284 20804 25342
rect 20748 25218 20804 25228
rect 20636 24894 20638 24946
rect 20690 24894 20692 24946
rect 20636 24882 20692 24894
rect 20748 24948 20804 24958
rect 20748 24854 20804 24892
rect 20860 24834 20916 26126
rect 21196 26180 21252 26238
rect 21196 26114 21252 26124
rect 21420 26290 21476 26302
rect 21420 26238 21422 26290
rect 21474 26238 21476 26290
rect 20860 24782 20862 24834
rect 20914 24782 20916 24834
rect 20860 24770 20916 24782
rect 21196 25284 21252 25294
rect 20076 23660 20244 23716
rect 19964 23650 20020 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 22878 19630 22930
rect 19682 22878 19684 22930
rect 19628 22866 19684 22878
rect 19852 23380 19908 23390
rect 19852 23042 19908 23324
rect 20188 23380 20244 23660
rect 20188 23314 20244 23324
rect 20356 23660 20468 23716
rect 20076 23268 20132 23278
rect 20076 23174 20132 23212
rect 20300 23268 20356 23660
rect 20300 23202 20356 23212
rect 20412 23492 20468 23502
rect 19852 22990 19854 23042
rect 19906 22990 19908 23042
rect 19852 22484 19908 22990
rect 19852 22418 19908 22428
rect 20412 22372 20468 23436
rect 20748 23380 20804 23390
rect 20748 23154 20804 23324
rect 21196 23380 21252 25228
rect 21420 25284 21476 26238
rect 21532 25508 21588 27468
rect 21756 27300 21812 28364
rect 22092 27524 22148 29374
rect 22764 29314 22820 29326
rect 22764 29262 22766 29314
rect 22818 29262 22820 29314
rect 22764 28644 22820 29262
rect 22764 28578 22820 28588
rect 22876 28418 22932 28430
rect 22876 28366 22878 28418
rect 22930 28366 22932 28418
rect 22092 27458 22148 27468
rect 22540 27746 22596 27758
rect 22540 27694 22542 27746
rect 22594 27694 22596 27746
rect 22540 27524 22596 27694
rect 22876 27748 22932 28366
rect 22988 27748 23044 27758
rect 22876 27692 22988 27748
rect 22988 27654 23044 27692
rect 22540 27458 22596 27468
rect 21644 27244 21812 27300
rect 21644 26516 21700 27244
rect 21644 26450 21700 26460
rect 21756 27074 21812 27086
rect 21756 27022 21758 27074
rect 21810 27022 21812 27074
rect 21756 26852 21812 27022
rect 22204 27074 22260 27086
rect 22204 27022 22206 27074
rect 22258 27022 22260 27074
rect 22204 26908 22260 27022
rect 22540 27076 22596 27114
rect 22540 27010 22596 27020
rect 23100 27074 23156 35420
rect 23324 35474 23380 35486
rect 23324 35422 23326 35474
rect 23378 35422 23380 35474
rect 23212 34914 23268 34926
rect 23212 34862 23214 34914
rect 23266 34862 23268 34914
rect 23212 34018 23268 34862
rect 23212 33966 23214 34018
rect 23266 33966 23268 34018
rect 23212 33124 23268 33966
rect 23324 33348 23380 35422
rect 23772 35140 23828 36206
rect 23884 36258 23940 36270
rect 23884 36206 23886 36258
rect 23938 36206 23940 36258
rect 23884 35924 23940 36206
rect 23884 35868 24052 35924
rect 23884 35700 23940 35710
rect 23884 35606 23940 35644
rect 23772 34244 23828 35084
rect 23884 35028 23940 35038
rect 23996 35028 24052 35868
rect 24444 35812 24500 37102
rect 24556 37044 24612 37436
rect 24668 37268 24724 37278
rect 25228 37268 25284 37278
rect 24668 37266 25284 37268
rect 24668 37214 24670 37266
rect 24722 37214 25230 37266
rect 25282 37214 25284 37266
rect 24668 37212 25284 37214
rect 24668 37202 24724 37212
rect 25228 37202 25284 37212
rect 25340 37044 25396 37996
rect 25564 37492 25620 40684
rect 25676 40290 25732 43148
rect 25788 41300 25844 41310
rect 25788 41186 25844 41244
rect 25788 41134 25790 41186
rect 25842 41134 25844 41186
rect 25788 41122 25844 41134
rect 25676 40238 25678 40290
rect 25730 40238 25732 40290
rect 25676 40226 25732 40238
rect 25676 39844 25732 39854
rect 25676 39618 25732 39788
rect 25676 39566 25678 39618
rect 25730 39566 25732 39618
rect 25676 39554 25732 39566
rect 24556 36978 24612 36988
rect 25116 36988 25396 37044
rect 25452 37436 25620 37492
rect 25900 37940 25956 43260
rect 26012 43092 26068 43484
rect 26012 43026 26068 43036
rect 26124 43538 26180 43550
rect 26124 43486 26126 43538
rect 26178 43486 26180 43538
rect 26124 42756 26180 43486
rect 26348 43540 26404 43550
rect 26348 42866 26404 43484
rect 26460 43538 26516 44044
rect 26684 43988 26740 43998
rect 26460 43486 26462 43538
rect 26514 43486 26516 43538
rect 26460 43474 26516 43486
rect 26572 43876 26628 43886
rect 26348 42814 26350 42866
rect 26402 42814 26404 42866
rect 26348 42802 26404 42814
rect 26124 42690 26180 42700
rect 26460 42756 26516 42766
rect 26460 42662 26516 42700
rect 26236 42644 26292 42654
rect 26236 42550 26292 42588
rect 26012 42532 26068 42542
rect 26012 41970 26068 42476
rect 26012 41918 26014 41970
rect 26066 41918 26068 41970
rect 26012 41906 26068 41918
rect 26460 41970 26516 41982
rect 26460 41918 26462 41970
rect 26514 41918 26516 41970
rect 26236 41746 26292 41758
rect 26236 41694 26238 41746
rect 26290 41694 26292 41746
rect 26012 41636 26068 41646
rect 26012 40402 26068 41580
rect 26236 41412 26292 41694
rect 26236 41346 26292 41356
rect 26236 41186 26292 41198
rect 26236 41134 26238 41186
rect 26290 41134 26292 41186
rect 26236 40628 26292 41134
rect 26236 40514 26292 40572
rect 26236 40462 26238 40514
rect 26290 40462 26292 40514
rect 26236 40450 26292 40462
rect 26012 40350 26014 40402
rect 26066 40350 26068 40402
rect 26012 40338 26068 40350
rect 26460 40404 26516 41918
rect 26572 41188 26628 43820
rect 26572 41122 26628 41132
rect 26460 40338 26516 40348
rect 26684 40180 26740 43932
rect 27356 43988 27412 43998
rect 26796 43876 26852 43886
rect 26796 43762 26852 43820
rect 26796 43710 26798 43762
rect 26850 43710 26852 43762
rect 26796 43698 26852 43710
rect 26908 43764 26964 43774
rect 26796 43316 26852 43326
rect 26796 42754 26852 43260
rect 26796 42702 26798 42754
rect 26850 42702 26852 42754
rect 26796 42690 26852 42702
rect 26908 42084 26964 43708
rect 27020 43652 27076 43662
rect 27020 43558 27076 43596
rect 27356 43538 27412 43932
rect 27356 43486 27358 43538
rect 27410 43486 27412 43538
rect 27132 43428 27188 43438
rect 27132 43334 27188 43372
rect 27356 42980 27412 43486
rect 27468 43092 27524 45054
rect 27580 43316 27636 45612
rect 27692 43540 27748 45724
rect 27804 45666 27860 45678
rect 27804 45614 27806 45666
rect 27858 45614 27860 45666
rect 27804 43988 27860 45614
rect 27916 45668 27972 46956
rect 28140 46788 28196 46798
rect 28252 46788 28308 48076
rect 28364 48066 28420 48076
rect 28476 47460 28532 49084
rect 29484 49140 29540 49150
rect 28588 49026 28644 49038
rect 28588 48974 28590 49026
rect 28642 48974 28644 49026
rect 28588 47572 28644 48974
rect 29148 49028 29204 49038
rect 29148 48934 29204 48972
rect 29484 49026 29540 49084
rect 29596 49138 29652 50372
rect 30156 49252 30212 55916
rect 30268 52836 30324 56030
rect 30716 55970 30772 56252
rect 30940 56308 30996 59200
rect 31388 56308 31444 59200
rect 32284 57092 32340 59200
rect 32284 57026 32340 57036
rect 31500 56308 31556 56318
rect 31388 56306 31556 56308
rect 31388 56254 31502 56306
rect 31554 56254 31556 56306
rect 31388 56252 31556 56254
rect 30940 56242 30996 56252
rect 31500 56242 31556 56252
rect 32620 56308 32676 56318
rect 32172 56084 32228 56094
rect 30716 55918 30718 55970
rect 30770 55918 30772 55970
rect 30716 55906 30772 55918
rect 32060 56082 32228 56084
rect 32060 56030 32174 56082
rect 32226 56030 32228 56082
rect 32060 56028 32228 56030
rect 32060 55410 32116 56028
rect 32172 56018 32228 56028
rect 32620 55970 32676 56252
rect 32620 55918 32622 55970
rect 32674 55918 32676 55970
rect 32620 55906 32676 55918
rect 32060 55358 32062 55410
rect 32114 55358 32116 55410
rect 32060 55346 32116 55358
rect 32508 55298 32564 55310
rect 32508 55246 32510 55298
rect 32562 55246 32564 55298
rect 30380 54514 30436 54526
rect 30380 54462 30382 54514
rect 30434 54462 30436 54514
rect 30380 53620 30436 54462
rect 30380 53554 30436 53564
rect 30940 54404 30996 54414
rect 30940 53730 30996 54348
rect 32060 54404 32116 54414
rect 32060 54310 32116 54348
rect 32508 54404 32564 55246
rect 32732 54740 32788 59200
rect 33628 56980 33684 59200
rect 33628 56914 33684 56924
rect 34076 56308 34132 59200
rect 34076 56242 34132 56252
rect 34188 57092 34244 57102
rect 33740 56084 33796 56094
rect 33628 56082 33796 56084
rect 33628 56030 33742 56082
rect 33794 56030 33796 56082
rect 33628 56028 33796 56030
rect 33180 55186 33236 55198
rect 33180 55134 33182 55186
rect 33234 55134 33236 55186
rect 33068 54740 33124 54750
rect 32732 54738 33124 54740
rect 32732 54686 33070 54738
rect 33122 54686 33124 54738
rect 32732 54684 33124 54686
rect 33068 54674 33124 54684
rect 32508 54310 32564 54348
rect 30940 53678 30942 53730
rect 30994 53678 30996 53730
rect 30828 53172 30884 53182
rect 30940 53172 30996 53678
rect 31612 53620 31668 53630
rect 31612 53618 32004 53620
rect 31612 53566 31614 53618
rect 31666 53566 32004 53618
rect 31612 53564 32004 53566
rect 31612 53554 31668 53564
rect 30492 53170 30996 53172
rect 30492 53118 30830 53170
rect 30882 53118 30996 53170
rect 30492 53116 30996 53118
rect 31948 53170 32004 53564
rect 31948 53118 31950 53170
rect 32002 53118 32004 53170
rect 30380 52836 30436 52846
rect 30268 52834 30436 52836
rect 30268 52782 30382 52834
rect 30434 52782 30436 52834
rect 30268 52780 30436 52782
rect 30380 52770 30436 52780
rect 30492 52162 30548 53116
rect 30828 53106 30884 53116
rect 31948 53106 32004 53118
rect 33180 53172 33236 55134
rect 33628 54292 33684 56028
rect 33740 56018 33796 56028
rect 33852 56084 33908 56094
rect 33852 54964 33908 56028
rect 34188 55970 34244 57036
rect 34972 57092 35028 59200
rect 35420 57316 35476 59200
rect 35420 57260 36260 57316
rect 34972 57026 35028 57036
rect 35308 56308 35364 56318
rect 35308 56214 35364 56252
rect 35980 56084 36036 56094
rect 35980 55990 36036 56028
rect 34188 55918 34190 55970
rect 34242 55918 34244 55970
rect 34188 55906 34244 55918
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35308 55524 35364 55534
rect 35308 55410 35364 55468
rect 35308 55358 35310 55410
rect 35362 55358 35364 55410
rect 35308 55346 35364 55358
rect 35980 55188 36036 55198
rect 36204 55188 36260 57260
rect 36316 55412 36372 59200
rect 36428 56980 36484 56990
rect 36428 55970 36484 56924
rect 36764 56308 36820 59200
rect 37660 56756 37716 59200
rect 38108 57316 38164 59200
rect 38108 57260 38612 57316
rect 37660 56690 37716 56700
rect 37996 57092 38052 57102
rect 36764 56242 36820 56252
rect 36428 55918 36430 55970
rect 36482 55918 36484 55970
rect 36428 55906 36484 55918
rect 37548 56082 37604 56094
rect 37548 56030 37550 56082
rect 37602 56030 37604 56082
rect 37548 55524 37604 56030
rect 37996 55970 38052 57036
rect 37996 55918 37998 55970
rect 38050 55918 38052 55970
rect 37996 55906 38052 55918
rect 37548 55458 37604 55468
rect 36316 55346 36372 55356
rect 37436 55412 37492 55422
rect 37436 55318 37492 55356
rect 38108 55300 38164 55310
rect 37772 55298 38164 55300
rect 37772 55246 38110 55298
rect 38162 55246 38164 55298
rect 37772 55244 38164 55246
rect 36316 55188 36372 55198
rect 35980 55186 36148 55188
rect 35980 55134 35982 55186
rect 36034 55134 36148 55186
rect 35980 55132 36148 55134
rect 36204 55186 36372 55188
rect 36204 55134 36318 55186
rect 36370 55134 36372 55186
rect 36204 55132 36372 55134
rect 35980 55122 36036 55132
rect 33180 53106 33236 53116
rect 33292 54236 33684 54292
rect 33740 54908 33908 54964
rect 35644 55074 35700 55086
rect 35644 55022 35646 55074
rect 35698 55022 35700 55074
rect 32284 52948 32340 52958
rect 32284 52854 32340 52892
rect 33292 52274 33348 54236
rect 33292 52222 33294 52274
rect 33346 52222 33348 52274
rect 33292 52210 33348 52222
rect 33516 54068 33572 54078
rect 30492 52110 30494 52162
rect 30546 52110 30548 52162
rect 30492 51604 30548 52110
rect 31164 52162 31220 52174
rect 31164 52110 31166 52162
rect 31218 52110 31220 52162
rect 31164 52052 31220 52110
rect 31164 51986 31220 51996
rect 30492 50428 30548 51548
rect 31836 51604 31892 51614
rect 33516 51604 33572 54012
rect 33740 53842 33796 54908
rect 35644 54626 35700 55022
rect 35644 54574 35646 54626
rect 35698 54574 35700 54626
rect 35644 54562 35700 54574
rect 34524 54516 34580 54526
rect 34860 54516 34916 54526
rect 34188 54514 34916 54516
rect 34188 54462 34526 54514
rect 34578 54462 34862 54514
rect 34914 54462 34916 54514
rect 34188 54460 34916 54462
rect 34188 54404 34244 54460
rect 34524 54450 34580 54460
rect 34860 54450 34916 54460
rect 34188 53844 34244 54348
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 36092 54068 36148 55132
rect 36316 55122 36372 55132
rect 37772 54402 37828 55244
rect 38108 55234 38164 55244
rect 38556 55186 38612 57260
rect 39004 56868 39060 59200
rect 39004 56802 39060 56812
rect 39228 56642 39284 56654
rect 39228 56590 39230 56642
rect 39282 56590 39284 56642
rect 39116 56308 39172 56318
rect 39116 56214 39172 56252
rect 39116 55300 39172 55310
rect 39228 55300 39284 56590
rect 39116 55298 39284 55300
rect 39116 55246 39118 55298
rect 39170 55246 39284 55298
rect 39116 55244 39284 55246
rect 39116 55234 39172 55244
rect 38556 55134 38558 55186
rect 38610 55134 38612 55186
rect 38556 55122 38612 55134
rect 39340 55074 39396 55086
rect 39340 55022 39342 55074
rect 39394 55022 39396 55074
rect 37772 54350 37774 54402
rect 37826 54350 37828 54402
rect 37772 54338 37828 54350
rect 39228 54514 39284 54526
rect 39228 54462 39230 54514
rect 39282 54462 39284 54514
rect 39116 54292 39172 54302
rect 39004 54236 39116 54292
rect 36092 54012 36932 54068
rect 35196 53844 35252 53854
rect 33740 53790 33742 53842
rect 33794 53790 33796 53842
rect 33740 53778 33796 53790
rect 33852 53842 34244 53844
rect 33852 53790 34190 53842
rect 34242 53790 34244 53842
rect 33852 53788 34244 53790
rect 33740 52276 33796 52286
rect 33852 52276 33908 53788
rect 34188 53778 34244 53788
rect 34300 53842 35252 53844
rect 34300 53790 35198 53842
rect 35250 53790 35252 53842
rect 34300 53788 35252 53790
rect 34076 53396 34132 53406
rect 33964 53172 34020 53182
rect 33964 53078 34020 53116
rect 34076 53170 34132 53340
rect 34076 53118 34078 53170
rect 34130 53118 34132 53170
rect 34076 53106 34132 53118
rect 34300 53170 34356 53788
rect 34748 53620 34804 53630
rect 34300 53118 34302 53170
rect 34354 53118 34356 53170
rect 34300 53106 34356 53118
rect 34524 53284 34580 53294
rect 33740 52274 33908 52276
rect 33740 52222 33742 52274
rect 33794 52222 33908 52274
rect 33740 52220 33908 52222
rect 34524 52946 34580 53228
rect 34748 53170 34804 53564
rect 34748 53118 34750 53170
rect 34802 53118 34804 53170
rect 34748 53106 34804 53118
rect 34524 52894 34526 52946
rect 34578 52894 34580 52946
rect 33740 52210 33796 52220
rect 33852 51604 33908 51614
rect 33516 51602 33908 51604
rect 33516 51550 33854 51602
rect 33906 51550 33908 51602
rect 33516 51548 33908 51550
rect 31836 51510 31892 51548
rect 33852 51538 33908 51548
rect 34188 51492 34244 51502
rect 34188 51398 34244 51436
rect 33964 51378 34020 51390
rect 33964 51326 33966 51378
rect 34018 51326 34020 51378
rect 31388 51268 31444 51278
rect 33964 51268 34020 51326
rect 34412 51380 34468 51390
rect 34412 51286 34468 51324
rect 31388 51266 31556 51268
rect 31388 51214 31390 51266
rect 31442 51214 31556 51266
rect 31388 51212 31556 51214
rect 31388 51202 31444 51212
rect 30716 50482 30772 50494
rect 30716 50430 30718 50482
rect 30770 50430 30772 50482
rect 30716 50428 30772 50430
rect 30492 50372 30772 50428
rect 30492 49700 30548 49710
rect 30492 49606 30548 49644
rect 30156 49186 30212 49196
rect 29596 49086 29598 49138
rect 29650 49086 29652 49138
rect 29596 49074 29652 49086
rect 30380 49140 30436 49150
rect 29484 48974 29486 49026
rect 29538 48974 29540 49026
rect 29484 48962 29540 48974
rect 28924 48916 28980 48926
rect 28812 48860 28924 48916
rect 28812 48466 28868 48860
rect 28924 48850 28980 48860
rect 30380 48914 30436 49084
rect 30380 48862 30382 48914
rect 30434 48862 30436 48914
rect 30380 48850 30436 48862
rect 28812 48414 28814 48466
rect 28866 48414 28868 48466
rect 28812 48402 28868 48414
rect 29372 48804 29428 48814
rect 28700 48244 28756 48254
rect 28700 47908 28756 48188
rect 28700 47842 28756 47852
rect 28924 48242 28980 48254
rect 28924 48190 28926 48242
rect 28978 48190 28980 48242
rect 28588 47516 28868 47572
rect 28476 47458 28756 47460
rect 28476 47406 28478 47458
rect 28530 47406 28756 47458
rect 28476 47404 28756 47406
rect 28476 47394 28532 47404
rect 28140 46786 28308 46788
rect 28140 46734 28142 46786
rect 28194 46734 28308 46786
rect 28140 46732 28308 46734
rect 28364 47346 28420 47358
rect 28364 47294 28366 47346
rect 28418 47294 28420 47346
rect 28140 46722 28196 46732
rect 28028 46676 28084 46686
rect 28028 46582 28084 46620
rect 28364 46340 28420 47294
rect 28028 46284 28420 46340
rect 28476 47236 28532 47246
rect 28476 46786 28532 47180
rect 28476 46734 28478 46786
rect 28530 46734 28532 46786
rect 28028 45892 28084 46284
rect 28476 46228 28532 46734
rect 28588 46788 28644 46798
rect 28588 46694 28644 46732
rect 28700 46676 28756 47404
rect 28812 46898 28868 47516
rect 28924 47460 28980 48190
rect 29372 48242 29428 48748
rect 29708 48804 29764 48814
rect 29708 48710 29764 48748
rect 30604 48356 30660 50372
rect 30716 49924 30772 49934
rect 30716 49026 30772 49868
rect 31164 49924 31220 49934
rect 30716 48974 30718 49026
rect 30770 48974 30772 49026
rect 30716 48962 30772 48974
rect 30828 49700 30884 49710
rect 30716 48356 30772 48366
rect 30604 48354 30772 48356
rect 30604 48302 30718 48354
rect 30770 48302 30772 48354
rect 30604 48300 30772 48302
rect 30716 48290 30772 48300
rect 29372 48190 29374 48242
rect 29426 48190 29428 48242
rect 29148 48132 29204 48142
rect 29148 48038 29204 48076
rect 29260 48020 29316 48030
rect 29036 47460 29092 47470
rect 28924 47404 29036 47460
rect 29036 47366 29092 47404
rect 28812 46846 28814 46898
rect 28866 46846 28868 46898
rect 28812 46834 28868 46846
rect 28924 47012 28980 47022
rect 29260 47012 29316 47964
rect 29372 47570 29428 48190
rect 29372 47518 29374 47570
rect 29426 47518 29428 47570
rect 29372 47506 29428 47518
rect 29596 48018 29652 48030
rect 29596 47966 29598 48018
rect 29650 47966 29652 48018
rect 29260 46956 29428 47012
rect 28924 46898 28980 46956
rect 28924 46846 28926 46898
rect 28978 46846 28980 46898
rect 28924 46834 28980 46846
rect 29148 46786 29204 46798
rect 29148 46734 29150 46786
rect 29202 46734 29204 46786
rect 29148 46676 29204 46734
rect 29260 46788 29316 46798
rect 29260 46694 29316 46732
rect 28700 46620 29204 46676
rect 28364 46172 28532 46228
rect 28028 45798 28084 45836
rect 28140 46004 28196 46014
rect 27916 45612 28084 45668
rect 27804 43922 27860 43932
rect 27916 45218 27972 45230
rect 27916 45166 27918 45218
rect 27970 45166 27972 45218
rect 27916 43764 27972 45166
rect 27916 43698 27972 43708
rect 28028 43652 28084 45612
rect 28140 43876 28196 45948
rect 28252 45778 28308 45790
rect 28252 45726 28254 45778
rect 28306 45726 28308 45778
rect 28252 45444 28308 45726
rect 28252 45378 28308 45388
rect 28364 44436 28420 46172
rect 29372 45892 29428 46956
rect 29484 46900 29540 46910
rect 29484 46564 29540 46844
rect 29484 46498 29540 46508
rect 29596 46788 29652 47966
rect 29708 47796 29764 47806
rect 29708 47570 29764 47740
rect 29708 47518 29710 47570
rect 29762 47518 29764 47570
rect 29708 47506 29764 47518
rect 29820 47572 29876 47582
rect 29820 47458 29876 47516
rect 29820 47406 29822 47458
rect 29874 47406 29876 47458
rect 29820 47394 29876 47406
rect 30828 47458 30884 49644
rect 30940 49586 30996 49598
rect 30940 49534 30942 49586
rect 30994 49534 30996 49586
rect 30940 48468 30996 49534
rect 30940 48402 30996 48412
rect 30828 47406 30830 47458
rect 30882 47406 30884 47458
rect 29708 46900 29764 46910
rect 30156 46900 30212 46910
rect 29708 46806 29764 46844
rect 29820 46844 30156 46900
rect 28588 45836 29204 45892
rect 28364 44370 28420 44380
rect 28476 44884 28532 44894
rect 28588 44884 28644 45836
rect 29148 45778 29204 45836
rect 29148 45726 29150 45778
rect 29202 45726 29204 45778
rect 29148 45714 29204 45726
rect 29260 45890 29428 45892
rect 29260 45838 29374 45890
rect 29426 45838 29428 45890
rect 29260 45836 29428 45838
rect 29260 45556 29316 45836
rect 29372 45826 29428 45836
rect 29484 46002 29540 46014
rect 29484 45950 29486 46002
rect 29538 45950 29540 46002
rect 28924 45500 29316 45556
rect 28924 45106 28980 45500
rect 29372 45444 29428 45454
rect 28924 45054 28926 45106
rect 28978 45054 28980 45106
rect 28924 45042 28980 45054
rect 29148 45332 29204 45342
rect 28532 44828 28644 44884
rect 28700 44994 28756 45006
rect 28700 44942 28702 44994
rect 28754 44942 28756 44994
rect 28252 44324 28308 44334
rect 28252 44230 28308 44268
rect 28476 44210 28532 44828
rect 28588 44548 28644 44558
rect 28588 44322 28644 44492
rect 28588 44270 28590 44322
rect 28642 44270 28644 44322
rect 28588 44258 28644 44270
rect 28476 44158 28478 44210
rect 28530 44158 28532 44210
rect 28476 44146 28532 44158
rect 28140 43810 28196 43820
rect 28700 43764 28756 44942
rect 29148 44546 29204 45276
rect 29260 45108 29316 45118
rect 29260 44994 29316 45052
rect 29260 44942 29262 44994
rect 29314 44942 29316 44994
rect 29260 44930 29316 44942
rect 29148 44494 29150 44546
rect 29202 44494 29204 44546
rect 29148 44482 29204 44494
rect 29372 44546 29428 45388
rect 29372 44494 29374 44546
rect 29426 44494 29428 44546
rect 29372 44482 29428 44494
rect 29484 44100 29540 45950
rect 29596 45890 29652 46732
rect 29820 46786 29876 46844
rect 30156 46806 30212 46844
rect 30828 46900 30884 47406
rect 30828 46834 30884 46844
rect 31052 47570 31108 47582
rect 31052 47518 31054 47570
rect 31106 47518 31108 47570
rect 29820 46734 29822 46786
rect 29874 46734 29876 46786
rect 29820 46722 29876 46734
rect 30492 46786 30548 46798
rect 30492 46734 30494 46786
rect 30546 46734 30548 46786
rect 30492 46676 30548 46734
rect 30940 46788 30996 46798
rect 30940 46694 30996 46732
rect 30828 46676 30884 46686
rect 30492 46674 30884 46676
rect 30492 46622 30830 46674
rect 30882 46622 30884 46674
rect 30492 46620 30884 46622
rect 29708 46452 29764 46462
rect 29708 46450 30100 46452
rect 29708 46398 29710 46450
rect 29762 46398 30100 46450
rect 29708 46396 30100 46398
rect 29708 46386 29764 46396
rect 29596 45838 29598 45890
rect 29650 45838 29652 45890
rect 29596 45826 29652 45838
rect 30044 45890 30100 46396
rect 30828 46228 30884 46620
rect 31052 46676 31108 47518
rect 31164 47458 31220 49868
rect 31500 49924 31556 51212
rect 33964 51202 34020 51212
rect 34412 50708 34468 50718
rect 34300 50596 34356 50606
rect 34300 50034 34356 50540
rect 34300 49982 34302 50034
rect 34354 49982 34356 50034
rect 34300 49970 34356 49982
rect 31836 49924 31892 49934
rect 31500 49922 31892 49924
rect 31500 49870 31502 49922
rect 31554 49870 31838 49922
rect 31890 49870 31892 49922
rect 31500 49868 31892 49870
rect 31500 49858 31556 49868
rect 31836 49858 31892 49868
rect 32172 49924 32228 49934
rect 32172 49830 32228 49868
rect 34188 49812 34244 49822
rect 34412 49812 34468 50652
rect 34524 50036 34580 52894
rect 34860 52052 34916 52062
rect 34860 51602 34916 51996
rect 34860 51550 34862 51602
rect 34914 51550 34916 51602
rect 34860 51538 34916 51550
rect 35084 51604 35140 53788
rect 35196 53778 35252 53788
rect 35980 53676 36372 53732
rect 35196 53620 35252 53630
rect 35196 52946 35252 53564
rect 35532 53618 35588 53630
rect 35532 53566 35534 53618
rect 35586 53566 35588 53618
rect 35196 52894 35198 52946
rect 35250 52894 35252 52946
rect 35196 52882 35252 52894
rect 35308 53506 35364 53518
rect 35308 53454 35310 53506
rect 35362 53454 35364 53506
rect 35308 53060 35364 53454
rect 35308 52724 35364 53004
rect 35308 52658 35364 52668
rect 35420 52836 35476 52846
rect 35420 52722 35476 52780
rect 35420 52670 35422 52722
rect 35474 52670 35476 52722
rect 35420 52658 35476 52670
rect 35532 52724 35588 53566
rect 35868 53618 35924 53630
rect 35868 53566 35870 53618
rect 35922 53566 35924 53618
rect 35868 53284 35924 53566
rect 35980 53618 36036 53676
rect 35980 53566 35982 53618
rect 36034 53566 36036 53618
rect 35980 53554 36036 53566
rect 35868 53218 35924 53228
rect 36204 53506 36260 53518
rect 36204 53454 36206 53506
rect 36258 53454 36260 53506
rect 36204 53060 36260 53454
rect 35644 53004 36260 53060
rect 35644 52946 35700 53004
rect 35644 52894 35646 52946
rect 35698 52894 35700 52946
rect 35644 52882 35700 52894
rect 36204 52946 36260 53004
rect 36204 52894 36206 52946
rect 36258 52894 36260 52946
rect 36204 52882 36260 52894
rect 35980 52834 36036 52846
rect 35980 52782 35982 52834
rect 36034 52782 36036 52834
rect 35980 52724 36036 52782
rect 36316 52724 36372 53676
rect 36876 53170 36932 54012
rect 38556 53844 38612 53854
rect 38556 53750 38612 53788
rect 37884 53732 37940 53742
rect 37772 53676 37884 53732
rect 37772 53618 37828 53676
rect 37884 53666 37940 53676
rect 38332 53732 38388 53742
rect 37772 53566 37774 53618
rect 37826 53566 37828 53618
rect 37772 53554 37828 53566
rect 37996 53620 38052 53630
rect 36876 53118 36878 53170
rect 36930 53118 36932 53170
rect 36876 53106 36932 53118
rect 37884 53506 37940 53518
rect 37884 53454 37886 53506
rect 37938 53454 37940 53506
rect 37212 52948 37268 52958
rect 37884 52948 37940 53454
rect 37212 52854 37268 52892
rect 37772 52892 37884 52948
rect 35532 52668 36148 52724
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35644 52500 35700 52510
rect 35532 52276 35588 52286
rect 35308 51940 35364 51950
rect 35196 51604 35252 51614
rect 35084 51602 35252 51604
rect 35084 51550 35198 51602
rect 35250 51550 35252 51602
rect 35084 51548 35252 51550
rect 35196 51538 35252 51548
rect 34636 51378 34692 51390
rect 34636 51326 34638 51378
rect 34690 51326 34692 51378
rect 34636 50818 34692 51326
rect 34972 51378 35028 51390
rect 34972 51326 34974 51378
rect 35026 51326 35028 51378
rect 34972 51268 35028 51326
rect 34972 51202 35028 51212
rect 34636 50766 34638 50818
rect 34690 50766 34692 50818
rect 34636 50754 34692 50766
rect 34748 51156 34804 51166
rect 35308 51156 35364 51884
rect 35532 51604 35588 52220
rect 35644 51828 35700 52444
rect 36092 52274 36148 52668
rect 36092 52222 36094 52274
rect 36146 52222 36148 52274
rect 36092 52210 36148 52222
rect 36204 52388 36260 52398
rect 35756 52052 35812 52062
rect 35756 51958 35812 51996
rect 36204 52050 36260 52332
rect 36316 52276 36372 52668
rect 36316 52210 36372 52220
rect 36428 52722 36484 52734
rect 36428 52670 36430 52722
rect 36482 52670 36484 52722
rect 36204 51998 36206 52050
rect 36258 51998 36260 52050
rect 36204 51986 36260 51998
rect 36316 52052 36372 52062
rect 35980 51940 36036 51950
rect 35868 51938 36036 51940
rect 35868 51886 35982 51938
rect 36034 51886 36036 51938
rect 35868 51884 36036 51886
rect 35644 51772 35812 51828
rect 35420 51492 35476 51502
rect 35420 51398 35476 51436
rect 34748 50482 34804 51100
rect 35084 51100 35364 51156
rect 34972 50820 35028 50830
rect 35084 50820 35140 51100
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 34972 50818 35364 50820
rect 34972 50766 34974 50818
rect 35026 50766 35364 50818
rect 34972 50764 35364 50766
rect 34972 50754 35028 50764
rect 34748 50430 34750 50482
rect 34802 50430 34804 50482
rect 34748 50418 34804 50430
rect 35084 50484 35140 50494
rect 34524 49980 34804 50036
rect 34524 49812 34580 49822
rect 34188 49810 34580 49812
rect 34188 49758 34190 49810
rect 34242 49758 34526 49810
rect 34578 49758 34580 49810
rect 34188 49756 34580 49758
rect 34188 49746 34244 49756
rect 34524 49746 34580 49756
rect 31276 49700 31332 49710
rect 31276 49606 31332 49644
rect 33964 49698 34020 49710
rect 33964 49646 33966 49698
rect 34018 49646 34020 49698
rect 31276 49028 31332 49038
rect 31276 48934 31332 48972
rect 33964 49028 34020 49646
rect 34748 49698 34804 49980
rect 35084 50034 35140 50428
rect 35308 50370 35364 50764
rect 35420 50596 35476 50606
rect 35420 50502 35476 50540
rect 35308 50318 35310 50370
rect 35362 50318 35364 50370
rect 35308 50306 35364 50318
rect 35084 49982 35086 50034
rect 35138 49982 35140 50034
rect 35084 49970 35140 49982
rect 34860 49812 34916 49822
rect 34860 49718 34916 49756
rect 35532 49810 35588 51548
rect 35644 51380 35700 51390
rect 35644 51044 35700 51324
rect 35644 50978 35700 50988
rect 35532 49758 35534 49810
rect 35586 49758 35588 49810
rect 35532 49746 35588 49758
rect 35644 50594 35700 50606
rect 35644 50542 35646 50594
rect 35698 50542 35700 50594
rect 35644 49812 35700 50542
rect 34748 49646 34750 49698
rect 34802 49646 34804 49698
rect 34748 49634 34804 49646
rect 34300 49476 34356 49486
rect 31948 48916 32004 48926
rect 31948 48822 32004 48860
rect 33404 48916 33460 48926
rect 33180 48356 33236 48366
rect 31836 48244 31892 48254
rect 31836 47570 31892 48188
rect 32508 48244 32564 48254
rect 32508 48150 32564 48188
rect 33068 47908 33124 47918
rect 33068 47682 33124 47852
rect 33068 47630 33070 47682
rect 33122 47630 33124 47682
rect 33068 47618 33124 47630
rect 31836 47518 31838 47570
rect 31890 47518 31892 47570
rect 31836 47506 31892 47518
rect 31164 47406 31166 47458
rect 31218 47406 31220 47458
rect 31164 46788 31220 47406
rect 31388 47460 31444 47470
rect 31388 47346 31444 47404
rect 31388 47294 31390 47346
rect 31442 47294 31444 47346
rect 31388 47282 31444 47294
rect 32172 47458 32228 47470
rect 32172 47406 32174 47458
rect 32226 47406 32228 47458
rect 32172 47012 32228 47406
rect 32732 47460 32788 47470
rect 33180 47460 33236 48300
rect 32788 47458 33236 47460
rect 32788 47406 33182 47458
rect 33234 47406 33236 47458
rect 32788 47404 33236 47406
rect 32732 47366 32788 47404
rect 33180 47394 33236 47404
rect 33292 48244 33348 48254
rect 33292 47124 33348 48188
rect 33292 47058 33348 47068
rect 31164 46694 31220 46732
rect 31948 46956 32228 47012
rect 32508 47012 32564 47022
rect 33068 47012 33124 47022
rect 32564 46956 32676 47012
rect 31052 46610 31108 46620
rect 31276 46676 31332 46686
rect 30828 46172 31220 46228
rect 30044 45838 30046 45890
rect 30098 45838 30100 45890
rect 30044 45826 30100 45838
rect 31052 45890 31108 45902
rect 31052 45838 31054 45890
rect 31106 45838 31108 45890
rect 30156 45780 30212 45790
rect 30716 45780 30772 45790
rect 31052 45780 31108 45838
rect 30156 45686 30212 45724
rect 30268 45778 31108 45780
rect 30268 45726 30718 45778
rect 30770 45726 31108 45778
rect 30268 45724 31108 45726
rect 30044 45220 30100 45230
rect 29820 45108 29876 45118
rect 29596 44994 29652 45006
rect 29596 44942 29598 44994
rect 29650 44942 29652 44994
rect 29596 44548 29652 44942
rect 29596 44482 29652 44492
rect 28364 43708 28756 43764
rect 29036 44044 29540 44100
rect 29596 44322 29652 44334
rect 29596 44270 29598 44322
rect 29650 44270 29652 44322
rect 28140 43652 28196 43662
rect 28028 43596 28140 43652
rect 28140 43586 28196 43596
rect 27804 43540 27860 43550
rect 27692 43538 27860 43540
rect 27692 43486 27806 43538
rect 27858 43486 27860 43538
rect 27692 43484 27860 43486
rect 27804 43474 27860 43484
rect 28252 43538 28308 43550
rect 28252 43486 28254 43538
rect 28306 43486 28308 43538
rect 27580 43260 28196 43316
rect 27468 43026 27524 43036
rect 27356 42868 27412 42924
rect 27580 42868 27636 42878
rect 27356 42866 27636 42868
rect 27356 42814 27582 42866
rect 27634 42814 27636 42866
rect 27356 42812 27636 42814
rect 27132 42756 27188 42766
rect 27132 42644 27188 42700
rect 27580 42644 27636 42812
rect 27132 42642 27412 42644
rect 27132 42590 27134 42642
rect 27186 42590 27412 42642
rect 27132 42588 27412 42590
rect 27132 42578 27188 42588
rect 27132 42084 27188 42094
rect 26908 42028 27132 42084
rect 27132 41990 27188 42028
rect 27244 42082 27300 42094
rect 27244 42030 27246 42082
rect 27298 42030 27300 42082
rect 26796 41860 26852 41870
rect 26796 41186 26852 41804
rect 27244 41860 27300 42030
rect 27356 41972 27412 42588
rect 27580 42578 27636 42588
rect 27916 42868 27972 42878
rect 27468 42196 27524 42206
rect 27468 42102 27524 42140
rect 27580 42028 27860 42084
rect 27580 41972 27636 42028
rect 27356 41916 27636 41972
rect 27804 41970 27860 42028
rect 27804 41918 27806 41970
rect 27858 41918 27860 41970
rect 27804 41906 27860 41918
rect 27244 41794 27300 41804
rect 27692 41860 27748 41870
rect 27692 41766 27748 41804
rect 27916 41636 27972 42812
rect 28028 42530 28084 42542
rect 28028 42478 28030 42530
rect 28082 42478 28084 42530
rect 28028 42420 28084 42478
rect 28140 42532 28196 43260
rect 28252 42754 28308 43486
rect 28252 42702 28254 42754
rect 28306 42702 28308 42754
rect 28252 42690 28308 42702
rect 28140 42476 28308 42532
rect 28028 42354 28084 42364
rect 27468 41580 27972 41636
rect 28140 41970 28196 41982
rect 28140 41918 28142 41970
rect 28194 41918 28196 41970
rect 26796 41134 26798 41186
rect 26850 41134 26852 41186
rect 26796 41122 26852 41134
rect 27132 41186 27188 41198
rect 27132 41134 27134 41186
rect 27186 41134 27188 41186
rect 27132 40740 27188 41134
rect 26684 40114 26740 40124
rect 26796 40684 27188 40740
rect 26796 40514 26852 40684
rect 26796 40462 26798 40514
rect 26850 40462 26852 40514
rect 26684 39844 26740 39854
rect 26796 39844 26852 40462
rect 26908 40516 26964 40526
rect 27356 40516 27412 40526
rect 26908 40514 27412 40516
rect 26908 40462 26910 40514
rect 26962 40462 27358 40514
rect 27410 40462 27412 40514
rect 26908 40460 27412 40462
rect 26908 40450 26964 40460
rect 27356 40450 27412 40460
rect 27468 40514 27524 41580
rect 27580 41412 27636 41422
rect 27580 41318 27636 41356
rect 27468 40462 27470 40514
rect 27522 40462 27524 40514
rect 26908 40292 26964 40302
rect 27468 40292 27524 40462
rect 27692 41186 27748 41198
rect 27692 41134 27694 41186
rect 27746 41134 27748 41186
rect 27692 40404 27748 41134
rect 28140 40404 28196 41918
rect 27692 40402 28196 40404
rect 27692 40350 28142 40402
rect 28194 40350 28196 40402
rect 27692 40348 28196 40350
rect 26908 40178 26964 40236
rect 26908 40126 26910 40178
rect 26962 40126 26964 40178
rect 26908 40114 26964 40126
rect 27244 40236 27524 40292
rect 26684 39842 26852 39844
rect 26684 39790 26686 39842
rect 26738 39790 26852 39842
rect 26684 39788 26852 39790
rect 26908 39956 26964 39966
rect 26684 39778 26740 39788
rect 26572 39620 26628 39630
rect 26572 39526 26628 39564
rect 26012 39508 26068 39518
rect 26012 39414 26068 39452
rect 26684 39394 26740 39406
rect 26684 39342 26686 39394
rect 26738 39342 26740 39394
rect 26684 39060 26740 39342
rect 26012 38724 26068 38762
rect 26460 38724 26516 38734
rect 26012 38722 26516 38724
rect 26012 38670 26014 38722
rect 26066 38670 26462 38722
rect 26514 38670 26516 38722
rect 26012 38668 26516 38670
rect 26012 38612 26068 38668
rect 26460 38658 26516 38668
rect 26012 38546 26068 38556
rect 24444 35746 24500 35756
rect 24556 36258 24612 36270
rect 24556 36206 24558 36258
rect 24610 36206 24612 36258
rect 24556 35140 24612 36206
rect 24892 36258 24948 36270
rect 24892 36206 24894 36258
rect 24946 36206 24948 36258
rect 24892 35924 24948 36206
rect 24892 35858 24948 35868
rect 24556 35074 24612 35084
rect 23884 35026 24052 35028
rect 23884 34974 23886 35026
rect 23938 34974 24052 35026
rect 23884 34972 24052 34974
rect 23884 34962 23940 34972
rect 23772 34178 23828 34188
rect 24668 34356 24724 34366
rect 24668 34130 24724 34300
rect 24668 34078 24670 34130
rect 24722 34078 24724 34130
rect 24668 34066 24724 34078
rect 24444 34018 24500 34030
rect 24444 33966 24446 34018
rect 24498 33966 24500 34018
rect 24332 33908 24388 33918
rect 24332 33814 24388 33852
rect 24444 33458 24500 33966
rect 24444 33406 24446 33458
rect 24498 33406 24500 33458
rect 24444 33394 24500 33406
rect 23324 33292 23492 33348
rect 23324 33124 23380 33134
rect 23212 33122 23380 33124
rect 23212 33070 23326 33122
rect 23378 33070 23380 33122
rect 23212 33068 23380 33070
rect 23324 33012 23380 33068
rect 23324 32946 23380 32956
rect 23324 30882 23380 30894
rect 23324 30830 23326 30882
rect 23378 30830 23380 30882
rect 23324 30436 23380 30830
rect 23324 30370 23380 30380
rect 23436 29764 23492 33292
rect 23660 33346 23716 33358
rect 23660 33294 23662 33346
rect 23714 33294 23716 33346
rect 23660 33012 23716 33294
rect 24892 33124 24948 33134
rect 23660 32946 23716 32956
rect 24444 33012 24500 33022
rect 23660 32564 23716 32574
rect 23660 32470 23716 32508
rect 24444 32562 24500 32956
rect 24444 32510 24446 32562
rect 24498 32510 24500 32562
rect 24444 31220 24500 32510
rect 24892 31890 24948 33068
rect 24892 31838 24894 31890
rect 24946 31838 24948 31890
rect 24892 31826 24948 31838
rect 25004 31668 25060 31678
rect 25004 31574 25060 31612
rect 24668 31220 24724 31230
rect 24444 31164 24668 31220
rect 24668 31126 24724 31164
rect 23436 29698 23492 29708
rect 24108 30770 24164 30782
rect 24108 30718 24110 30770
rect 24162 30718 24164 30770
rect 24108 30100 24164 30718
rect 23660 29540 23716 29550
rect 23660 29538 23828 29540
rect 23660 29486 23662 29538
rect 23714 29486 23828 29538
rect 23660 29484 23828 29486
rect 23660 29474 23716 29484
rect 23436 28644 23492 28654
rect 23436 28550 23492 28588
rect 23436 27748 23492 27758
rect 23436 27076 23492 27692
rect 23100 27022 23102 27074
rect 23154 27022 23156 27074
rect 23100 26908 23156 27022
rect 23324 27074 23492 27076
rect 23324 27022 23438 27074
rect 23490 27022 23492 27074
rect 23324 27020 23492 27022
rect 22204 26852 22596 26908
rect 21644 26290 21700 26302
rect 21644 26238 21646 26290
rect 21698 26238 21700 26290
rect 21644 26068 21700 26238
rect 21644 26002 21700 26012
rect 21644 25508 21700 25518
rect 21532 25506 21700 25508
rect 21532 25454 21646 25506
rect 21698 25454 21700 25506
rect 21532 25452 21700 25454
rect 21420 25218 21476 25228
rect 21644 24724 21700 25452
rect 21756 25284 21812 26796
rect 22428 26628 22484 26638
rect 22316 26572 22428 26628
rect 22540 26628 22596 26852
rect 22652 26852 22708 26862
rect 22652 26758 22708 26796
rect 22876 26850 22932 26862
rect 23100 26852 23268 26908
rect 22876 26798 22878 26850
rect 22930 26798 22932 26850
rect 22876 26740 22932 26798
rect 22876 26684 23156 26740
rect 22540 26572 22820 26628
rect 21868 26404 21924 26414
rect 22316 26404 22372 26572
rect 22428 26562 22484 26572
rect 22764 26514 22820 26572
rect 23100 26516 23156 26684
rect 23212 26628 23268 26852
rect 23212 26562 23268 26572
rect 22764 26462 22766 26514
rect 22818 26462 22820 26514
rect 22764 26450 22820 26462
rect 22988 26460 23156 26516
rect 21868 26402 22372 26404
rect 21868 26350 21870 26402
rect 21922 26350 22372 26402
rect 21868 26348 22372 26350
rect 21868 26338 21924 26348
rect 22316 26290 22372 26348
rect 22540 26404 22596 26414
rect 22540 26310 22596 26348
rect 22988 26402 23044 26460
rect 22988 26350 22990 26402
rect 23042 26350 23044 26402
rect 22316 26238 22318 26290
rect 22370 26238 22372 26290
rect 22316 26226 22372 26238
rect 22988 26068 23044 26350
rect 23100 26292 23156 26302
rect 23100 26198 23156 26236
rect 22988 26002 23044 26012
rect 22540 25396 22596 25406
rect 21980 25284 22036 25294
rect 21756 25228 21980 25284
rect 21980 24948 22036 25228
rect 22316 24948 22372 24958
rect 21980 24946 22372 24948
rect 21980 24894 22318 24946
rect 22370 24894 22372 24946
rect 21980 24892 22372 24894
rect 22540 24948 22596 25340
rect 22652 25284 22708 25294
rect 23100 25284 23156 25294
rect 23324 25284 23380 27020
rect 23436 27010 23492 27020
rect 23772 26908 23828 29484
rect 23996 29426 24052 29438
rect 23996 29374 23998 29426
rect 24050 29374 24052 29426
rect 23996 27860 24052 29374
rect 23996 27766 24052 27804
rect 24108 28644 24164 30044
rect 24668 29428 24724 29466
rect 24668 29362 24724 29372
rect 24332 29204 24388 29214
rect 24668 29204 24724 29214
rect 24332 29202 24500 29204
rect 24332 29150 24334 29202
rect 24386 29150 24500 29202
rect 24332 29148 24500 29150
rect 24332 29138 24388 29148
rect 24108 27746 24164 28588
rect 24332 28868 24388 28878
rect 24332 27858 24388 28812
rect 24332 27806 24334 27858
rect 24386 27806 24388 27858
rect 24332 27794 24388 27806
rect 24108 27694 24110 27746
rect 24162 27694 24164 27746
rect 24108 27682 24164 27694
rect 23660 26852 23828 26908
rect 24220 26962 24276 26974
rect 24220 26910 24222 26962
rect 24274 26910 24276 26962
rect 23548 26516 23604 26526
rect 23548 26290 23604 26460
rect 23548 26238 23550 26290
rect 23602 26238 23604 26290
rect 23548 26226 23604 26238
rect 23548 25620 23604 25630
rect 23660 25620 23716 26852
rect 24220 26514 24276 26910
rect 24444 26908 24500 29148
rect 24668 29110 24724 29148
rect 24892 28644 24948 28654
rect 24556 28642 24948 28644
rect 24556 28590 24894 28642
rect 24946 28590 24948 28642
rect 24556 28588 24948 28590
rect 24556 27746 24612 28588
rect 24892 28578 24948 28588
rect 24556 27694 24558 27746
rect 24610 27694 24612 27746
rect 24556 27682 24612 27694
rect 25116 26908 25172 36988
rect 25228 36820 25284 36830
rect 25228 36370 25284 36764
rect 25228 36318 25230 36370
rect 25282 36318 25284 36370
rect 25228 36306 25284 36318
rect 25452 36036 25508 37436
rect 25564 37268 25620 37278
rect 25564 36260 25620 37212
rect 25900 37266 25956 37884
rect 26572 37940 26628 37950
rect 26684 37940 26740 39004
rect 26572 37938 26740 37940
rect 26572 37886 26574 37938
rect 26626 37886 26740 37938
rect 26572 37884 26740 37886
rect 26572 37874 26628 37884
rect 26012 37828 26068 37838
rect 26236 37828 26292 37838
rect 26012 37826 26292 37828
rect 26012 37774 26014 37826
rect 26066 37774 26238 37826
rect 26290 37774 26292 37826
rect 26012 37772 26292 37774
rect 26012 37762 26068 37772
rect 25900 37214 25902 37266
rect 25954 37214 25956 37266
rect 25900 37202 25956 37214
rect 26124 37156 26180 37166
rect 26236 37156 26292 37772
rect 26684 37156 26740 37166
rect 26124 37154 26740 37156
rect 26124 37102 26126 37154
rect 26178 37102 26686 37154
rect 26738 37102 26740 37154
rect 26124 37100 26740 37102
rect 26124 37090 26180 37100
rect 25900 36372 25956 36382
rect 25956 36316 26068 36372
rect 25900 36306 25956 36316
rect 25564 36258 25732 36260
rect 25564 36206 25566 36258
rect 25618 36206 25732 36258
rect 25564 36204 25732 36206
rect 25564 36194 25620 36204
rect 25228 35980 25508 36036
rect 25228 35922 25284 35980
rect 25228 35870 25230 35922
rect 25282 35870 25284 35922
rect 25228 35252 25284 35870
rect 25564 35924 25620 35934
rect 25564 35830 25620 35868
rect 25228 35186 25284 35196
rect 25676 35028 25732 36204
rect 26012 35588 26068 36316
rect 26124 35700 26180 35710
rect 26180 35644 26516 35700
rect 26124 35606 26180 35644
rect 26012 35252 26068 35532
rect 26012 35196 26180 35252
rect 26012 35028 26068 35038
rect 25676 35026 26068 35028
rect 25676 34974 26014 35026
rect 26066 34974 26068 35026
rect 25676 34972 26068 34974
rect 26012 34962 26068 34972
rect 26124 34804 26180 35196
rect 26460 34914 26516 35644
rect 26460 34862 26462 34914
rect 26514 34862 26516 34914
rect 26460 34850 26516 34862
rect 25900 34748 26180 34804
rect 25452 34356 25508 34366
rect 25452 34262 25508 34300
rect 25900 34242 25956 34748
rect 25900 34190 25902 34242
rect 25954 34190 25956 34242
rect 25900 34178 25956 34190
rect 25340 34132 25396 34142
rect 25340 32002 25396 34076
rect 26460 34132 26516 34142
rect 26460 34038 26516 34076
rect 26012 33908 26068 33918
rect 26012 33814 26068 33852
rect 25340 31950 25342 32002
rect 25394 31950 25396 32002
rect 25340 31938 25396 31950
rect 25676 31892 25732 31902
rect 26460 31892 26516 31902
rect 25676 31890 26516 31892
rect 25676 31838 25678 31890
rect 25730 31838 26462 31890
rect 26514 31838 26516 31890
rect 25676 31836 26516 31838
rect 25676 31826 25732 31836
rect 25564 31666 25620 31678
rect 26012 31668 26068 31678
rect 26236 31668 26292 31678
rect 25564 31614 25566 31666
rect 25618 31614 25620 31666
rect 25564 31556 25620 31614
rect 25788 31612 26012 31668
rect 25676 31556 25732 31566
rect 25564 31500 25676 31556
rect 25676 31490 25732 31500
rect 25228 30882 25284 30894
rect 25228 30830 25230 30882
rect 25282 30830 25284 30882
rect 25228 30436 25284 30830
rect 25228 30370 25284 30380
rect 25788 30210 25844 31612
rect 26012 31574 26068 31612
rect 26124 31666 26292 31668
rect 26124 31614 26238 31666
rect 26290 31614 26292 31666
rect 26124 31612 26292 31614
rect 26124 31556 26180 31612
rect 26236 31602 26292 31612
rect 26124 30324 26180 31500
rect 26348 30434 26404 31836
rect 26460 31826 26516 31836
rect 26348 30382 26350 30434
rect 26402 30382 26404 30434
rect 26348 30370 26404 30382
rect 26460 31554 26516 31566
rect 26460 31502 26462 31554
rect 26514 31502 26516 31554
rect 26124 30212 26180 30268
rect 25788 30158 25790 30210
rect 25842 30158 25844 30210
rect 25788 30146 25844 30158
rect 25900 30210 26180 30212
rect 25900 30158 26126 30210
rect 26178 30158 26180 30210
rect 25900 30156 26180 30158
rect 25340 29988 25396 29998
rect 25228 29314 25284 29326
rect 25228 29262 25230 29314
rect 25282 29262 25284 29314
rect 25228 28868 25284 29262
rect 25228 28802 25284 28812
rect 25340 28754 25396 29932
rect 25340 28702 25342 28754
rect 25394 28702 25396 28754
rect 25340 28690 25396 28702
rect 25452 29428 25508 29438
rect 25228 28644 25284 28654
rect 25228 28550 25284 28588
rect 25452 28644 25508 29372
rect 25900 29426 25956 30156
rect 26124 30146 26180 30156
rect 25900 29374 25902 29426
rect 25954 29374 25956 29426
rect 25900 29362 25956 29374
rect 24220 26462 24222 26514
rect 24274 26462 24276 26514
rect 24220 26450 24276 26462
rect 24332 26852 24500 26908
rect 25004 26852 25172 26908
rect 24108 26290 24164 26302
rect 24108 26238 24110 26290
rect 24162 26238 24164 26290
rect 23884 26180 23940 26190
rect 23884 26086 23940 26124
rect 23604 25564 23716 25620
rect 23548 25506 23604 25564
rect 23548 25454 23550 25506
rect 23602 25454 23604 25506
rect 23548 25442 23604 25454
rect 23996 25508 24052 25518
rect 24108 25508 24164 26238
rect 24332 26292 24388 26852
rect 24332 26198 24388 26236
rect 24892 26068 24948 26078
rect 24444 25620 24500 25630
rect 24332 25508 24388 25518
rect 24108 25506 24388 25508
rect 24108 25454 24334 25506
rect 24386 25454 24388 25506
rect 24108 25452 24388 25454
rect 23996 25414 24052 25452
rect 24332 25396 24388 25452
rect 24332 25330 24388 25340
rect 22652 25282 23380 25284
rect 22652 25230 22654 25282
rect 22706 25230 23102 25282
rect 23154 25230 23380 25282
rect 22652 25228 23380 25230
rect 22652 25218 22708 25228
rect 23100 25218 23156 25228
rect 22764 24948 22820 24958
rect 22540 24946 22820 24948
rect 22540 24894 22766 24946
rect 22818 24894 22820 24946
rect 22540 24892 22820 24894
rect 22316 24882 22372 24892
rect 22764 24882 22820 24892
rect 23100 24836 23156 24846
rect 21644 24722 22036 24724
rect 21644 24670 21646 24722
rect 21698 24670 22036 24722
rect 21644 24668 22036 24670
rect 21644 24658 21700 24668
rect 21308 24610 21364 24622
rect 21308 24558 21310 24610
rect 21362 24558 21364 24610
rect 21308 23492 21364 24558
rect 21980 23938 22036 24668
rect 21980 23886 21982 23938
rect 22034 23886 22036 23938
rect 21980 23874 22036 23886
rect 22092 24498 22148 24510
rect 22092 24446 22094 24498
rect 22146 24446 22148 24498
rect 21532 23828 21588 23838
rect 21532 23734 21588 23772
rect 21868 23828 21924 23838
rect 21308 23426 21364 23436
rect 21196 23314 21252 23324
rect 21756 23380 21812 23390
rect 20748 23102 20750 23154
rect 20802 23102 20804 23154
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19516 21756 19908 21812
rect 19852 21698 19908 21756
rect 19852 21646 19854 21698
rect 19906 21646 19908 21698
rect 19852 21634 19908 21646
rect 19964 21700 20020 21710
rect 19180 20638 19182 20690
rect 19234 20638 19236 20690
rect 18620 20580 18676 20590
rect 18620 20486 18676 20524
rect 18620 20020 18676 20030
rect 19068 20020 19124 20030
rect 18620 20018 19124 20020
rect 18620 19966 18622 20018
rect 18674 19966 19070 20018
rect 19122 19966 19124 20018
rect 18620 19964 19124 19966
rect 18620 19954 18676 19964
rect 19068 19954 19124 19964
rect 19180 19796 19236 20638
rect 19964 20692 20020 21644
rect 20188 21588 20244 21598
rect 20188 21494 20244 21532
rect 20412 20914 20468 22316
rect 20636 22372 20692 22382
rect 20748 22372 20804 23102
rect 20636 22370 20804 22372
rect 20636 22318 20638 22370
rect 20690 22318 20804 22370
rect 20636 22316 20804 22318
rect 20524 21924 20580 21934
rect 20636 21924 20692 22316
rect 20580 21868 20692 21924
rect 21532 21924 21588 21934
rect 20524 21586 20580 21868
rect 20524 21534 20526 21586
rect 20578 21534 20580 21586
rect 20524 21522 20580 21534
rect 20860 21588 20916 21598
rect 20860 21494 20916 21532
rect 20636 21362 20692 21374
rect 20636 21310 20638 21362
rect 20690 21310 20692 21362
rect 20524 21028 20580 21038
rect 20636 21028 20692 21310
rect 21308 21364 21364 21374
rect 21308 21362 21476 21364
rect 21308 21310 21310 21362
rect 21362 21310 21476 21362
rect 21308 21308 21476 21310
rect 21308 21298 21364 21308
rect 20524 21026 20692 21028
rect 20524 20974 20526 21026
rect 20578 20974 20692 21026
rect 20524 20972 20692 20974
rect 20524 20962 20580 20972
rect 20412 20862 20414 20914
rect 20466 20862 20468 20914
rect 20412 20850 20468 20862
rect 19964 20626 20020 20636
rect 20300 20804 20356 20814
rect 19628 20468 19684 20478
rect 19628 20132 19684 20412
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19964 20132 20020 20142
rect 19628 20130 20020 20132
rect 19628 20078 19966 20130
rect 20018 20078 20020 20130
rect 19628 20076 20020 20078
rect 19964 20066 20020 20076
rect 20188 20132 20244 20142
rect 20188 20018 20244 20076
rect 20188 19966 20190 20018
rect 20242 19966 20244 20018
rect 20188 19954 20244 19966
rect 18844 19740 19236 19796
rect 19404 19796 19460 19806
rect 18732 15874 18788 15886
rect 18732 15822 18734 15874
rect 18786 15822 18788 15874
rect 18732 15764 18788 15822
rect 18732 15698 18788 15708
rect 18508 14466 18564 14476
rect 15708 14418 15988 14420
rect 15708 14366 15934 14418
rect 15986 14366 15988 14418
rect 15708 14364 15988 14366
rect 15820 11788 15876 14364
rect 15932 14354 15988 14364
rect 16044 14364 16324 14420
rect 15932 13972 15988 13982
rect 16044 13972 16100 14364
rect 15932 13970 16100 13972
rect 15932 13918 15934 13970
rect 15986 13918 16100 13970
rect 15932 13916 16100 13918
rect 17164 14306 17220 14318
rect 17164 14254 17166 14306
rect 17218 14254 17220 14306
rect 15932 13906 15988 13916
rect 16604 13636 16660 13646
rect 16492 13580 16604 13636
rect 15596 11732 15876 11788
rect 16380 12516 16436 12526
rect 15372 11620 15428 11630
rect 15372 10724 15428 11564
rect 15372 9042 15428 10668
rect 15484 11396 15540 11406
rect 15596 11396 15652 11732
rect 15540 11340 15652 11396
rect 15708 11508 15764 11518
rect 15708 11394 15764 11452
rect 16380 11506 16436 12460
rect 16492 12290 16548 13580
rect 16604 13570 16660 13580
rect 17164 13076 17220 14254
rect 17164 13010 17220 13020
rect 17388 13858 17444 13870
rect 17388 13806 17390 13858
rect 17442 13806 17444 13858
rect 16492 12238 16494 12290
rect 16546 12238 16548 12290
rect 16492 12226 16548 12238
rect 16604 12962 16660 12974
rect 16604 12910 16606 12962
rect 16658 12910 16660 12962
rect 16380 11454 16382 11506
rect 16434 11454 16436 11506
rect 16380 11442 16436 11454
rect 16604 11508 16660 12910
rect 17276 12852 17332 12862
rect 16828 12850 17332 12852
rect 16828 12798 17278 12850
rect 17330 12798 17332 12850
rect 16828 12796 17332 12798
rect 16828 12402 16884 12796
rect 17276 12786 17332 12796
rect 17388 12516 17444 13806
rect 17724 13748 17780 13758
rect 17724 13746 18116 13748
rect 17724 13694 17726 13746
rect 17778 13694 18116 13746
rect 17724 13692 18116 13694
rect 17724 13682 17780 13692
rect 17388 12450 17444 12460
rect 16828 12350 16830 12402
rect 16882 12350 16884 12402
rect 16828 12338 16884 12350
rect 18060 12402 18116 13692
rect 18284 13636 18340 13646
rect 18284 13542 18340 13580
rect 18620 13522 18676 13534
rect 18620 13470 18622 13522
rect 18674 13470 18676 13522
rect 18620 12740 18676 13470
rect 18620 12674 18676 12684
rect 18060 12350 18062 12402
rect 18114 12350 18116 12402
rect 18060 12338 18116 12350
rect 18396 12180 18452 12190
rect 18452 12124 18564 12180
rect 18396 12086 18452 12124
rect 16604 11442 16660 11452
rect 17276 11508 17332 11518
rect 15708 11342 15710 11394
rect 15762 11342 15764 11394
rect 15484 10500 15540 11340
rect 15708 11330 15764 11342
rect 16268 10722 16324 10734
rect 16268 10670 16270 10722
rect 16322 10670 16324 10722
rect 15484 10498 15652 10500
rect 15484 10446 15486 10498
rect 15538 10446 15652 10498
rect 15484 10444 15652 10446
rect 15484 10434 15540 10444
rect 15484 9380 15540 9390
rect 15484 9154 15540 9324
rect 15484 9102 15486 9154
rect 15538 9102 15540 9154
rect 15484 9090 15540 9102
rect 15372 8990 15374 9042
rect 15426 8990 15428 9042
rect 15372 8978 15428 8990
rect 14812 6638 14814 6690
rect 14866 6638 14868 6690
rect 14812 6626 14868 6638
rect 15148 6748 15316 6804
rect 15036 6580 15092 6590
rect 15036 6486 15092 6524
rect 14028 6468 14084 6478
rect 13804 6466 14084 6468
rect 13804 6414 14030 6466
rect 14082 6414 14084 6466
rect 13804 6412 14084 6414
rect 13468 6020 13524 6030
rect 13356 6018 13524 6020
rect 13356 5966 13470 6018
rect 13522 5966 13524 6018
rect 13356 5964 13524 5966
rect 12236 4562 12628 4564
rect 12236 4510 12238 4562
rect 12290 4510 12628 4562
rect 12236 4508 12628 4510
rect 12236 4498 12292 4508
rect 12572 4338 12628 4508
rect 13356 4450 13412 5964
rect 13468 5954 13524 5964
rect 13804 6018 13860 6412
rect 14028 6402 14084 6412
rect 15148 6356 15204 6748
rect 14924 6300 15204 6356
rect 15260 6580 15316 6590
rect 14924 6130 14980 6300
rect 14924 6078 14926 6130
rect 14978 6078 14980 6130
rect 14924 6066 14980 6078
rect 13804 5966 13806 6018
rect 13858 5966 13860 6018
rect 13804 5954 13860 5966
rect 15260 5908 15316 6524
rect 15596 5908 15652 10444
rect 16268 8820 16324 10670
rect 16604 10612 16660 10622
rect 16604 10610 16996 10612
rect 16604 10558 16606 10610
rect 16658 10558 16996 10610
rect 16604 10556 16996 10558
rect 16604 10546 16660 10556
rect 16380 9940 16436 9950
rect 16380 9846 16436 9884
rect 16940 9940 16996 10556
rect 16940 9846 16996 9884
rect 17276 9826 17332 11452
rect 17836 11508 17892 11518
rect 17836 10834 17892 11452
rect 18508 11506 18564 12124
rect 18508 11454 18510 11506
rect 18562 11454 18564 11506
rect 18508 11442 18564 11454
rect 18844 11508 18900 19740
rect 19404 19702 19460 19740
rect 20300 19460 20356 20748
rect 21308 20692 21364 20702
rect 21308 20598 21364 20636
rect 20860 20244 20916 20254
rect 20860 20130 20916 20188
rect 20860 20078 20862 20130
rect 20914 20078 20916 20130
rect 20860 20066 20916 20078
rect 21084 20244 21140 20254
rect 20300 19394 20356 19404
rect 20412 19796 20468 19806
rect 20412 19348 20468 19740
rect 21084 19348 21140 20188
rect 21308 20132 21364 20142
rect 21308 20038 21364 20076
rect 20412 19346 20916 19348
rect 20412 19294 20414 19346
rect 20466 19294 20916 19346
rect 20412 19292 20916 19294
rect 20412 19282 20468 19292
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20860 18562 20916 19292
rect 21084 19282 21140 19292
rect 21308 19234 21364 19246
rect 21308 19182 21310 19234
rect 21362 19182 21364 19234
rect 20860 18510 20862 18562
rect 20914 18510 20916 18562
rect 20860 18498 20916 18510
rect 21196 18676 21252 18686
rect 21196 18452 21252 18620
rect 20972 18450 21252 18452
rect 20972 18398 21198 18450
rect 21250 18398 21252 18450
rect 20972 18396 21252 18398
rect 19516 17554 19572 17566
rect 19516 17502 19518 17554
rect 19570 17502 19572 17554
rect 19180 17444 19236 17454
rect 19068 17442 19236 17444
rect 19068 17390 19182 17442
rect 19234 17390 19236 17442
rect 19068 17388 19236 17390
rect 19068 16994 19124 17388
rect 19180 17378 19236 17388
rect 19068 16942 19070 16994
rect 19122 16942 19124 16994
rect 19068 16930 19124 16942
rect 18956 16772 19012 16782
rect 19012 16716 19124 16772
rect 18956 16706 19012 16716
rect 19068 16100 19124 16716
rect 19516 16322 19572 17502
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19516 16270 19518 16322
rect 19570 16270 19572 16322
rect 19516 16258 19572 16270
rect 19852 16548 19908 16558
rect 19852 16322 19908 16492
rect 19852 16270 19854 16322
rect 19906 16270 19908 16322
rect 19852 16258 19908 16270
rect 20972 16324 21028 18396
rect 21196 18386 21252 18396
rect 21308 18452 21364 19182
rect 21308 18386 21364 18396
rect 21196 18228 21252 18238
rect 21196 18134 21252 18172
rect 21420 18004 21476 21308
rect 21532 20802 21588 21868
rect 21644 21364 21700 21374
rect 21644 21026 21700 21308
rect 21644 20974 21646 21026
rect 21698 20974 21700 21026
rect 21644 20962 21700 20974
rect 21532 20750 21534 20802
rect 21586 20750 21588 20802
rect 21532 20738 21588 20750
rect 21756 20802 21812 23324
rect 21868 22932 21924 23772
rect 21868 22876 22036 22932
rect 21868 22258 21924 22270
rect 21868 22206 21870 22258
rect 21922 22206 21924 22258
rect 21868 21588 21924 22206
rect 21980 21698 22036 22876
rect 21980 21646 21982 21698
rect 22034 21646 22036 21698
rect 21980 21634 22036 21646
rect 21868 21522 21924 21532
rect 22092 21588 22148 24446
rect 22428 24498 22484 24510
rect 22428 24446 22430 24498
rect 22482 24446 22484 24498
rect 22204 23268 22260 23278
rect 22204 23174 22260 23212
rect 22316 21924 22372 21934
rect 22204 21588 22260 21598
rect 22092 21586 22260 21588
rect 22092 21534 22206 21586
rect 22258 21534 22260 21586
rect 22092 21532 22260 21534
rect 22092 21364 22148 21532
rect 22204 21522 22260 21532
rect 22092 21298 22148 21308
rect 21756 20750 21758 20802
rect 21810 20750 21812 20802
rect 21756 20738 21812 20750
rect 22316 20802 22372 21868
rect 22428 21588 22484 24446
rect 23100 24164 23156 24780
rect 22652 24108 23156 24164
rect 22540 23940 22596 23950
rect 22652 23940 22708 24108
rect 22540 23938 22708 23940
rect 22540 23886 22542 23938
rect 22594 23886 22708 23938
rect 22540 23884 22708 23886
rect 23100 23940 23156 23950
rect 22540 23156 22596 23884
rect 23100 23846 23156 23884
rect 22764 23828 22820 23838
rect 22540 23090 22596 23100
rect 22652 23492 22708 23502
rect 22652 23154 22708 23436
rect 22652 23102 22654 23154
rect 22706 23102 22708 23154
rect 22652 23090 22708 23102
rect 22764 22370 22820 23772
rect 22876 23716 22932 23726
rect 22876 23622 22932 23660
rect 22988 23714 23044 23726
rect 22988 23662 22990 23714
rect 23042 23662 23044 23714
rect 22764 22318 22766 22370
rect 22818 22318 22820 22370
rect 22764 22306 22820 22318
rect 22988 21588 23044 23662
rect 23100 23380 23156 23390
rect 23100 23266 23156 23324
rect 23324 23380 23380 25228
rect 23548 24836 23604 24846
rect 23548 24742 23604 24780
rect 23660 24836 23716 24846
rect 23660 24834 23828 24836
rect 23660 24782 23662 24834
rect 23714 24782 23828 24834
rect 23660 24780 23828 24782
rect 23660 24770 23716 24780
rect 23772 24612 23828 24780
rect 24220 24612 24276 24622
rect 23772 24610 24276 24612
rect 23772 24558 24222 24610
rect 24274 24558 24276 24610
rect 23772 24556 24276 24558
rect 23660 24500 23716 24510
rect 23660 24406 23716 24444
rect 23324 23314 23380 23324
rect 23548 24050 23604 24062
rect 23548 23998 23550 24050
rect 23602 23998 23604 24050
rect 23100 23214 23102 23266
rect 23154 23214 23156 23266
rect 23100 23202 23156 23214
rect 23436 23042 23492 23054
rect 23436 22990 23438 23042
rect 23490 22990 23492 23042
rect 23100 22484 23156 22494
rect 23100 22390 23156 22428
rect 23324 22146 23380 22158
rect 23324 22094 23326 22146
rect 23378 22094 23380 22146
rect 23324 21924 23380 22094
rect 23324 21858 23380 21868
rect 23212 21700 23268 21710
rect 23212 21606 23268 21644
rect 22428 21532 22708 21588
rect 22540 21362 22596 21374
rect 22540 21310 22542 21362
rect 22594 21310 22596 21362
rect 22540 20916 22596 21310
rect 22652 21028 22708 21532
rect 22988 21586 23156 21588
rect 22988 21534 22990 21586
rect 23042 21534 23156 21586
rect 22988 21532 23156 21534
rect 22988 21522 23044 21532
rect 22652 20972 23044 21028
rect 22540 20860 22932 20916
rect 22316 20750 22318 20802
rect 22370 20750 22372 20802
rect 22316 20738 22372 20750
rect 21980 20578 22036 20590
rect 21980 20526 21982 20578
rect 22034 20526 22036 20578
rect 21980 20132 22036 20526
rect 22204 20578 22260 20590
rect 22204 20526 22206 20578
rect 22258 20526 22260 20578
rect 22204 20244 22260 20526
rect 22204 20178 22260 20188
rect 22764 20578 22820 20590
rect 22764 20526 22766 20578
rect 22818 20526 22820 20578
rect 22764 20244 22820 20526
rect 22764 20178 22820 20188
rect 21980 20066 22036 20076
rect 22428 20132 22484 20142
rect 22428 20038 22484 20076
rect 21756 20020 21812 20030
rect 21644 19794 21700 19806
rect 21644 19742 21646 19794
rect 21698 19742 21700 19794
rect 21644 19348 21700 19742
rect 21644 19282 21700 19292
rect 21644 18452 21700 18462
rect 20636 16212 20692 16222
rect 20524 16156 20636 16212
rect 19068 16098 19460 16100
rect 19068 16046 19070 16098
rect 19122 16046 19460 16098
rect 19068 16044 19460 16046
rect 19068 16034 19124 16044
rect 18956 15988 19012 15998
rect 18956 12290 19012 15932
rect 19180 15764 19236 15774
rect 19180 15428 19236 15708
rect 19404 15538 19460 16044
rect 20524 16098 20580 16156
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 20524 16034 20580 16046
rect 20412 15988 20468 15998
rect 20412 15894 20468 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19404 15486 19406 15538
rect 19458 15486 19460 15538
rect 19404 15474 19460 15486
rect 19180 13858 19236 15372
rect 20076 15426 20132 15438
rect 20076 15374 20078 15426
rect 20130 15374 20132 15426
rect 19852 15316 19908 15326
rect 19852 15222 19908 15260
rect 20076 14644 20132 15374
rect 20524 15428 20580 15438
rect 20524 15334 20580 15372
rect 20636 15314 20692 16156
rect 20636 15262 20638 15314
rect 20690 15262 20692 15314
rect 20636 15250 20692 15262
rect 20972 15148 21028 16268
rect 20076 14578 20132 14588
rect 20860 15092 21028 15148
rect 21084 17948 21476 18004
rect 21532 18396 21644 18452
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19180 13806 19182 13858
rect 19234 13806 19236 13858
rect 19180 13794 19236 13806
rect 19516 13804 19796 13860
rect 19404 13748 19460 13758
rect 19516 13748 19572 13804
rect 18956 12238 18958 12290
rect 19010 12238 19012 12290
rect 18956 12226 19012 12238
rect 19292 13746 19572 13748
rect 19292 13694 19406 13746
rect 19458 13694 19572 13746
rect 19292 13692 19572 13694
rect 19180 12180 19236 12190
rect 19292 12180 19348 13692
rect 19404 13682 19460 13692
rect 19628 13636 19684 13646
rect 19404 13074 19460 13086
rect 19404 13022 19406 13074
rect 19458 13022 19460 13074
rect 19404 12740 19460 13022
rect 19404 12674 19460 12684
rect 19180 12178 19348 12180
rect 19180 12126 19182 12178
rect 19234 12126 19348 12178
rect 19180 12124 19348 12126
rect 19180 12114 19236 12124
rect 19628 12068 19684 13580
rect 19740 13186 19796 13804
rect 20860 13746 20916 15092
rect 20860 13694 20862 13746
rect 20914 13694 20916 13746
rect 20860 13682 20916 13694
rect 19740 13134 19742 13186
rect 19794 13134 19796 13186
rect 19740 13122 19796 13134
rect 20524 13522 20580 13534
rect 20524 13470 20526 13522
rect 20578 13470 20580 13522
rect 20076 12964 20132 12974
rect 20076 12962 20244 12964
rect 20076 12910 20078 12962
rect 20130 12910 20244 12962
rect 20076 12908 20244 12910
rect 20076 12898 20132 12908
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19740 12068 19796 12078
rect 19628 12066 20020 12068
rect 19628 12014 19742 12066
rect 19794 12014 20020 12066
rect 19628 12012 20020 12014
rect 19740 12002 19796 12012
rect 19292 11956 19348 11966
rect 18844 11452 19236 11508
rect 19068 11170 19124 11182
rect 19068 11118 19070 11170
rect 19122 11118 19124 11170
rect 17836 10782 17838 10834
rect 17890 10782 17892 10834
rect 17836 10770 17892 10782
rect 18956 10836 19012 10846
rect 18172 10724 18228 10734
rect 17948 10722 18228 10724
rect 17948 10670 18174 10722
rect 18226 10670 18228 10722
rect 17948 10668 18228 10670
rect 17948 9938 18004 10668
rect 18172 10658 18228 10668
rect 17948 9886 17950 9938
rect 18002 9886 18004 9938
rect 17948 9874 18004 9886
rect 18396 10610 18452 10622
rect 18396 10558 18398 10610
rect 18450 10558 18452 10610
rect 17276 9774 17278 9826
rect 17330 9774 17332 9826
rect 17276 9762 17332 9774
rect 18396 9266 18452 10558
rect 18396 9214 18398 9266
rect 18450 9214 18452 9266
rect 18396 9202 18452 9214
rect 18956 9154 19012 10780
rect 19068 10610 19124 11118
rect 19068 10558 19070 10610
rect 19122 10558 19124 10610
rect 19068 10276 19124 10558
rect 19068 10210 19124 10220
rect 18956 9102 18958 9154
rect 19010 9102 19012 9154
rect 18956 9090 19012 9102
rect 16268 8754 16324 8764
rect 18060 8820 18116 8830
rect 17836 8260 17892 8270
rect 17724 8148 17780 8158
rect 17724 8054 17780 8092
rect 16492 7586 16548 7598
rect 16492 7534 16494 7586
rect 16546 7534 16548 7586
rect 16380 6804 16436 6814
rect 16492 6804 16548 7534
rect 16828 7476 16884 7486
rect 16828 7382 16884 7420
rect 17500 7476 17556 7486
rect 17500 7382 17556 7420
rect 17836 7476 17892 8204
rect 17836 7382 17892 7420
rect 16380 6802 16548 6804
rect 16380 6750 16382 6802
rect 16434 6750 16548 6802
rect 16380 6748 16548 6750
rect 16380 6738 16436 6748
rect 15708 6692 15764 6702
rect 15708 6598 15764 6636
rect 16604 6692 16660 6702
rect 16044 6020 16100 6030
rect 16044 5926 16100 5964
rect 15932 5908 15988 5918
rect 15260 5906 15540 5908
rect 15260 5854 15262 5906
rect 15314 5854 15540 5906
rect 15260 5852 15540 5854
rect 15596 5906 15988 5908
rect 15596 5854 15934 5906
rect 15986 5854 15988 5906
rect 15596 5852 15988 5854
rect 15260 5842 15316 5852
rect 13356 4398 13358 4450
rect 13410 4398 13412 4450
rect 13356 4386 13412 4398
rect 12572 4286 12574 4338
rect 12626 4286 12628 4338
rect 12572 4274 12628 4286
rect 15484 4226 15540 5852
rect 15932 5236 15988 5852
rect 16492 5908 16548 5918
rect 16492 5814 16548 5852
rect 16268 5236 16324 5246
rect 15932 5234 16324 5236
rect 15932 5182 16270 5234
rect 16322 5182 16324 5234
rect 15932 5180 16324 5182
rect 16268 5170 16324 5180
rect 16604 5122 16660 6636
rect 16828 6020 16884 6030
rect 16828 6018 17332 6020
rect 16828 5966 16830 6018
rect 16882 5966 17332 6018
rect 16828 5964 17332 5966
rect 16828 5954 16884 5964
rect 17276 5234 17332 5964
rect 17612 5908 17668 5918
rect 17612 5814 17668 5852
rect 17948 5908 18004 5918
rect 18060 5908 18116 8764
rect 18732 8820 18788 8830
rect 18732 8726 18788 8764
rect 18284 8260 18340 8270
rect 18284 8166 18340 8204
rect 18508 8258 18564 8270
rect 18508 8206 18510 8258
rect 18562 8206 18564 8258
rect 18508 8036 18564 8206
rect 19180 8260 19236 11452
rect 19292 10498 19348 11900
rect 19852 11620 19908 11630
rect 19292 10446 19294 10498
rect 19346 10446 19348 10498
rect 19292 8932 19348 10446
rect 19292 8866 19348 8876
rect 19404 11618 19908 11620
rect 19404 11566 19854 11618
rect 19906 11566 19908 11618
rect 19404 11564 19908 11566
rect 19180 8166 19236 8204
rect 18508 7970 18564 7980
rect 18844 8146 18900 8158
rect 18844 8094 18846 8146
rect 18898 8094 18900 8146
rect 18844 7812 18900 8094
rect 18396 7756 18900 7812
rect 19180 8036 19236 8046
rect 18284 7476 18340 7486
rect 18396 7476 18452 7756
rect 19180 7700 19236 7980
rect 19180 7606 19236 7644
rect 18284 7474 18452 7476
rect 18284 7422 18286 7474
rect 18338 7422 18452 7474
rect 18284 7420 18452 7422
rect 18508 7588 18564 7598
rect 18284 6018 18340 7420
rect 18508 6802 18564 7532
rect 19404 7476 19460 11564
rect 19852 11554 19908 11564
rect 19964 11508 20020 12012
rect 20076 11956 20132 11966
rect 20188 11956 20244 12908
rect 20132 11900 20244 11956
rect 20300 12850 20356 12862
rect 20300 12798 20302 12850
rect 20354 12798 20356 12850
rect 20076 11890 20132 11900
rect 20300 11844 20356 12798
rect 20524 12180 20580 13470
rect 20860 13522 20916 13534
rect 20860 13470 20862 13522
rect 20914 13470 20916 13522
rect 20860 13188 20916 13470
rect 20860 13122 20916 13132
rect 20524 12114 20580 12124
rect 20748 12740 20804 12750
rect 21084 12740 21140 17948
rect 21532 16996 21588 18396
rect 21644 18358 21700 18396
rect 21644 17332 21700 17342
rect 21644 17106 21700 17276
rect 21644 17054 21646 17106
rect 21698 17054 21700 17106
rect 21644 17042 21700 17054
rect 21420 16882 21476 16894
rect 21420 16830 21422 16882
rect 21474 16830 21476 16882
rect 21196 16770 21252 16782
rect 21196 16718 21198 16770
rect 21250 16718 21252 16770
rect 21196 16548 21252 16718
rect 21196 16482 21252 16492
rect 21420 16212 21476 16830
rect 21420 16146 21476 16156
rect 21532 16210 21588 16940
rect 21756 16994 21812 19964
rect 22652 20018 22708 20030
rect 22652 19966 22654 20018
rect 22706 19966 22708 20018
rect 21980 19908 22036 19918
rect 21980 19814 22036 19852
rect 22652 19908 22708 19966
rect 22652 19842 22708 19852
rect 22204 19572 22260 19582
rect 22092 19124 22148 19134
rect 22092 19030 22148 19068
rect 21980 18116 22036 18126
rect 21980 17332 22036 18060
rect 21756 16942 21758 16994
rect 21810 16942 21812 16994
rect 21756 16930 21812 16942
rect 21868 17108 21924 17118
rect 21532 16158 21534 16210
rect 21586 16158 21588 16210
rect 21532 16146 21588 16158
rect 21644 15316 21700 15326
rect 21644 15222 21700 15260
rect 21308 15090 21364 15102
rect 21308 15038 21310 15090
rect 21362 15038 21364 15090
rect 21308 14532 21364 15038
rect 21308 14466 21364 14476
rect 21420 14530 21476 14542
rect 21420 14478 21422 14530
rect 21474 14478 21476 14530
rect 21196 13746 21252 13758
rect 21196 13694 21198 13746
rect 21250 13694 21252 13746
rect 21196 13524 21252 13694
rect 21420 13636 21476 14478
rect 21420 13570 21476 13580
rect 21196 13458 21252 13468
rect 21868 13524 21924 17052
rect 21980 15874 22036 17276
rect 21980 15822 21982 15874
rect 22034 15822 22036 15874
rect 21980 15204 22036 15822
rect 21980 15138 22036 15148
rect 22092 14644 22148 14654
rect 22092 14550 22148 14588
rect 21868 13458 21924 13468
rect 21868 13300 21924 13310
rect 20748 12738 21140 12740
rect 20748 12686 20750 12738
rect 20802 12686 21140 12738
rect 20748 12684 21140 12686
rect 21644 12850 21700 12862
rect 21644 12798 21646 12850
rect 21698 12798 21700 12850
rect 20748 11956 20804 12684
rect 21644 12402 21700 12798
rect 21644 12350 21646 12402
rect 21698 12350 21700 12402
rect 21644 12338 21700 12350
rect 20748 11890 20804 11900
rect 21532 12066 21588 12078
rect 21532 12014 21534 12066
rect 21586 12014 21588 12066
rect 20300 11778 20356 11788
rect 20020 11452 20132 11508
rect 19964 11442 20020 11452
rect 20076 11396 20132 11452
rect 20076 11340 20244 11396
rect 19516 11170 19572 11182
rect 19516 11118 19518 11170
rect 19570 11118 19572 11170
rect 19516 10612 19572 11118
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10836 20244 11340
rect 20076 10780 20244 10836
rect 19516 10556 19684 10612
rect 19628 9828 19684 10556
rect 20076 10610 20132 10780
rect 20076 10558 20078 10610
rect 20130 10558 20132 10610
rect 20076 10546 20132 10558
rect 19628 9762 19684 9772
rect 20076 10388 20132 10398
rect 20076 9938 20132 10332
rect 20076 9886 20078 9938
rect 20130 9886 20132 9938
rect 20076 9604 20132 9886
rect 19516 9548 20132 9604
rect 20188 10052 20244 10780
rect 20300 11394 20356 11406
rect 20300 11342 20302 11394
rect 20354 11342 20356 11394
rect 20300 10836 20356 11342
rect 20636 11284 20692 11294
rect 20636 11190 20692 11228
rect 20300 10770 20356 10780
rect 19516 9154 19572 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9380 20244 9996
rect 20748 10498 20804 10510
rect 20748 10446 20750 10498
rect 20802 10446 20804 10498
rect 20412 9828 20468 9838
rect 20412 9734 20468 9772
rect 20748 9714 20804 10446
rect 21532 10388 21588 12014
rect 21532 10322 21588 10332
rect 20748 9662 20750 9714
rect 20802 9662 20804 9714
rect 20748 9650 20804 9662
rect 20188 9324 20580 9380
rect 19516 9102 19518 9154
rect 19570 9102 19572 9154
rect 19516 9090 19572 9102
rect 20076 8932 20132 8942
rect 20076 8838 20132 8876
rect 19628 8260 19684 8270
rect 20076 8260 20132 8270
rect 19628 8258 20132 8260
rect 19628 8206 19630 8258
rect 19682 8206 20078 8258
rect 20130 8206 20132 8258
rect 19628 8204 20132 8206
rect 19628 8194 19684 8204
rect 20076 8036 20132 8204
rect 20076 7970 20132 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19404 7410 19460 7420
rect 20300 7474 20356 9324
rect 20524 9266 20580 9324
rect 20524 9214 20526 9266
rect 20578 9214 20580 9266
rect 20524 9202 20580 9214
rect 21308 8932 21364 8942
rect 21308 8838 21364 8876
rect 21756 8930 21812 8942
rect 21756 8878 21758 8930
rect 21810 8878 21812 8930
rect 20412 8820 20468 8830
rect 20412 8258 20468 8764
rect 21756 8484 21812 8878
rect 21756 8418 21812 8428
rect 20412 8206 20414 8258
rect 20466 8206 20468 8258
rect 20412 8194 20468 8206
rect 21868 8258 21924 13244
rect 22092 13188 22148 13198
rect 22092 13094 22148 13132
rect 21980 12962 22036 12974
rect 21980 12910 21982 12962
rect 22034 12910 22036 12962
rect 21980 12628 22036 12910
rect 21980 12562 22036 12572
rect 22092 11732 22148 11742
rect 22204 11732 22260 19516
rect 22652 17108 22708 17118
rect 22652 16882 22708 17052
rect 22652 16830 22654 16882
rect 22706 16830 22708 16882
rect 22652 16818 22708 16830
rect 22764 16436 22820 16446
rect 22764 16098 22820 16380
rect 22764 16046 22766 16098
rect 22818 16046 22820 16098
rect 22764 16034 22820 16046
rect 22876 14644 22932 20860
rect 22988 20132 23044 20972
rect 23100 20692 23156 21532
rect 23324 21140 23380 21150
rect 23324 21026 23380 21084
rect 23324 20974 23326 21026
rect 23378 20974 23380 21026
rect 23324 20962 23380 20974
rect 23212 20692 23268 20702
rect 23100 20690 23268 20692
rect 23100 20638 23214 20690
rect 23266 20638 23268 20690
rect 23100 20636 23268 20638
rect 23212 20626 23268 20636
rect 23436 20356 23492 22990
rect 23548 21586 23604 23998
rect 24220 23940 24276 24556
rect 24220 23874 24276 23884
rect 23996 23826 24052 23838
rect 23996 23774 23998 23826
rect 24050 23774 24052 23826
rect 23996 23492 24052 23774
rect 24444 23716 24500 25564
rect 24892 25506 24948 26012
rect 24892 25454 24894 25506
rect 24946 25454 24948 25506
rect 24892 25442 24948 25454
rect 24668 24948 24724 24958
rect 24668 24854 24724 24892
rect 24052 23436 24388 23492
rect 23996 23426 24052 23436
rect 24332 23266 24388 23436
rect 24444 23378 24500 23660
rect 24444 23326 24446 23378
rect 24498 23326 24500 23378
rect 24444 23314 24500 23326
rect 24556 24836 24612 24846
rect 24332 23214 24334 23266
rect 24386 23214 24388 23266
rect 24332 23202 24388 23214
rect 23996 22596 24052 22606
rect 23996 21700 24052 22540
rect 24444 22596 24500 22606
rect 24444 22482 24500 22540
rect 24444 22430 24446 22482
rect 24498 22430 24500 22482
rect 24444 22418 24500 22430
rect 24556 22372 24612 24780
rect 24892 23940 24948 23950
rect 24892 23846 24948 23884
rect 24668 23156 24724 23166
rect 24668 23154 24948 23156
rect 24668 23102 24670 23154
rect 24722 23102 24948 23154
rect 24668 23100 24948 23102
rect 24668 23090 24724 23100
rect 24892 22482 24948 23100
rect 24892 22430 24894 22482
rect 24946 22430 24948 22482
rect 24780 22372 24836 22382
rect 24556 22370 24836 22372
rect 24556 22318 24782 22370
rect 24834 22318 24836 22370
rect 24556 22316 24836 22318
rect 24780 22306 24836 22316
rect 24556 21812 24612 21822
rect 23996 21698 24276 21700
rect 23996 21646 23998 21698
rect 24050 21646 24276 21698
rect 23996 21644 24276 21646
rect 23996 21634 24052 21644
rect 23548 21534 23550 21586
rect 23602 21534 23604 21586
rect 23548 20580 23604 21534
rect 23660 21362 23716 21374
rect 23660 21310 23662 21362
rect 23714 21310 23716 21362
rect 23660 20804 23716 21310
rect 24220 20914 24276 21644
rect 24556 21588 24612 21756
rect 24668 21700 24724 21710
rect 24668 21606 24724 21644
rect 24220 20862 24222 20914
rect 24274 20862 24276 20914
rect 24220 20850 24276 20862
rect 24332 21586 24612 21588
rect 24332 21534 24558 21586
rect 24610 21534 24612 21586
rect 24332 21532 24612 21534
rect 23660 20748 23940 20804
rect 23772 20580 23828 20590
rect 23548 20578 23828 20580
rect 23548 20526 23774 20578
rect 23826 20526 23828 20578
rect 23548 20524 23828 20526
rect 23436 20290 23492 20300
rect 23212 20244 23268 20254
rect 23212 20150 23268 20188
rect 23100 20132 23156 20142
rect 22988 20130 23156 20132
rect 22988 20078 23102 20130
rect 23154 20078 23156 20130
rect 22988 20076 23156 20078
rect 22988 20020 23044 20076
rect 23100 20066 23156 20076
rect 22988 19954 23044 19964
rect 23436 20020 23492 20030
rect 23436 19926 23492 19964
rect 23212 17892 23268 17902
rect 23212 17666 23268 17836
rect 23212 17614 23214 17666
rect 23266 17614 23268 17666
rect 23212 17602 23268 17614
rect 23548 17556 23604 17566
rect 23548 17462 23604 17500
rect 23660 17332 23716 20524
rect 23772 20514 23828 20524
rect 23772 20132 23828 20142
rect 23772 20038 23828 20076
rect 23548 17276 23716 17332
rect 23772 18340 23828 18350
rect 23884 18340 23940 20748
rect 24220 19348 24276 19358
rect 24220 18788 24276 19292
rect 24220 18722 24276 18732
rect 24332 18450 24388 21532
rect 24556 21522 24612 21532
rect 24892 21588 24948 22430
rect 24892 21522 24948 21532
rect 25004 20914 25060 26852
rect 25116 26292 25172 26302
rect 25116 26198 25172 26236
rect 25452 26290 25508 28588
rect 25564 29314 25620 29326
rect 25564 29262 25566 29314
rect 25618 29262 25620 29314
rect 25564 27746 25620 29262
rect 26460 28868 26516 31502
rect 26572 31556 26628 37100
rect 26684 37090 26740 37100
rect 26908 37044 26964 39900
rect 27244 39842 27300 40236
rect 27244 39790 27246 39842
rect 27298 39790 27300 39842
rect 27244 39778 27300 39790
rect 27692 39618 27748 39630
rect 27692 39566 27694 39618
rect 27746 39566 27748 39618
rect 27692 39060 27748 39566
rect 27916 39620 27972 39630
rect 27916 39526 27972 39564
rect 28140 39508 28196 40348
rect 28252 40068 28308 42476
rect 28364 42420 28420 43708
rect 28476 43540 28532 43550
rect 28476 43446 28532 43484
rect 28700 43538 28756 43550
rect 28700 43486 28702 43538
rect 28754 43486 28756 43538
rect 28700 43428 28756 43486
rect 28924 43540 28980 43550
rect 28924 43446 28980 43484
rect 28588 43204 28644 43214
rect 28588 42754 28644 43148
rect 28588 42702 28590 42754
rect 28642 42702 28644 42754
rect 28588 42690 28644 42702
rect 28476 42644 28532 42654
rect 28476 42550 28532 42588
rect 28364 42354 28420 42364
rect 28364 42196 28420 42206
rect 28364 42102 28420 42140
rect 28588 42196 28644 42206
rect 28700 42196 28756 43372
rect 28812 43316 28868 43326
rect 28812 43222 28868 43260
rect 29036 43092 29092 44044
rect 29596 43650 29652 44270
rect 29820 44322 29876 45052
rect 30044 45106 30100 45164
rect 30044 45054 30046 45106
rect 30098 45054 30100 45106
rect 30044 45042 30100 45054
rect 30268 44436 30324 45724
rect 30716 45714 30772 45724
rect 30716 45556 30772 45566
rect 30716 45106 30772 45500
rect 30716 45054 30718 45106
rect 30770 45054 30772 45106
rect 30716 45042 30772 45054
rect 30940 45108 30996 45118
rect 29820 44270 29822 44322
rect 29874 44270 29876 44322
rect 29820 44258 29876 44270
rect 30044 44380 30324 44436
rect 30940 44434 30996 45052
rect 30940 44382 30942 44434
rect 30994 44382 30996 44434
rect 30044 44322 30100 44380
rect 30940 44370 30996 44382
rect 30380 44324 30436 44334
rect 30044 44270 30046 44322
rect 30098 44270 30100 44322
rect 30044 44258 30100 44270
rect 30268 44322 30436 44324
rect 30268 44270 30382 44322
rect 30434 44270 30436 44322
rect 30268 44268 30436 44270
rect 31052 44324 31108 45724
rect 31164 45780 31220 46172
rect 31276 45892 31332 46620
rect 31724 46676 31780 46686
rect 31948 46676 32004 46956
rect 32508 46946 32564 46956
rect 31724 46674 32004 46676
rect 31724 46622 31726 46674
rect 31778 46622 32004 46674
rect 31724 46620 32004 46622
rect 32060 46786 32116 46798
rect 32060 46734 32062 46786
rect 32114 46734 32116 46786
rect 32060 46676 32116 46734
rect 32396 46788 32452 46798
rect 32396 46694 32452 46732
rect 31724 46564 31780 46620
rect 32060 46610 32116 46620
rect 31724 46498 31780 46508
rect 32508 46450 32564 46462
rect 32508 46398 32510 46450
rect 32562 46398 32564 46450
rect 31388 46114 31444 46126
rect 31388 46062 31390 46114
rect 31442 46062 31444 46114
rect 31388 46004 31444 46062
rect 31836 46004 31892 46014
rect 31388 46002 31892 46004
rect 31388 45950 31838 46002
rect 31890 45950 31892 46002
rect 31388 45948 31892 45950
rect 31836 45938 31892 45948
rect 32060 45892 32116 45902
rect 32508 45892 32564 46398
rect 31276 45836 31444 45892
rect 31164 45714 31220 45724
rect 31276 45666 31332 45678
rect 31276 45614 31278 45666
rect 31330 45614 31332 45666
rect 31276 45332 31332 45614
rect 31276 45266 31332 45276
rect 31388 45220 31444 45836
rect 32060 45890 32564 45892
rect 32060 45838 32062 45890
rect 32114 45838 32510 45890
rect 32562 45838 32564 45890
rect 32060 45836 32564 45838
rect 32060 45826 32116 45836
rect 32508 45826 32564 45836
rect 31724 45780 31780 45790
rect 31724 45686 31780 45724
rect 31388 45126 31444 45164
rect 31948 45388 32452 45444
rect 31276 45106 31332 45118
rect 31276 45054 31278 45106
rect 31330 45054 31332 45106
rect 31276 44548 31332 45054
rect 31276 44482 31332 44492
rect 31388 44994 31444 45006
rect 31388 44942 31390 44994
rect 31442 44942 31444 44994
rect 31276 44324 31332 44334
rect 31052 44268 31220 44324
rect 29932 44100 29988 44110
rect 29932 44006 29988 44044
rect 30044 43988 30100 43998
rect 29596 43598 29598 43650
rect 29650 43598 29652 43650
rect 29596 43316 29652 43598
rect 29708 43652 29764 43662
rect 29708 43538 29764 43596
rect 29708 43486 29710 43538
rect 29762 43486 29764 43538
rect 29708 43474 29764 43486
rect 29596 43260 29876 43316
rect 28588 42194 28756 42196
rect 28588 42142 28590 42194
rect 28642 42142 28756 42194
rect 28588 42140 28756 42142
rect 28812 43036 29092 43092
rect 28588 42130 28644 42140
rect 28812 41970 28868 43036
rect 29148 42868 29204 42878
rect 29148 42774 29204 42812
rect 29484 42866 29540 42878
rect 29484 42814 29486 42866
rect 29538 42814 29540 42866
rect 29484 42756 29540 42814
rect 29484 42690 29540 42700
rect 29708 42868 29764 42878
rect 29372 42530 29428 42542
rect 29372 42478 29374 42530
rect 29426 42478 29428 42530
rect 29036 41972 29092 41982
rect 28812 41918 28814 41970
rect 28866 41918 28868 41970
rect 28812 41906 28868 41918
rect 28924 41970 29092 41972
rect 28924 41918 29038 41970
rect 29090 41918 29092 41970
rect 28924 41916 29092 41918
rect 28588 41748 28644 41758
rect 28588 40964 28644 41692
rect 28700 41748 28756 41758
rect 28924 41748 28980 41916
rect 29036 41906 29092 41916
rect 29372 41972 29428 42478
rect 29708 42194 29764 42812
rect 29820 42756 29876 43260
rect 30044 42978 30100 43932
rect 30044 42926 30046 42978
rect 30098 42926 30100 42978
rect 30044 42914 30100 42926
rect 30156 43876 30212 43886
rect 29932 42756 29988 42766
rect 29820 42754 29988 42756
rect 29820 42702 29934 42754
rect 29986 42702 29988 42754
rect 29820 42700 29988 42702
rect 29932 42420 29988 42700
rect 29932 42354 29988 42364
rect 29708 42142 29710 42194
rect 29762 42142 29764 42194
rect 29708 42130 29764 42142
rect 29484 41972 29540 41982
rect 29372 41970 29540 41972
rect 29372 41918 29486 41970
rect 29538 41918 29540 41970
rect 29372 41916 29540 41918
rect 28700 41746 28980 41748
rect 28700 41694 28702 41746
rect 28754 41694 28980 41746
rect 28700 41692 28980 41694
rect 28700 41682 28756 41692
rect 28588 40628 28644 40908
rect 29148 40962 29204 40974
rect 29148 40910 29150 40962
rect 29202 40910 29204 40962
rect 28700 40628 28756 40638
rect 28588 40626 28756 40628
rect 28588 40574 28702 40626
rect 28754 40574 28756 40626
rect 28588 40572 28756 40574
rect 28700 40562 28756 40572
rect 28364 40514 28420 40526
rect 29036 40516 29092 40526
rect 28364 40462 28366 40514
rect 28418 40462 28420 40514
rect 28364 40292 28420 40462
rect 28364 40226 28420 40236
rect 28924 40514 29092 40516
rect 28924 40462 29038 40514
rect 29090 40462 29092 40514
rect 28924 40460 29092 40462
rect 28924 40068 28980 40460
rect 29036 40450 29092 40460
rect 29148 40404 29204 40910
rect 29148 40338 29204 40348
rect 29260 40962 29316 40974
rect 29260 40910 29262 40962
rect 29314 40910 29316 40962
rect 28252 40012 28420 40068
rect 28252 39508 28308 39518
rect 28140 39452 28252 39508
rect 28252 39414 28308 39452
rect 27692 38994 27748 39004
rect 27692 38722 27748 38734
rect 27692 38670 27694 38722
rect 27746 38670 27748 38722
rect 27692 38668 27748 38670
rect 28364 38668 28420 40012
rect 28924 40002 28980 40012
rect 29036 40180 29092 40190
rect 28588 39844 28644 39882
rect 28588 39778 28644 39788
rect 28924 39844 28980 39854
rect 28588 39620 28644 39630
rect 28588 39526 28644 39564
rect 28924 38946 28980 39788
rect 29036 39618 29092 40124
rect 29036 39566 29038 39618
rect 29090 39566 29092 39618
rect 29036 39554 29092 39566
rect 29148 40068 29204 40078
rect 29036 39060 29092 39070
rect 29036 38966 29092 39004
rect 28924 38894 28926 38946
rect 28978 38894 28980 38946
rect 28924 38882 28980 38894
rect 27244 38612 27748 38668
rect 28252 38612 28420 38668
rect 27020 38276 27076 38286
rect 27020 38182 27076 38220
rect 27244 37828 27300 38612
rect 27916 38388 27972 38398
rect 27356 38164 27412 38174
rect 27356 38162 27860 38164
rect 27356 38110 27358 38162
rect 27410 38110 27860 38162
rect 27356 38108 27860 38110
rect 27356 38098 27412 38108
rect 27244 37826 27524 37828
rect 27244 37774 27246 37826
rect 27298 37774 27524 37826
rect 27244 37772 27524 37774
rect 27244 37762 27300 37772
rect 27244 37268 27300 37278
rect 27244 37174 27300 37212
rect 26908 36978 26964 36988
rect 27356 36596 27412 36606
rect 27356 36482 27412 36540
rect 27356 36430 27358 36482
rect 27410 36430 27412 36482
rect 27356 36418 27412 36430
rect 27468 36372 27524 37772
rect 27804 37380 27860 38108
rect 27916 38162 27972 38332
rect 27916 38110 27918 38162
rect 27970 38110 27972 38162
rect 27916 38098 27972 38110
rect 28252 37826 28308 38612
rect 28476 38388 28532 38398
rect 28532 38332 28644 38388
rect 28476 38322 28532 38332
rect 28588 38052 28644 38332
rect 28588 37958 28644 37996
rect 28252 37774 28254 37826
rect 28306 37774 28308 37826
rect 27916 37380 27972 37390
rect 27804 37378 27972 37380
rect 27804 37326 27918 37378
rect 27970 37326 27972 37378
rect 27804 37324 27972 37326
rect 27916 37314 27972 37324
rect 28028 36932 28084 36942
rect 27692 36372 27748 36382
rect 27468 36316 27692 36372
rect 27020 34914 27076 34926
rect 27020 34862 27022 34914
rect 27074 34862 27076 34914
rect 27020 34804 27076 34862
rect 27020 34738 27076 34748
rect 27132 34692 27188 34702
rect 27132 34242 27188 34636
rect 27468 34356 27524 36316
rect 27692 36278 27748 36316
rect 28028 35922 28084 36876
rect 28140 36596 28196 36606
rect 28252 36596 28308 37774
rect 28196 36540 28308 36596
rect 28588 36596 28644 36606
rect 28140 36502 28196 36540
rect 28588 36502 28644 36540
rect 28028 35870 28030 35922
rect 28082 35870 28084 35922
rect 28028 35858 28084 35870
rect 28812 35924 28868 35934
rect 29148 35924 29204 40012
rect 29260 39620 29316 40910
rect 29372 40962 29428 41916
rect 29484 41906 29540 41916
rect 30044 41970 30100 41982
rect 30044 41918 30046 41970
rect 30098 41918 30100 41970
rect 29596 41860 29652 41870
rect 29596 41766 29652 41804
rect 30044 41748 30100 41918
rect 30044 41682 30100 41692
rect 30156 41524 30212 43820
rect 30268 43540 30324 44268
rect 30380 44258 30436 44268
rect 30828 44100 30884 44110
rect 30716 44098 30884 44100
rect 30716 44046 30830 44098
rect 30882 44046 30884 44098
rect 30716 44044 30884 44046
rect 30604 43764 30660 43774
rect 30268 41636 30324 43484
rect 30268 41570 30324 41580
rect 30380 43538 30436 43550
rect 30380 43486 30382 43538
rect 30434 43486 30436 43538
rect 30380 42530 30436 43486
rect 30380 42478 30382 42530
rect 30434 42478 30436 42530
rect 30380 42082 30436 42478
rect 30380 42030 30382 42082
rect 30434 42030 30436 42082
rect 30380 41972 30436 42030
rect 29708 41468 30212 41524
rect 29484 41076 29540 41086
rect 29484 40982 29540 41020
rect 29372 40910 29374 40962
rect 29426 40910 29428 40962
rect 29372 40852 29428 40910
rect 29372 40796 29652 40852
rect 29372 40404 29428 40414
rect 29372 39732 29428 40348
rect 29596 40292 29652 40796
rect 29708 40626 29764 41468
rect 29932 41188 29988 41198
rect 30380 41188 30436 41916
rect 29932 41186 30436 41188
rect 29932 41134 29934 41186
rect 29986 41134 30436 41186
rect 29932 41132 30436 41134
rect 30492 43426 30548 43438
rect 30492 43374 30494 43426
rect 30546 43374 30548 43426
rect 29932 41122 29988 41132
rect 30268 40964 30324 40974
rect 30268 40870 30324 40908
rect 29708 40574 29710 40626
rect 29762 40574 29764 40626
rect 29708 40562 29764 40574
rect 29932 40404 29988 40414
rect 29932 40402 30100 40404
rect 29932 40350 29934 40402
rect 29986 40350 30100 40402
rect 29932 40348 30100 40350
rect 29932 40338 29988 40348
rect 29596 39844 29652 40236
rect 29820 40292 29876 40302
rect 29820 40198 29876 40236
rect 29932 39844 29988 39854
rect 29596 39842 29988 39844
rect 29596 39790 29934 39842
rect 29986 39790 29988 39842
rect 29596 39788 29988 39790
rect 29932 39778 29988 39788
rect 29372 39676 29652 39732
rect 29260 39564 29540 39620
rect 29372 39394 29428 39406
rect 29372 39342 29374 39394
rect 29426 39342 29428 39394
rect 29260 39060 29316 39070
rect 29372 39060 29428 39342
rect 29260 39058 29428 39060
rect 29260 39006 29262 39058
rect 29314 39006 29428 39058
rect 29260 39004 29428 39006
rect 29260 38994 29316 39004
rect 29484 38668 29540 39564
rect 29596 39506 29652 39676
rect 30044 39730 30100 40348
rect 30044 39678 30046 39730
rect 30098 39678 30100 39730
rect 30044 39666 30100 39678
rect 29596 39454 29598 39506
rect 29650 39454 29652 39506
rect 29596 39442 29652 39454
rect 29708 39396 29764 39406
rect 29708 39302 29764 39340
rect 30156 39394 30212 39406
rect 30156 39342 30158 39394
rect 30210 39342 30212 39394
rect 30156 39060 30212 39342
rect 30156 38994 30212 39004
rect 30492 38668 30548 43374
rect 30604 42754 30660 43708
rect 30604 42702 30606 42754
rect 30658 42702 30660 42754
rect 30604 42690 30660 42702
rect 30604 41636 30660 41646
rect 30604 41074 30660 41580
rect 30716 41412 30772 44044
rect 30828 44034 30884 44044
rect 31052 44100 31108 44110
rect 31052 44006 31108 44044
rect 31164 43876 31220 44268
rect 31276 44230 31332 44268
rect 31052 43820 31220 43876
rect 31052 43540 31108 43820
rect 30828 43538 31108 43540
rect 30828 43486 31054 43538
rect 31106 43486 31108 43538
rect 30828 43484 31108 43486
rect 30828 42754 30884 43484
rect 31052 43474 31108 43484
rect 31164 43540 31220 43550
rect 31388 43540 31444 44942
rect 31612 44660 31668 44670
rect 31612 44322 31668 44604
rect 31612 44270 31614 44322
rect 31666 44270 31668 44322
rect 31612 44258 31668 44270
rect 31948 44322 32004 45388
rect 32284 45220 32340 45230
rect 32396 45220 32452 45388
rect 32508 45220 32564 45230
rect 32620 45220 32676 46956
rect 33068 46898 33124 46956
rect 33068 46846 33070 46898
rect 33122 46846 33124 46898
rect 33068 46834 33124 46846
rect 33292 46674 33348 46686
rect 33292 46622 33294 46674
rect 33346 46622 33348 46674
rect 32396 45218 32676 45220
rect 32396 45166 32510 45218
rect 32562 45166 32676 45218
rect 32396 45164 32676 45166
rect 32956 46002 33012 46014
rect 32956 45950 32958 46002
rect 33010 45950 33012 46002
rect 32284 45126 32340 45164
rect 32508 45154 32564 45164
rect 31948 44270 31950 44322
rect 32002 44270 32004 44322
rect 31948 44258 32004 44270
rect 32172 44882 32228 44894
rect 32172 44830 32174 44882
rect 32226 44830 32228 44882
rect 31164 43538 31444 43540
rect 31164 43486 31166 43538
rect 31218 43486 31444 43538
rect 31164 43484 31444 43486
rect 31612 44098 31668 44110
rect 31612 44046 31614 44098
rect 31666 44046 31668 44098
rect 31164 43204 31220 43484
rect 31164 43138 31220 43148
rect 31612 42980 31668 44046
rect 32172 43764 32228 44830
rect 32508 44660 32564 44670
rect 32508 44546 32564 44604
rect 32508 44494 32510 44546
rect 32562 44494 32564 44546
rect 32508 44482 32564 44494
rect 32956 44548 33012 45950
rect 33292 45780 33348 46622
rect 33404 46228 33460 48860
rect 33964 48132 34020 48972
rect 34076 49138 34132 49150
rect 34076 49086 34078 49138
rect 34130 49086 34132 49138
rect 34076 48356 34132 49086
rect 34300 49026 34356 49420
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 34300 48974 34302 49026
rect 34354 48974 34356 49026
rect 34300 48962 34356 48974
rect 34748 48916 34804 48926
rect 34748 48822 34804 48860
rect 34972 48916 35028 48926
rect 34972 48822 35028 48860
rect 34076 48290 34132 48300
rect 34636 48802 34692 48814
rect 34636 48750 34638 48802
rect 34690 48750 34692 48802
rect 34300 48132 34356 48142
rect 33740 48130 34468 48132
rect 33740 48078 34302 48130
rect 34354 48078 34468 48130
rect 33740 48076 34468 48078
rect 33516 47460 33572 47470
rect 33740 47460 33796 48076
rect 34300 48066 34356 48076
rect 33516 47458 33796 47460
rect 33516 47406 33518 47458
rect 33570 47406 33796 47458
rect 33516 47404 33796 47406
rect 33516 47394 33572 47404
rect 34300 47346 34356 47358
rect 34300 47294 34302 47346
rect 34354 47294 34356 47346
rect 33404 46162 33460 46172
rect 33628 47124 33684 47134
rect 33292 45714 33348 45724
rect 32956 44482 33012 44492
rect 33404 44994 33460 45006
rect 33404 44942 33406 44994
rect 33458 44942 33460 44994
rect 33404 44884 33460 44942
rect 32844 44436 32900 44446
rect 32844 44342 32900 44380
rect 32172 43698 32228 43708
rect 32396 44324 32452 44334
rect 31612 42924 31780 42980
rect 30940 42868 30996 42878
rect 30940 42866 31668 42868
rect 30940 42814 30942 42866
rect 30994 42814 31668 42866
rect 30940 42812 31668 42814
rect 30940 42802 30996 42812
rect 30828 42702 30830 42754
rect 30882 42702 30884 42754
rect 30828 42690 30884 42702
rect 31388 42530 31444 42542
rect 31388 42478 31390 42530
rect 31442 42478 31444 42530
rect 31388 42420 31444 42478
rect 31388 42354 31444 42364
rect 31276 42196 31332 42206
rect 31276 42102 31332 42140
rect 30828 42084 30884 42094
rect 30828 41748 30884 42028
rect 30940 41972 30996 41982
rect 30940 41878 30996 41916
rect 31612 41970 31668 42812
rect 31612 41918 31614 41970
rect 31666 41918 31668 41970
rect 31612 41906 31668 41918
rect 30828 41692 30996 41748
rect 30828 41412 30884 41422
rect 30716 41356 30828 41412
rect 30828 41346 30884 41356
rect 30940 41188 30996 41692
rect 30604 41022 30606 41074
rect 30658 41022 30660 41074
rect 30604 40404 30660 41022
rect 30604 40338 30660 40348
rect 30828 41132 30996 41188
rect 30828 40402 30884 41132
rect 30940 40516 30996 40526
rect 31724 40516 31780 42924
rect 32284 42196 32340 42206
rect 32284 42102 32340 42140
rect 32060 42084 32116 42094
rect 32060 41990 32116 42028
rect 31948 41972 32004 41982
rect 31836 41858 31892 41870
rect 31836 41806 31838 41858
rect 31890 41806 31892 41858
rect 31836 41412 31892 41806
rect 31948 41524 32004 41916
rect 32172 41858 32228 41870
rect 32172 41806 32174 41858
rect 32226 41806 32228 41858
rect 32172 41748 32228 41806
rect 32172 41682 32228 41692
rect 31948 41458 32004 41468
rect 31836 41346 31892 41356
rect 32060 41300 32116 41310
rect 32060 41186 32116 41244
rect 32060 41134 32062 41186
rect 32114 41134 32116 41186
rect 32060 41122 32116 41134
rect 32284 40628 32340 40638
rect 32284 40534 32340 40572
rect 30940 40514 31780 40516
rect 30940 40462 30942 40514
rect 30994 40462 31780 40514
rect 30940 40460 31780 40462
rect 30940 40450 30996 40460
rect 30828 40350 30830 40402
rect 30882 40350 30884 40402
rect 30828 40338 30884 40350
rect 31948 40402 32004 40414
rect 31948 40350 31950 40402
rect 32002 40350 32004 40402
rect 31948 39844 32004 40350
rect 31948 39778 32004 39788
rect 32284 39508 32340 39518
rect 32396 39508 32452 44268
rect 33404 44324 33460 44828
rect 33404 44258 33460 44268
rect 33516 44548 33572 44558
rect 33516 44322 33572 44492
rect 33516 44270 33518 44322
rect 33570 44270 33572 44322
rect 33516 44258 33572 44270
rect 32732 44098 32788 44110
rect 32732 44046 32734 44098
rect 32786 44046 32788 44098
rect 32732 43540 32788 44046
rect 33404 44100 33460 44110
rect 33404 43650 33460 44044
rect 33404 43598 33406 43650
rect 33458 43598 33460 43650
rect 33068 43540 33124 43550
rect 32732 43538 33124 43540
rect 32732 43486 33070 43538
rect 33122 43486 33124 43538
rect 32732 43484 33124 43486
rect 32620 42530 32676 42542
rect 32620 42478 32622 42530
rect 32674 42478 32676 42530
rect 32620 42084 32676 42478
rect 32620 42018 32676 42028
rect 33068 41972 33124 43484
rect 33068 41906 33124 41916
rect 33292 42082 33348 42094
rect 33292 42030 33294 42082
rect 33346 42030 33348 42082
rect 33292 41972 33348 42030
rect 33292 41906 33348 41916
rect 33180 41858 33236 41870
rect 33180 41806 33182 41858
rect 33234 41806 33236 41858
rect 33068 41748 33124 41758
rect 33068 41654 33124 41692
rect 33180 41412 33236 41806
rect 32732 41356 33236 41412
rect 32732 41298 32788 41356
rect 32732 41246 32734 41298
rect 32786 41246 32788 41298
rect 32732 41234 32788 41246
rect 32508 40516 32564 40526
rect 33404 40516 33460 43598
rect 32508 40514 33460 40516
rect 32508 40462 32510 40514
rect 32562 40462 33460 40514
rect 32508 40460 33460 40462
rect 33516 41972 33572 41982
rect 33516 41188 33572 41916
rect 32508 40450 32564 40460
rect 32508 40292 32564 40302
rect 32508 39618 32564 40236
rect 32508 39566 32510 39618
rect 32562 39566 32564 39618
rect 32508 39554 32564 39566
rect 33180 39620 33236 40460
rect 33404 39620 33460 39630
rect 33180 39618 33460 39620
rect 33180 39566 33406 39618
rect 33458 39566 33460 39618
rect 33180 39564 33460 39566
rect 33404 39554 33460 39564
rect 32284 39506 32452 39508
rect 32284 39454 32286 39506
rect 32338 39454 32452 39506
rect 32284 39452 32452 39454
rect 32844 39508 32900 39518
rect 33068 39508 33124 39518
rect 32844 39506 33124 39508
rect 32844 39454 32846 39506
rect 32898 39454 33070 39506
rect 33122 39454 33124 39506
rect 32844 39452 33124 39454
rect 31948 39396 32004 39406
rect 32284 39396 32340 39452
rect 32844 39442 32900 39452
rect 33068 39442 33124 39452
rect 31948 39394 32340 39396
rect 31948 39342 31950 39394
rect 32002 39342 32340 39394
rect 31948 39340 32340 39342
rect 32620 39394 32676 39406
rect 32620 39342 32622 39394
rect 32674 39342 32676 39394
rect 31276 38834 31332 38846
rect 31276 38782 31278 38834
rect 31330 38782 31332 38834
rect 30828 38724 30884 38762
rect 31276 38668 31332 38782
rect 29484 38612 29764 38668
rect 30492 38612 30660 38668
rect 30828 38658 30884 38668
rect 29484 38052 29540 38062
rect 29484 37958 29540 37996
rect 29484 36596 29540 36606
rect 29484 36482 29540 36540
rect 29484 36430 29486 36482
rect 29538 36430 29540 36482
rect 29484 36418 29540 36430
rect 29260 35924 29316 35934
rect 29148 35868 29260 35924
rect 28588 35810 28644 35822
rect 28588 35758 28590 35810
rect 28642 35758 28644 35810
rect 28252 35700 28308 35710
rect 28588 35700 28644 35758
rect 28252 35698 28756 35700
rect 28252 35646 28254 35698
rect 28306 35646 28756 35698
rect 28252 35644 28756 35646
rect 28252 35634 28308 35644
rect 27916 35588 27972 35598
rect 27916 35494 27972 35532
rect 28700 35028 28756 35644
rect 28812 35698 28868 35868
rect 29260 35830 29316 35868
rect 29372 35924 29428 35934
rect 29372 35922 29652 35924
rect 29372 35870 29374 35922
rect 29426 35870 29652 35922
rect 29372 35868 29652 35870
rect 29372 35858 29428 35868
rect 28812 35646 28814 35698
rect 28866 35646 28868 35698
rect 28812 35634 28868 35646
rect 29484 35698 29540 35710
rect 29484 35646 29486 35698
rect 29538 35646 29540 35698
rect 29484 35476 29540 35646
rect 29260 35420 29540 35476
rect 29260 35028 29316 35420
rect 29484 35140 29540 35150
rect 29596 35140 29652 35868
rect 29708 35922 29764 38612
rect 30268 38052 30324 38062
rect 30268 37958 30324 37996
rect 29820 37940 29876 37950
rect 29820 37846 29876 37884
rect 30492 37268 30548 37278
rect 30492 37174 30548 37212
rect 30044 37156 30100 37166
rect 30044 37062 30100 37100
rect 30044 36596 30100 36606
rect 30044 36502 30100 36540
rect 29708 35870 29710 35922
rect 29762 35870 29764 35922
rect 29708 35858 29764 35870
rect 30268 35924 30324 35934
rect 30604 35924 30660 38612
rect 31052 38612 31332 38668
rect 31948 38724 32004 39340
rect 32620 38668 32676 39342
rect 31948 38658 32004 38668
rect 32508 38612 32676 38668
rect 33292 39394 33348 39406
rect 33292 39342 33294 39394
rect 33346 39342 33348 39394
rect 30716 37940 30772 37950
rect 30716 37846 30772 37884
rect 31052 37938 31108 38612
rect 32508 38162 32564 38612
rect 33292 38276 33348 39342
rect 33292 38210 33348 38220
rect 33404 39284 33460 39294
rect 32508 38110 32510 38162
rect 32562 38110 32564 38162
rect 32508 38098 32564 38110
rect 31724 38050 31780 38062
rect 31724 37998 31726 38050
rect 31778 37998 31780 38050
rect 31052 37886 31054 37938
rect 31106 37886 31108 37938
rect 30940 37156 30996 37166
rect 30940 37062 30996 37100
rect 30828 36258 30884 36270
rect 30828 36206 30830 36258
rect 30882 36206 30884 36258
rect 30828 36036 30884 36206
rect 30828 35970 30884 35980
rect 30716 35924 30772 35934
rect 30604 35922 30772 35924
rect 30604 35870 30718 35922
rect 30770 35870 30772 35922
rect 30604 35868 30772 35870
rect 30268 35830 30324 35868
rect 30716 35858 30772 35868
rect 30492 35812 30548 35822
rect 30492 35718 30548 35756
rect 29484 35138 29652 35140
rect 29484 35086 29486 35138
rect 29538 35086 29652 35138
rect 29484 35084 29652 35086
rect 30380 35586 30436 35598
rect 30380 35534 30382 35586
rect 30434 35534 30436 35586
rect 30380 35140 30436 35534
rect 30604 35140 30660 35150
rect 30380 35138 30660 35140
rect 30380 35086 30606 35138
rect 30658 35086 30660 35138
rect 30380 35084 30660 35086
rect 29484 35074 29540 35084
rect 30604 35074 30660 35084
rect 28700 34972 29204 35028
rect 29148 34916 29204 34972
rect 29148 34822 29204 34860
rect 27468 34290 27524 34300
rect 27132 34190 27134 34242
rect 27186 34190 27188 34242
rect 27132 34178 27188 34190
rect 29260 34018 29316 34972
rect 29484 34916 29540 34926
rect 29372 34692 29428 34702
rect 29372 34598 29428 34636
rect 29260 33966 29262 34018
rect 29314 33966 29316 34018
rect 29260 33954 29316 33966
rect 27132 33908 27188 33918
rect 26684 33124 26740 33134
rect 26684 33122 26852 33124
rect 26684 33070 26686 33122
rect 26738 33070 26852 33122
rect 26684 33068 26852 33070
rect 26684 33058 26740 33068
rect 26684 31892 26740 31902
rect 26684 31778 26740 31836
rect 26684 31726 26686 31778
rect 26738 31726 26740 31778
rect 26684 31714 26740 31726
rect 26796 31780 26852 33068
rect 26796 31724 27076 31780
rect 26572 31500 26852 31556
rect 26684 30884 26740 30894
rect 26572 30212 26628 30222
rect 26572 30118 26628 30156
rect 26572 29988 26628 29998
rect 26684 29988 26740 30828
rect 26572 29986 26740 29988
rect 26572 29934 26574 29986
rect 26626 29934 26740 29986
rect 26572 29932 26740 29934
rect 26572 29922 26628 29932
rect 26796 29876 26852 31500
rect 26908 30324 26964 30334
rect 26908 30098 26964 30268
rect 26908 30046 26910 30098
rect 26962 30046 26964 30098
rect 26908 30034 26964 30046
rect 26796 29820 26964 29876
rect 26460 28802 26516 28812
rect 26684 29764 26740 29774
rect 25564 27694 25566 27746
rect 25618 27694 25620 27746
rect 25564 26908 25620 27694
rect 26236 28530 26292 28542
rect 26236 28478 26238 28530
rect 26290 28478 26292 28530
rect 26236 27860 26292 28478
rect 26236 27188 26292 27804
rect 26348 27188 26404 27198
rect 26236 27186 26404 27188
rect 26236 27134 26350 27186
rect 26402 27134 26404 27186
rect 26236 27132 26404 27134
rect 26348 27122 26404 27132
rect 26684 26908 26740 29708
rect 26908 29652 26964 29820
rect 27020 29764 27076 31724
rect 27132 30660 27188 33852
rect 29484 33346 29540 34860
rect 30268 34916 30324 34926
rect 30268 34822 30324 34860
rect 30492 34690 30548 34702
rect 30492 34638 30494 34690
rect 30546 34638 30548 34690
rect 30380 34244 30436 34254
rect 30492 34244 30548 34638
rect 30380 34242 30548 34244
rect 30380 34190 30382 34242
rect 30434 34190 30548 34242
rect 30380 34188 30548 34190
rect 30380 34178 30436 34188
rect 29596 34132 29652 34142
rect 29652 34076 29988 34132
rect 29596 34038 29652 34076
rect 29932 33460 29988 34076
rect 30380 33460 30436 33470
rect 29932 33458 30380 33460
rect 29932 33406 29934 33458
rect 29986 33406 30380 33458
rect 29932 33404 30380 33406
rect 29932 33394 29988 33404
rect 29484 33294 29486 33346
rect 29538 33294 29540 33346
rect 29484 33282 29540 33294
rect 29148 33234 29204 33246
rect 29148 33182 29150 33234
rect 29202 33182 29204 33234
rect 27244 32452 27300 32462
rect 27244 32358 27300 32396
rect 29148 32452 29204 33182
rect 30044 33236 30100 33246
rect 29260 33122 29316 33134
rect 29260 33070 29262 33122
rect 29314 33070 29316 33122
rect 29260 32676 29316 33070
rect 29708 32788 29764 32798
rect 29372 32676 29428 32686
rect 29260 32674 29428 32676
rect 29260 32622 29374 32674
rect 29426 32622 29428 32674
rect 29260 32620 29428 32622
rect 29372 32610 29428 32620
rect 27356 31892 27412 31902
rect 27356 31798 27412 31836
rect 28252 31780 28308 31790
rect 28140 31724 28252 31780
rect 28028 31220 28084 31230
rect 28028 30994 28084 31164
rect 28028 30942 28030 30994
rect 28082 30942 28084 30994
rect 27356 30884 27412 30894
rect 27356 30790 27412 30828
rect 27132 30604 27300 30660
rect 27132 30436 27188 30446
rect 27132 30210 27188 30380
rect 27132 30158 27134 30210
rect 27186 30158 27188 30210
rect 27132 30146 27188 30158
rect 27020 29698 27076 29708
rect 26796 29596 26964 29652
rect 26796 28644 26852 29596
rect 26796 28588 26964 28644
rect 25564 26852 26404 26908
rect 25676 26292 25732 26302
rect 25452 26238 25454 26290
rect 25506 26238 25508 26290
rect 25340 26180 25396 26190
rect 25340 26086 25396 26124
rect 25340 25396 25396 25406
rect 25116 25284 25172 25294
rect 25116 21476 25172 25228
rect 25340 25282 25396 25340
rect 25340 25230 25342 25282
rect 25394 25230 25396 25282
rect 25228 24610 25284 24622
rect 25228 24558 25230 24610
rect 25282 24558 25284 24610
rect 25228 24500 25284 24558
rect 25340 24612 25396 25230
rect 25452 24836 25508 26238
rect 25452 24770 25508 24780
rect 25564 26290 25732 26292
rect 25564 26238 25678 26290
rect 25730 26238 25732 26290
rect 25564 26236 25732 26238
rect 25564 25508 25620 26236
rect 25676 26226 25732 26236
rect 26124 26068 26180 26078
rect 26124 25974 26180 26012
rect 26348 26068 26404 26852
rect 26572 26852 26740 26908
rect 26460 26068 26516 26078
rect 26348 26066 26516 26068
rect 26348 26014 26462 26066
rect 26514 26014 26516 26066
rect 26348 26012 26516 26014
rect 25564 24722 25620 25452
rect 25676 25618 25732 25630
rect 25676 25566 25678 25618
rect 25730 25566 25732 25618
rect 25676 25284 25732 25566
rect 25676 25218 25732 25228
rect 25564 24670 25566 24722
rect 25618 24670 25620 24722
rect 25340 24556 25508 24612
rect 25228 24444 25396 24500
rect 25340 24052 25396 24444
rect 25340 23986 25396 23996
rect 25228 23940 25284 23950
rect 25228 21698 25284 23884
rect 25340 23380 25396 23390
rect 25340 23042 25396 23324
rect 25340 22990 25342 23042
rect 25394 22990 25396 23042
rect 25340 21812 25396 22990
rect 25452 22148 25508 24556
rect 25564 23938 25620 24670
rect 26124 25172 26180 25182
rect 25564 23886 25566 23938
rect 25618 23886 25620 23938
rect 25564 22370 25620 23886
rect 25788 24610 25844 24622
rect 25788 24558 25790 24610
rect 25842 24558 25844 24610
rect 25788 24500 25844 24558
rect 25676 23044 25732 23054
rect 25676 22950 25732 22988
rect 25788 22594 25844 24444
rect 25788 22542 25790 22594
rect 25842 22542 25844 22594
rect 25788 22530 25844 22542
rect 25564 22318 25566 22370
rect 25618 22318 25620 22370
rect 25564 22306 25620 22318
rect 25452 22092 25732 22148
rect 25340 21756 25620 21812
rect 25228 21646 25230 21698
rect 25282 21646 25284 21698
rect 25228 21634 25284 21646
rect 25452 21588 25508 21598
rect 25452 21494 25508 21532
rect 25116 21410 25172 21420
rect 25004 20862 25006 20914
rect 25058 20862 25060 20914
rect 25004 20850 25060 20862
rect 25452 21364 25508 21374
rect 24556 20804 24612 20814
rect 24556 20710 24612 20748
rect 25452 20692 25508 21308
rect 25228 20690 25508 20692
rect 25228 20638 25454 20690
rect 25506 20638 25508 20690
rect 25228 20636 25508 20638
rect 24668 19908 24724 19918
rect 24668 19012 24724 19852
rect 25004 19236 25060 19246
rect 25004 19142 25060 19180
rect 25228 19124 25284 20636
rect 25452 20626 25508 20636
rect 25564 20018 25620 21756
rect 25676 21140 25732 22092
rect 26124 22146 26180 25116
rect 26348 24948 26404 26012
rect 26460 26002 26516 26012
rect 26348 24854 26404 24892
rect 26124 22094 26126 22146
rect 26178 22094 26180 22146
rect 25788 21364 25844 21374
rect 25788 21270 25844 21308
rect 25676 21084 25956 21140
rect 25676 20804 25732 20814
rect 25676 20802 25844 20804
rect 25676 20750 25678 20802
rect 25730 20750 25844 20802
rect 25676 20748 25844 20750
rect 25676 20738 25732 20748
rect 25564 19966 25566 20018
rect 25618 19966 25620 20018
rect 25564 19908 25620 19966
rect 25564 19842 25620 19852
rect 25676 20244 25732 20254
rect 25676 19572 25732 20188
rect 24668 19010 24836 19012
rect 24668 18958 24670 19010
rect 24722 18958 24836 19010
rect 24668 18956 24836 18958
rect 24668 18946 24724 18956
rect 24332 18398 24334 18450
rect 24386 18398 24388 18450
rect 24332 18386 24388 18398
rect 24108 18340 24164 18350
rect 23772 18338 24164 18340
rect 23772 18286 23774 18338
rect 23826 18286 24110 18338
rect 24162 18286 24164 18338
rect 23772 18284 24164 18286
rect 23436 16436 23492 16446
rect 23436 16098 23492 16380
rect 23436 16046 23438 16098
rect 23490 16046 23492 16098
rect 23436 16034 23492 16046
rect 23100 15874 23156 15886
rect 23100 15822 23102 15874
rect 23154 15822 23156 15874
rect 23100 15204 23156 15822
rect 23100 15138 23156 15148
rect 23324 15652 23380 15662
rect 23324 15538 23380 15596
rect 23324 15486 23326 15538
rect 23378 15486 23380 15538
rect 22876 14578 22932 14588
rect 22316 13636 22372 13646
rect 22316 13542 22372 13580
rect 22316 13188 22372 13198
rect 22988 13188 23044 13198
rect 22316 12962 22372 13132
rect 22316 12910 22318 12962
rect 22370 12910 22372 12962
rect 22316 12898 22372 12910
rect 22428 13186 23044 13188
rect 22428 13134 22990 13186
rect 23042 13134 23044 13186
rect 22428 13132 23044 13134
rect 22428 12738 22484 13132
rect 22988 13122 23044 13132
rect 22764 12964 22820 12974
rect 22764 12870 22820 12908
rect 23324 12962 23380 15486
rect 23436 13860 23492 13870
rect 23436 13074 23492 13804
rect 23548 13300 23604 17276
rect 23772 17220 23828 18284
rect 24108 18274 24164 18284
rect 24668 18340 24724 18350
rect 24668 18246 24724 18284
rect 23884 17892 23940 17902
rect 23884 17666 23940 17836
rect 23884 17614 23886 17666
rect 23938 17614 23940 17666
rect 23884 17602 23940 17614
rect 24668 17666 24724 17678
rect 24668 17614 24670 17666
rect 24722 17614 24724 17666
rect 24220 17444 24276 17454
rect 24668 17444 24724 17614
rect 24220 17442 24724 17444
rect 24220 17390 24222 17442
rect 24274 17390 24724 17442
rect 24220 17388 24724 17390
rect 24220 17378 24276 17388
rect 24668 17332 24724 17388
rect 24668 17266 24724 17276
rect 23772 17154 23828 17164
rect 24332 17220 24388 17230
rect 23884 16996 23940 17006
rect 23884 16902 23940 16940
rect 23660 16772 23716 16782
rect 23660 15540 23716 16716
rect 24220 16660 24276 16670
rect 24220 16210 24276 16604
rect 24220 16158 24222 16210
rect 24274 16158 24276 16210
rect 24220 16146 24276 16158
rect 23660 15446 23716 15484
rect 23772 16100 23828 16110
rect 23772 15874 23828 16044
rect 24332 16098 24388 17164
rect 24668 16996 24724 17006
rect 24780 16996 24836 18956
rect 25228 18452 25284 19068
rect 25228 18386 25284 18396
rect 25340 19516 25732 19572
rect 24892 18228 24948 18238
rect 24892 17890 24948 18172
rect 24892 17838 24894 17890
rect 24946 17838 24948 17890
rect 24892 17826 24948 17838
rect 25340 17666 25396 19516
rect 25452 19348 25508 19358
rect 25452 19254 25508 19292
rect 25676 19124 25732 19134
rect 25676 19030 25732 19068
rect 25676 18900 25732 18910
rect 25564 18844 25676 18900
rect 25564 18674 25620 18844
rect 25676 18834 25732 18844
rect 25564 18622 25566 18674
rect 25618 18622 25620 18674
rect 25564 18610 25620 18622
rect 25452 18450 25508 18462
rect 25452 18398 25454 18450
rect 25506 18398 25508 18450
rect 25452 18228 25508 18398
rect 25452 18162 25508 18172
rect 25564 17892 25620 17902
rect 25340 17614 25342 17666
rect 25394 17614 25396 17666
rect 25340 17602 25396 17614
rect 25452 17836 25564 17892
rect 25116 17554 25172 17566
rect 25116 17502 25118 17554
rect 25170 17502 25172 17554
rect 24724 16940 24836 16996
rect 25004 17442 25060 17454
rect 25004 17390 25006 17442
rect 25058 17390 25060 17442
rect 24668 16930 24724 16940
rect 24332 16046 24334 16098
rect 24386 16046 24388 16098
rect 24332 16034 24388 16046
rect 24556 16884 24612 16894
rect 24220 15988 24276 15998
rect 23772 15822 23774 15874
rect 23826 15822 23828 15874
rect 23548 13234 23604 13244
rect 23436 13022 23438 13074
rect 23490 13022 23492 13074
rect 23436 13010 23492 13022
rect 23324 12910 23326 12962
rect 23378 12910 23380 12962
rect 23324 12898 23380 12910
rect 22428 12686 22430 12738
rect 22482 12686 22484 12738
rect 22428 12674 22484 12686
rect 22988 12852 23044 12862
rect 22988 12402 23044 12796
rect 23548 12850 23604 12862
rect 23548 12798 23550 12850
rect 23602 12798 23604 12850
rect 22988 12350 22990 12402
rect 23042 12350 23044 12402
rect 22988 12338 23044 12350
rect 23436 12404 23492 12414
rect 23436 12310 23492 12348
rect 22148 11676 22260 11732
rect 22876 12066 22932 12078
rect 22876 12014 22878 12066
rect 22930 12014 22932 12066
rect 22092 11666 22148 11676
rect 22876 11284 22932 12014
rect 23436 11508 23492 11518
rect 23436 11414 23492 11452
rect 22876 10498 22932 11228
rect 22876 10446 22878 10498
rect 22930 10446 22932 10498
rect 22876 10434 22932 10446
rect 23324 10498 23380 10510
rect 23324 10446 23326 10498
rect 23378 10446 23380 10498
rect 23324 10052 23380 10446
rect 23324 9986 23380 9996
rect 22316 9828 22372 9838
rect 22092 9772 22316 9828
rect 21980 9602 22036 9614
rect 21980 9550 21982 9602
rect 22034 9550 22036 9602
rect 21980 8820 22036 9550
rect 21980 8754 22036 8764
rect 21868 8206 21870 8258
rect 21922 8206 21924 8258
rect 20748 8036 20804 8046
rect 20748 8034 21028 8036
rect 20748 7982 20750 8034
rect 20802 7982 21028 8034
rect 20748 7980 21028 7982
rect 20748 7970 20804 7980
rect 20972 7586 21028 7980
rect 20972 7534 20974 7586
rect 21026 7534 21028 7586
rect 20972 7522 21028 7534
rect 21868 7700 21924 8206
rect 20300 7422 20302 7474
rect 20354 7422 20356 7474
rect 18508 6750 18510 6802
rect 18562 6750 18564 6802
rect 18508 6738 18564 6750
rect 18956 6692 19012 6702
rect 18956 6598 19012 6636
rect 19628 6692 19684 6702
rect 18284 5966 18286 6018
rect 18338 5966 18340 6018
rect 18284 5954 18340 5966
rect 18508 6020 18564 6030
rect 18508 5926 18564 5964
rect 19404 6020 19460 6030
rect 17948 5906 18116 5908
rect 17948 5854 17950 5906
rect 18002 5854 18116 5906
rect 17948 5852 18116 5854
rect 17948 5842 18004 5852
rect 17276 5182 17278 5234
rect 17330 5182 17332 5234
rect 17276 5170 17332 5182
rect 19404 5234 19460 5964
rect 19404 5182 19406 5234
rect 19458 5182 19460 5234
rect 19404 5170 19460 5182
rect 19628 5236 19684 6636
rect 20300 6692 20356 7422
rect 21868 6804 21924 7644
rect 21868 6738 21924 6748
rect 20300 6626 20356 6636
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 21868 5908 21924 5918
rect 22092 5908 22148 9772
rect 22316 9734 22372 9772
rect 22540 9716 22596 9726
rect 22428 9714 22596 9716
rect 22428 9662 22542 9714
rect 22594 9662 22596 9714
rect 22428 9660 22596 9662
rect 22316 8932 22372 8942
rect 22316 8258 22372 8876
rect 22428 8372 22484 9660
rect 22540 9650 22596 9660
rect 23100 9714 23156 9726
rect 23100 9662 23102 9714
rect 23154 9662 23156 9714
rect 22428 8370 23044 8372
rect 22428 8318 22430 8370
rect 22482 8318 23044 8370
rect 22428 8316 23044 8318
rect 22428 8306 22484 8316
rect 22316 8206 22318 8258
rect 22370 8206 22372 8258
rect 22316 7812 22372 8206
rect 22988 8258 23044 8316
rect 22988 8206 22990 8258
rect 23042 8206 23044 8258
rect 22988 8194 23044 8206
rect 22876 8148 22932 8158
rect 22876 8054 22932 8092
rect 22316 7746 22372 7756
rect 23100 7362 23156 9662
rect 23100 7310 23102 7362
rect 23154 7310 23156 7362
rect 23100 6916 23156 7310
rect 23548 7252 23604 12798
rect 23772 12628 23828 15822
rect 24108 15874 24164 15886
rect 24108 15822 24110 15874
rect 24162 15822 24164 15874
rect 24108 13860 24164 15822
rect 24220 15538 24276 15932
rect 24556 15988 24612 16828
rect 25004 16436 25060 17390
rect 25004 16370 25060 16380
rect 25116 17444 25172 17502
rect 25004 16100 25060 16110
rect 25116 16100 25172 17388
rect 25228 17220 25284 17230
rect 25228 17106 25284 17164
rect 25228 17054 25230 17106
rect 25282 17054 25284 17106
rect 25228 17042 25284 17054
rect 25228 16884 25284 16894
rect 25228 16790 25284 16828
rect 25452 16324 25508 17836
rect 25564 17826 25620 17836
rect 25788 17890 25844 20748
rect 25900 18116 25956 21084
rect 26124 20132 26180 22094
rect 26460 23044 26516 23054
rect 26460 22372 26516 22988
rect 26460 21698 26516 22316
rect 26460 21646 26462 21698
rect 26514 21646 26516 21698
rect 26460 21634 26516 21646
rect 26572 21812 26628 26852
rect 26684 26178 26740 26190
rect 26684 26126 26686 26178
rect 26738 26126 26740 26178
rect 26684 25620 26740 26126
rect 26684 25554 26740 25564
rect 26684 24836 26740 24846
rect 26684 24742 26740 24780
rect 26796 24052 26852 24062
rect 26684 22258 26740 22270
rect 26684 22206 26686 22258
rect 26738 22206 26740 22258
rect 26684 21924 26740 22206
rect 26684 21858 26740 21868
rect 26796 22258 26852 23996
rect 26796 22206 26798 22258
rect 26850 22206 26852 22258
rect 26348 21476 26404 21486
rect 26236 21474 26404 21476
rect 26236 21422 26350 21474
rect 26402 21422 26404 21474
rect 26236 21420 26404 21422
rect 26236 20244 26292 21420
rect 26348 21410 26404 21420
rect 26572 21476 26628 21756
rect 26572 21410 26628 21420
rect 26796 21252 26852 22206
rect 26908 22148 26964 28588
rect 27132 28532 27188 28542
rect 27244 28532 27300 30604
rect 27692 29652 27748 29662
rect 28028 29652 28084 30942
rect 27692 29650 28084 29652
rect 27692 29598 27694 29650
rect 27746 29598 28084 29650
rect 27692 29596 28084 29598
rect 27692 29586 27748 29596
rect 28028 29426 28084 29596
rect 28028 29374 28030 29426
rect 28082 29374 28084 29426
rect 28028 29362 28084 29374
rect 28140 30212 28196 31724
rect 28252 31714 28308 31724
rect 29148 31108 29204 32396
rect 27580 29204 27636 29214
rect 28140 29204 28196 30156
rect 28364 31106 29204 31108
rect 28364 31054 29150 31106
rect 29202 31054 29204 31106
rect 28364 31052 29204 31054
rect 28364 30210 28420 31052
rect 29148 31042 29204 31052
rect 29596 32004 29652 32014
rect 29260 30996 29316 31006
rect 29260 30770 29316 30940
rect 29260 30718 29262 30770
rect 29314 30718 29316 30770
rect 29260 30436 29316 30718
rect 28364 30158 28366 30210
rect 28418 30158 28420 30210
rect 28364 30146 28420 30158
rect 28588 30380 29316 30436
rect 29484 30772 29540 30782
rect 28476 30100 28532 30110
rect 28476 30006 28532 30044
rect 27580 28866 27636 29148
rect 27916 29148 28196 29204
rect 28252 29652 28308 29662
rect 27580 28814 27582 28866
rect 27634 28814 27636 28866
rect 27580 28802 27636 28814
rect 27804 28868 27860 28878
rect 27356 28644 27412 28654
rect 27356 28550 27412 28588
rect 27132 28530 27300 28532
rect 27132 28478 27134 28530
rect 27186 28478 27300 28530
rect 27132 28476 27300 28478
rect 27132 28466 27188 28476
rect 27580 28418 27636 28430
rect 27580 28366 27582 28418
rect 27634 28366 27636 28418
rect 27580 27972 27636 28366
rect 27692 27972 27748 27982
rect 27580 27970 27748 27972
rect 27580 27918 27694 27970
rect 27746 27918 27748 27970
rect 27580 27916 27748 27918
rect 27692 27906 27748 27916
rect 27804 25618 27860 28812
rect 27916 28642 27972 29148
rect 28252 28868 28308 29596
rect 28588 28980 28644 30380
rect 28700 30212 28756 30222
rect 29036 30212 29092 30222
rect 28700 30210 29092 30212
rect 28700 30158 28702 30210
rect 28754 30158 29038 30210
rect 29090 30158 29092 30210
rect 28700 30156 29092 30158
rect 28700 30146 28756 30156
rect 29036 30146 29092 30156
rect 29484 30210 29540 30716
rect 29484 30158 29486 30210
rect 29538 30158 29540 30210
rect 29484 30146 29540 30158
rect 29596 30212 29652 31948
rect 29708 31220 29764 32732
rect 30044 32004 30100 33180
rect 30156 32562 30212 33404
rect 30380 33366 30436 33404
rect 30156 32510 30158 32562
rect 30210 32510 30212 32562
rect 30156 32498 30212 32510
rect 30828 32564 30884 32574
rect 31052 32564 31108 37886
rect 31164 37940 31220 37950
rect 31164 37266 31220 37884
rect 31500 37492 31556 37502
rect 31500 37398 31556 37436
rect 31164 37214 31166 37266
rect 31218 37214 31220 37266
rect 31164 36484 31220 37214
rect 31724 37268 31780 37998
rect 31724 37202 31780 37212
rect 32396 37266 32452 37278
rect 32396 37214 32398 37266
rect 32450 37214 32452 37266
rect 32060 37156 32116 37166
rect 32060 37062 32116 37100
rect 31500 36484 31556 36494
rect 31164 36482 31556 36484
rect 31164 36430 31166 36482
rect 31218 36430 31502 36482
rect 31554 36430 31556 36482
rect 31164 36428 31556 36430
rect 31164 36418 31220 36428
rect 31500 36418 31556 36428
rect 31836 36260 31892 36270
rect 31892 36204 32004 36260
rect 31836 36166 31892 36204
rect 30828 32562 31108 32564
rect 30828 32510 30830 32562
rect 30882 32510 31108 32562
rect 30828 32508 31108 32510
rect 31276 35140 31332 35150
rect 31276 32562 31332 35084
rect 31948 33236 32004 36204
rect 32172 36258 32228 36270
rect 32172 36206 32174 36258
rect 32226 36206 32228 36258
rect 32172 36036 32228 36206
rect 32396 36260 32452 37214
rect 33068 37268 33124 37278
rect 33068 37174 33124 37212
rect 33404 36932 33460 39228
rect 33404 36866 33460 36876
rect 32508 36484 32564 36494
rect 32508 36370 32564 36428
rect 33516 36484 33572 41132
rect 33516 36418 33572 36428
rect 32508 36318 32510 36370
rect 32562 36318 32564 36370
rect 32508 36306 32564 36318
rect 32396 36194 32452 36204
rect 32172 35970 32228 35980
rect 33404 34914 33460 34926
rect 33404 34862 33406 34914
rect 33458 34862 33460 34914
rect 33180 34804 33236 34814
rect 33404 34804 33460 34862
rect 33236 34748 33460 34804
rect 33180 34710 33236 34748
rect 33180 34130 33236 34142
rect 33180 34078 33182 34130
rect 33234 34078 33236 34130
rect 32508 34018 32564 34030
rect 32508 33966 32510 34018
rect 32562 33966 32564 34018
rect 32508 33908 32564 33966
rect 32508 33842 32564 33852
rect 32732 33460 32788 33470
rect 32732 33366 32788 33404
rect 33180 33460 33236 34078
rect 33516 34132 33572 34142
rect 33516 33684 33572 34076
rect 33628 34020 33684 47068
rect 33964 46676 34020 46686
rect 33852 46620 33964 46676
rect 33740 45106 33796 45118
rect 33740 45054 33742 45106
rect 33794 45054 33796 45106
rect 33740 44884 33796 45054
rect 33740 44818 33796 44828
rect 33740 44436 33796 44446
rect 33740 44322 33796 44380
rect 33740 44270 33742 44322
rect 33794 44270 33796 44322
rect 33740 44258 33796 44270
rect 33852 43876 33908 46620
rect 33964 46582 34020 46620
rect 34300 46562 34356 47294
rect 34412 47012 34468 48076
rect 34412 46946 34468 46956
rect 34412 46786 34468 46798
rect 34412 46734 34414 46786
rect 34466 46734 34468 46786
rect 34412 46676 34468 46734
rect 34636 46786 34692 48750
rect 35420 48804 35476 48814
rect 35644 48804 35700 49756
rect 35756 49586 35812 51772
rect 35868 51380 35924 51884
rect 35980 51874 36036 51884
rect 35980 51604 36036 51614
rect 35980 51510 36036 51548
rect 35980 51380 36036 51390
rect 36204 51380 36260 51390
rect 35868 51324 35980 51380
rect 35868 51156 35924 51166
rect 35868 51062 35924 51100
rect 35980 50594 36036 51324
rect 35980 50542 35982 50594
rect 36034 50542 36036 50594
rect 35980 50530 36036 50542
rect 36092 51378 36260 51380
rect 36092 51326 36206 51378
rect 36258 51326 36260 51378
rect 36092 51324 36260 51326
rect 36092 50428 36148 51324
rect 36204 51314 36260 51324
rect 36204 50820 36260 50830
rect 36316 50820 36372 51996
rect 36428 51940 36484 52670
rect 37660 52722 37716 52734
rect 37660 52670 37662 52722
rect 37714 52670 37716 52722
rect 37660 52276 37716 52670
rect 37660 52210 37716 52220
rect 36428 51884 36820 51940
rect 36204 50818 36372 50820
rect 36204 50766 36206 50818
rect 36258 50766 36372 50818
rect 36204 50764 36372 50766
rect 36428 51378 36484 51390
rect 36652 51380 36708 51390
rect 36428 51326 36430 51378
rect 36482 51326 36484 51378
rect 36204 50754 36260 50764
rect 36092 50372 36260 50428
rect 36204 49812 36260 50372
rect 36428 50372 36484 51326
rect 36428 50306 36484 50316
rect 36540 51378 36708 51380
rect 36540 51326 36654 51378
rect 36706 51326 36708 51378
rect 36540 51324 36708 51326
rect 36204 49718 36260 49756
rect 36540 49588 36596 51324
rect 36652 51314 36708 51324
rect 36764 51268 36820 51884
rect 37100 51492 37156 51502
rect 36988 51378 37044 51390
rect 36988 51326 36990 51378
rect 37042 51326 37044 51378
rect 36876 51268 36932 51278
rect 36764 51266 36932 51268
rect 36764 51214 36878 51266
rect 36930 51214 36932 51266
rect 36764 51212 36932 51214
rect 36876 51202 36932 51212
rect 36988 51044 37044 51326
rect 36988 50978 37044 50988
rect 36988 50596 37044 50606
rect 36988 50502 37044 50540
rect 37100 50482 37156 51436
rect 37212 51492 37268 51502
rect 37212 51490 37380 51492
rect 37212 51438 37214 51490
rect 37266 51438 37380 51490
rect 37212 51436 37380 51438
rect 37212 51426 37268 51436
rect 37100 50430 37102 50482
rect 37154 50430 37156 50482
rect 37100 50418 37156 50430
rect 37212 50820 37268 50830
rect 35756 49534 35758 49586
rect 35810 49534 35812 49586
rect 35756 49522 35812 49534
rect 36092 49532 36596 49588
rect 36652 50372 36708 50382
rect 36652 49922 36708 50316
rect 36876 50260 36932 50270
rect 36652 49870 36654 49922
rect 36706 49870 36708 49922
rect 36652 49588 36708 49870
rect 36092 49250 36148 49532
rect 36652 49522 36708 49532
rect 36764 50148 36820 50158
rect 36092 49198 36094 49250
rect 36146 49198 36148 49250
rect 36092 49186 36148 49198
rect 36204 49028 36260 49038
rect 36204 48934 36260 48972
rect 36428 48916 36484 48926
rect 36764 48916 36820 50092
rect 36876 49810 36932 50204
rect 37212 50036 37268 50764
rect 37324 50260 37380 51436
rect 37772 51380 37828 52892
rect 37884 52882 37940 52892
rect 37884 52722 37940 52734
rect 37884 52670 37886 52722
rect 37938 52670 37940 52722
rect 37884 51604 37940 52670
rect 37996 52388 38052 53564
rect 38108 53508 38164 53518
rect 38108 53414 38164 53452
rect 38108 53060 38164 53070
rect 38108 52946 38164 53004
rect 38108 52894 38110 52946
rect 38162 52894 38164 52946
rect 38108 52882 38164 52894
rect 37996 52294 38052 52332
rect 38220 52836 38276 52846
rect 38108 52050 38164 52062
rect 38108 51998 38110 52050
rect 38162 51998 38164 52050
rect 37884 51538 37940 51548
rect 37996 51940 38052 51950
rect 37324 50194 37380 50204
rect 37660 50594 37716 50606
rect 37660 50542 37662 50594
rect 37714 50542 37716 50594
rect 37548 50036 37604 50046
rect 37212 50034 37604 50036
rect 37212 49982 37550 50034
rect 37602 49982 37604 50034
rect 37212 49980 37604 49982
rect 37548 49970 37604 49980
rect 36876 49758 36878 49810
rect 36930 49758 36932 49810
rect 36876 49746 36932 49758
rect 37100 49924 37156 49934
rect 36484 48860 36820 48916
rect 36876 49252 36932 49262
rect 36092 48804 36148 48814
rect 35644 48748 36092 48804
rect 35420 48710 35476 48748
rect 36092 48710 36148 48748
rect 36204 48244 36260 48254
rect 36204 48150 36260 48188
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 36428 47570 36484 48860
rect 36428 47518 36430 47570
rect 36482 47518 36484 47570
rect 36428 47506 36484 47518
rect 34636 46734 34638 46786
rect 34690 46734 34692 46786
rect 34636 46722 34692 46734
rect 34748 47012 34804 47022
rect 34412 46610 34468 46620
rect 34300 46510 34302 46562
rect 34354 46510 34356 46562
rect 34300 46498 34356 46510
rect 33964 45108 34020 45118
rect 33964 45014 34020 45052
rect 34412 45108 34468 45118
rect 34748 45108 34804 46956
rect 35756 47012 35812 47022
rect 35756 46898 35812 46956
rect 35756 46846 35758 46898
rect 35810 46846 35812 46898
rect 35756 46834 35812 46846
rect 36316 47012 36372 47022
rect 36316 46674 36372 46956
rect 36316 46622 36318 46674
rect 36370 46622 36372 46674
rect 36316 46610 36372 46622
rect 35420 46562 35476 46574
rect 35420 46510 35422 46562
rect 35474 46510 35476 46562
rect 35420 46450 35476 46510
rect 35420 46398 35422 46450
rect 35474 46398 35476 46450
rect 35420 46386 35476 46398
rect 35980 46452 36036 46462
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34412 45106 34692 45108
rect 34412 45054 34414 45106
rect 34466 45054 34692 45106
rect 34412 45052 34692 45054
rect 34412 45042 34468 45052
rect 34188 44996 34244 45006
rect 34188 44902 34244 44940
rect 34636 44546 34692 45052
rect 34748 45106 35140 45108
rect 34748 45054 34750 45106
rect 34802 45054 35140 45106
rect 34748 45052 35140 45054
rect 34748 45042 34804 45052
rect 34636 44494 34638 44546
rect 34690 44494 34692 44546
rect 34636 44482 34692 44494
rect 34076 44434 34132 44446
rect 34076 44382 34078 44434
rect 34130 44382 34132 44434
rect 34076 44324 34132 44382
rect 34076 44268 34468 44324
rect 33964 44212 34020 44222
rect 33964 44118 34020 44156
rect 34076 44100 34132 44110
rect 34076 44006 34132 44044
rect 33852 43820 34356 43876
rect 34188 42530 34244 42542
rect 34188 42478 34190 42530
rect 34242 42478 34244 42530
rect 34188 42308 34244 42478
rect 34188 42242 34244 42252
rect 34188 40180 34244 40190
rect 33740 39396 33796 39406
rect 33740 39058 33796 39340
rect 33740 39006 33742 39058
rect 33794 39006 33796 39058
rect 33740 38994 33796 39006
rect 34188 39058 34244 40124
rect 34188 39006 34190 39058
rect 34242 39006 34244 39058
rect 34188 38994 34244 39006
rect 33964 38834 34020 38846
rect 33964 38782 33966 38834
rect 34018 38782 34020 38834
rect 33964 37716 34020 38782
rect 33964 37650 34020 37660
rect 34076 38722 34132 38734
rect 34076 38670 34078 38722
rect 34130 38670 34132 38722
rect 34076 37492 34132 38670
rect 33740 37436 34132 37492
rect 33740 36706 33796 37436
rect 33740 36654 33742 36706
rect 33794 36654 33796 36706
rect 33740 36642 33796 36654
rect 33852 37154 33908 37166
rect 33852 37102 33854 37154
rect 33906 37102 33908 37154
rect 33852 36594 33908 37102
rect 33852 36542 33854 36594
rect 33906 36542 33908 36594
rect 33852 36530 33908 36542
rect 34300 36596 34356 43820
rect 34412 43650 34468 44268
rect 34524 44210 34580 44222
rect 34524 44158 34526 44210
rect 34578 44158 34580 44210
rect 34524 43988 34580 44158
rect 34636 44100 34692 44110
rect 34636 44006 34692 44044
rect 34524 43922 34580 43932
rect 34412 43598 34414 43650
rect 34466 43598 34468 43650
rect 34412 43586 34468 43598
rect 34636 43650 34692 43662
rect 34636 43598 34638 43650
rect 34690 43598 34692 43650
rect 34524 43316 34580 43326
rect 34524 42978 34580 43260
rect 34524 42926 34526 42978
rect 34578 42926 34580 42978
rect 34524 42914 34580 42926
rect 34636 41188 34692 43598
rect 35084 43538 35140 45052
rect 35420 44996 35476 45006
rect 35420 44902 35476 44940
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35084 43486 35086 43538
rect 35138 43486 35140 43538
rect 35084 43474 35140 43486
rect 34748 43428 34804 43438
rect 34748 43334 34804 43372
rect 35868 43428 35924 43438
rect 35868 43334 35924 43372
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34748 42756 34804 42766
rect 34748 42662 34804 42700
rect 34972 42532 35028 42542
rect 34972 42438 35028 42476
rect 35084 42530 35140 42542
rect 35084 42478 35086 42530
rect 35138 42478 35140 42530
rect 34748 42084 34804 42094
rect 34748 41412 34804 42028
rect 34972 41970 35028 41982
rect 34972 41918 34974 41970
rect 35026 41918 35028 41970
rect 34860 41412 34916 41422
rect 34748 41356 34860 41412
rect 34860 41298 34916 41356
rect 34860 41246 34862 41298
rect 34914 41246 34916 41298
rect 34860 41234 34916 41246
rect 34636 41122 34692 41132
rect 34972 41076 35028 41918
rect 35084 41972 35140 42478
rect 35196 42530 35252 42542
rect 35196 42478 35198 42530
rect 35250 42478 35252 42530
rect 35196 42196 35252 42478
rect 35644 42530 35700 42542
rect 35644 42478 35646 42530
rect 35698 42478 35700 42530
rect 35644 42308 35700 42478
rect 35644 42242 35700 42252
rect 35252 42140 35476 42196
rect 35196 42102 35252 42140
rect 35420 42084 35476 42140
rect 35532 42084 35588 42094
rect 35420 42028 35532 42084
rect 35532 41990 35588 42028
rect 35084 41906 35140 41916
rect 35308 41970 35364 41982
rect 35308 41918 35310 41970
rect 35362 41918 35364 41970
rect 35308 41748 35364 41918
rect 35868 41972 35924 41982
rect 35868 41878 35924 41916
rect 35420 41858 35476 41870
rect 35420 41806 35422 41858
rect 35474 41806 35476 41858
rect 35420 41748 35476 41806
rect 35756 41860 35812 41870
rect 35420 41692 35588 41748
rect 35308 41682 35364 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35532 41412 35588 41692
rect 35308 41356 35588 41412
rect 34972 41010 35028 41020
rect 35084 41300 35140 41310
rect 35084 40402 35140 41244
rect 35308 41186 35364 41356
rect 35308 41134 35310 41186
rect 35362 41134 35364 41186
rect 35308 41122 35364 41134
rect 35756 41186 35812 41804
rect 35756 41134 35758 41186
rect 35810 41134 35812 41186
rect 35756 41122 35812 41134
rect 35084 40350 35086 40402
rect 35138 40350 35140 40402
rect 35084 40338 35140 40350
rect 35420 41074 35476 41086
rect 35420 41022 35422 41074
rect 35474 41022 35476 41074
rect 35420 40180 35476 41022
rect 35644 40962 35700 40974
rect 35644 40910 35646 40962
rect 35698 40910 35700 40962
rect 35644 40516 35700 40910
rect 35756 40516 35812 40526
rect 35644 40514 35812 40516
rect 35644 40462 35758 40514
rect 35810 40462 35812 40514
rect 35644 40460 35812 40462
rect 35756 40450 35812 40460
rect 35420 40114 35476 40124
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35980 39284 36036 46396
rect 36876 44660 36932 49196
rect 37100 49028 37156 49868
rect 37324 49810 37380 49822
rect 37324 49758 37326 49810
rect 37378 49758 37380 49810
rect 37324 49028 37380 49758
rect 37548 49812 37604 49822
rect 37548 49138 37604 49756
rect 37660 49700 37716 50542
rect 37772 49812 37828 51324
rect 37996 50148 38052 51884
rect 38108 51716 38164 51998
rect 38108 51650 38164 51660
rect 38220 52052 38276 52780
rect 38220 51492 38276 51996
rect 38220 51426 38276 51436
rect 38332 50820 38388 53676
rect 38668 53732 38724 53742
rect 38668 53638 38724 53676
rect 38780 53730 38836 53742
rect 38780 53678 38782 53730
rect 38834 53678 38836 53730
rect 38444 53506 38500 53518
rect 38444 53454 38446 53506
rect 38498 53454 38500 53506
rect 38444 53396 38500 53454
rect 38780 53396 38836 53678
rect 38500 53340 38612 53396
rect 38444 53330 38500 53340
rect 38444 52834 38500 52846
rect 38444 52782 38446 52834
rect 38498 52782 38500 52834
rect 38444 52724 38500 52782
rect 38444 52658 38500 52668
rect 38556 52500 38612 53340
rect 38668 53340 38836 53396
rect 38892 53732 38948 53742
rect 38668 53284 38724 53340
rect 38892 53284 38948 53676
rect 38668 53218 38724 53228
rect 38780 53228 38948 53284
rect 38668 52948 38724 52958
rect 38780 52948 38836 53228
rect 39004 53172 39060 54236
rect 39116 54198 39172 54236
rect 39116 53732 39172 53742
rect 39116 53638 39172 53676
rect 39228 53172 39284 54462
rect 39340 53732 39396 55022
rect 39452 54740 39508 59200
rect 39900 56644 39956 59200
rect 40348 56980 40404 59200
rect 40796 57092 40852 59200
rect 41020 57092 41076 57102
rect 40796 57036 41020 57092
rect 41020 57026 41076 57036
rect 40348 56924 40964 56980
rect 40460 56756 40516 56766
rect 39900 56642 40292 56644
rect 39900 56590 39902 56642
rect 39954 56590 40292 56642
rect 39900 56588 40292 56590
rect 39900 56578 39956 56588
rect 39788 56084 39844 56094
rect 39676 56082 39844 56084
rect 39676 56030 39790 56082
rect 39842 56030 39844 56082
rect 39676 56028 39844 56030
rect 39676 55410 39732 56028
rect 39788 56018 39844 56028
rect 39676 55358 39678 55410
rect 39730 55358 39732 55410
rect 39676 55346 39732 55358
rect 39676 54740 39732 54750
rect 39452 54738 39732 54740
rect 39452 54686 39678 54738
rect 39730 54686 39732 54738
rect 39452 54684 39732 54686
rect 39676 54674 39732 54684
rect 40236 54738 40292 56588
rect 40460 55970 40516 56700
rect 40460 55918 40462 55970
rect 40514 55918 40516 55970
rect 40460 55906 40516 55918
rect 40236 54686 40238 54738
rect 40290 54686 40292 54738
rect 40236 54674 40292 54686
rect 40908 54738 40964 56924
rect 41692 56308 41748 59200
rect 42140 56980 42196 59200
rect 42140 56914 42196 56924
rect 42924 57092 42980 57102
rect 41692 56242 41748 56252
rect 42028 56868 42084 56878
rect 42028 55970 42084 56812
rect 42588 56084 42644 56094
rect 42588 56082 42756 56084
rect 42588 56030 42590 56082
rect 42642 56030 42756 56082
rect 42588 56028 42756 56030
rect 42588 56018 42644 56028
rect 42028 55918 42030 55970
rect 42082 55918 42084 55970
rect 42028 55906 42084 55918
rect 42588 55298 42644 55310
rect 42588 55246 42590 55298
rect 42642 55246 42644 55298
rect 41804 55188 41860 55198
rect 41804 55094 41860 55132
rect 40908 54686 40910 54738
rect 40962 54686 40964 54738
rect 40908 54674 40964 54686
rect 39452 54292 39508 54302
rect 39508 54236 39732 54292
rect 39452 54226 39508 54236
rect 39564 53844 39620 53854
rect 39564 53750 39620 53788
rect 39340 53666 39396 53676
rect 39452 53620 39508 53630
rect 39452 53526 39508 53564
rect 39676 53618 39732 54236
rect 41804 53732 41860 53742
rect 39676 53566 39678 53618
rect 39730 53566 39732 53618
rect 39676 53554 39732 53566
rect 39788 53618 39844 53630
rect 39788 53566 39790 53618
rect 39842 53566 39844 53618
rect 39004 53116 39172 53172
rect 38668 52946 38836 52948
rect 38668 52894 38670 52946
rect 38722 52894 38836 52946
rect 38668 52892 38836 52894
rect 38668 52882 38724 52892
rect 38556 52444 38724 52500
rect 38444 52276 38500 52286
rect 38444 52182 38500 52220
rect 38556 52050 38612 52062
rect 38556 51998 38558 52050
rect 38610 51998 38612 52050
rect 38556 51828 38612 51998
rect 38668 52052 38724 52444
rect 38780 52388 38836 52892
rect 38892 53058 38948 53070
rect 38892 53006 38894 53058
rect 38946 53006 38948 53058
rect 38892 52836 38948 53006
rect 38892 52770 38948 52780
rect 39004 52946 39060 52958
rect 39004 52894 39006 52946
rect 39058 52894 39060 52946
rect 38892 52388 38948 52398
rect 38780 52332 38892 52388
rect 38892 52322 38948 52332
rect 39004 52164 39060 52894
rect 38892 52108 39060 52164
rect 38780 52052 38836 52062
rect 38668 51996 38780 52052
rect 38780 51958 38836 51996
rect 38780 51828 38836 51838
rect 38556 51772 38780 51828
rect 38780 51762 38836 51772
rect 38556 51604 38612 51614
rect 38892 51604 38948 52108
rect 38556 51510 38612 51548
rect 38780 51548 38948 51604
rect 39004 51938 39060 51950
rect 39004 51886 39006 51938
rect 39058 51886 39060 51938
rect 38444 51492 38500 51502
rect 38444 51398 38500 51436
rect 38668 51490 38724 51502
rect 38668 51438 38670 51490
rect 38722 51438 38724 51490
rect 38220 50708 38276 50718
rect 38220 50594 38276 50652
rect 38220 50542 38222 50594
rect 38274 50542 38276 50594
rect 38220 50484 38276 50542
rect 38220 50418 38276 50428
rect 38332 50484 38388 50764
rect 38444 50484 38500 50494
rect 38332 50482 38444 50484
rect 38332 50430 38334 50482
rect 38386 50430 38444 50482
rect 38332 50428 38444 50430
rect 38332 50418 38388 50428
rect 38444 50418 38500 50428
rect 38668 50484 38724 51438
rect 38668 50418 38724 50428
rect 38780 51434 38836 51548
rect 38780 51382 38782 51434
rect 38834 51382 38836 51434
rect 37996 50082 38052 50092
rect 38668 50036 38724 50046
rect 37884 49812 37940 49822
rect 38668 49812 38724 49980
rect 37772 49810 37940 49812
rect 37772 49758 37886 49810
rect 37938 49758 37940 49810
rect 37772 49756 37940 49758
rect 37884 49746 37940 49756
rect 38332 49810 38724 49812
rect 38332 49758 38670 49810
rect 38722 49758 38724 49810
rect 38332 49756 38724 49758
rect 37660 49644 37828 49700
rect 37548 49086 37550 49138
rect 37602 49086 37604 49138
rect 37548 49074 37604 49086
rect 37436 49028 37492 49038
rect 37324 48972 37436 49028
rect 37100 48934 37156 48972
rect 37436 48934 37492 48972
rect 37660 48916 37716 48926
rect 37660 48822 37716 48860
rect 37772 48804 37828 49644
rect 38332 49026 38388 49756
rect 38668 49746 38724 49756
rect 38668 49588 38724 49598
rect 38780 49588 38836 51382
rect 39004 51268 39060 51886
rect 39004 51202 39060 51212
rect 38668 49586 38836 49588
rect 38668 49534 38670 49586
rect 38722 49534 38836 49586
rect 38668 49532 38836 49534
rect 38892 51156 38948 51166
rect 38668 49522 38724 49532
rect 38892 49252 38948 51100
rect 39116 51044 39172 53116
rect 39228 53106 39284 53116
rect 39340 53508 39396 53518
rect 39228 52724 39284 52734
rect 39228 51378 39284 52668
rect 39340 52386 39396 53452
rect 39564 53508 39620 53518
rect 39452 53172 39508 53182
rect 39564 53172 39620 53452
rect 39788 53396 39844 53566
rect 39900 53618 39956 53630
rect 39900 53566 39902 53618
rect 39954 53566 39956 53618
rect 39900 53508 39956 53566
rect 39900 53442 39956 53452
rect 39788 53330 39844 53340
rect 40908 53284 40964 53294
rect 39452 53170 39620 53172
rect 39452 53118 39454 53170
rect 39506 53118 39620 53170
rect 39452 53116 39620 53118
rect 40236 53172 40292 53182
rect 39452 53106 39508 53116
rect 40236 53058 40292 53116
rect 40236 53006 40238 53058
rect 40290 53006 40292 53058
rect 39788 52948 39844 52958
rect 39676 52836 39732 52846
rect 39676 52742 39732 52780
rect 39340 52334 39342 52386
rect 39394 52334 39396 52386
rect 39340 52322 39396 52334
rect 39452 52164 39508 52202
rect 39452 52098 39508 52108
rect 39788 52050 39844 52892
rect 40012 52722 40068 52734
rect 40012 52670 40014 52722
rect 40066 52670 40068 52722
rect 40012 52164 40068 52670
rect 40012 52098 40068 52108
rect 40124 52164 40180 52174
rect 40236 52164 40292 53006
rect 40908 52948 40964 53228
rect 41020 53172 41076 53182
rect 41020 53170 41300 53172
rect 41020 53118 41022 53170
rect 41074 53118 41300 53170
rect 41020 53116 41300 53118
rect 41020 53106 41076 53116
rect 41132 52948 41188 52958
rect 40908 52892 41132 52948
rect 41132 52854 41188 52892
rect 41020 52724 41076 52734
rect 41020 52630 41076 52668
rect 40796 52388 40852 52398
rect 41244 52388 41300 53116
rect 41804 53060 41860 53676
rect 42252 53732 42308 53742
rect 42252 53638 42308 53676
rect 42588 53732 42644 55246
rect 42700 54402 42756 56028
rect 42924 55970 42980 57036
rect 43036 56196 43092 59200
rect 43036 56140 43428 56196
rect 42924 55918 42926 55970
rect 42978 55918 42980 55970
rect 42924 55906 42980 55918
rect 42924 55188 42980 55198
rect 42924 55094 42980 55132
rect 43036 55186 43092 55198
rect 43036 55134 43038 55186
rect 43090 55134 43092 55186
rect 42700 54350 42702 54402
rect 42754 54350 42756 54402
rect 42700 54338 42756 54350
rect 43036 54292 43092 55134
rect 43372 55186 43428 56140
rect 43484 55972 43540 59200
rect 44380 57090 44436 59200
rect 44380 57038 44382 57090
rect 44434 57038 44436 57090
rect 44380 57026 44436 57038
rect 44044 56980 44100 56990
rect 43596 56308 43652 56318
rect 43596 56214 43652 56252
rect 43484 55906 43540 55916
rect 44044 55970 44100 56924
rect 44044 55918 44046 55970
rect 44098 55918 44100 55970
rect 44044 55906 44100 55918
rect 44492 55972 44548 55982
rect 44492 55878 44548 55916
rect 44828 55860 44884 59200
rect 44940 57090 44996 57102
rect 44940 57038 44942 57090
rect 44994 57038 44996 57090
rect 44940 56306 44996 57038
rect 44940 56254 44942 56306
rect 44994 56254 44996 56306
rect 44940 56242 44996 56254
rect 45724 56308 45780 59200
rect 45948 56308 46004 56318
rect 45724 56306 46004 56308
rect 45724 56254 45950 56306
rect 46002 56254 46004 56306
rect 45724 56252 46004 56254
rect 45948 56242 46004 56252
rect 46172 55972 46228 59200
rect 47068 57764 47124 59200
rect 47068 57708 47460 57764
rect 47404 56306 47460 57708
rect 47404 56254 47406 56306
rect 47458 56254 47460 56306
rect 47404 56242 47460 56254
rect 46396 55972 46452 55982
rect 46172 55970 46452 55972
rect 46172 55918 46398 55970
rect 46450 55918 46452 55970
rect 46172 55916 46452 55918
rect 47516 55972 47572 59200
rect 48412 56308 48468 59200
rect 48636 56308 48692 56318
rect 48412 56306 48692 56308
rect 48412 56254 48638 56306
rect 48690 56254 48692 56306
rect 48412 56252 48692 56254
rect 48636 56242 48692 56252
rect 47852 55972 47908 55982
rect 47516 55970 47908 55972
rect 47516 55918 47854 55970
rect 47906 55918 47908 55970
rect 47516 55916 47908 55918
rect 48860 55972 48916 59200
rect 49756 56308 49812 59200
rect 49980 56308 50036 56318
rect 49756 56306 50036 56308
rect 49756 56254 49982 56306
rect 50034 56254 50036 56306
rect 49756 56252 50036 56254
rect 49980 56242 50036 56252
rect 49084 55972 49140 55982
rect 48860 55970 49140 55972
rect 48860 55918 49086 55970
rect 49138 55918 49140 55970
rect 48860 55916 49140 55918
rect 50204 55972 50260 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 51100 56308 51156 59200
rect 51324 56308 51380 56318
rect 51100 56306 51380 56308
rect 51100 56254 51326 56306
rect 51378 56254 51380 56306
rect 51100 56252 51380 56254
rect 51324 56242 51380 56252
rect 50428 55972 50484 55982
rect 50204 55970 50484 55972
rect 50204 55918 50430 55970
rect 50482 55918 50484 55970
rect 50204 55916 50484 55918
rect 51548 55972 51604 59200
rect 52444 56308 52500 59200
rect 52668 56308 52724 56318
rect 52444 56306 52724 56308
rect 52444 56254 52670 56306
rect 52722 56254 52724 56306
rect 52444 56252 52724 56254
rect 52668 56242 52724 56252
rect 51772 55972 51828 55982
rect 51548 55970 51828 55972
rect 51548 55918 51774 55970
rect 51826 55918 51828 55970
rect 51548 55916 51828 55918
rect 52892 55972 52948 59200
rect 53788 56308 53844 59200
rect 54236 56642 54292 59200
rect 54236 56590 54238 56642
rect 54290 56590 54292 56642
rect 54236 56578 54292 56590
rect 55020 56642 55076 56654
rect 55020 56590 55022 56642
rect 55074 56590 55076 56642
rect 54012 56308 54068 56318
rect 53788 56306 54068 56308
rect 53788 56254 54014 56306
rect 54066 56254 54068 56306
rect 53788 56252 54068 56254
rect 54012 56242 54068 56252
rect 53116 55972 53172 55982
rect 52892 55970 53172 55972
rect 52892 55918 53118 55970
rect 53170 55918 53172 55970
rect 52892 55916 53172 55918
rect 46396 55906 46452 55916
rect 47852 55906 47908 55916
rect 49084 55906 49140 55916
rect 50428 55906 50484 55916
rect 51772 55906 51828 55916
rect 53116 55906 53172 55916
rect 55020 55970 55076 56590
rect 55132 56308 55188 59200
rect 55580 57540 55636 59200
rect 55580 57484 55972 57540
rect 55468 56308 55524 56318
rect 55132 56306 55524 56308
rect 55132 56254 55470 56306
rect 55522 56254 55524 56306
rect 55132 56252 55524 56254
rect 55468 56242 55524 56252
rect 55020 55918 55022 55970
rect 55074 55918 55076 55970
rect 55020 55906 55076 55918
rect 55916 55970 55972 57484
rect 55916 55918 55918 55970
rect 55970 55918 55972 55970
rect 55916 55906 55972 55918
rect 44828 55794 44884 55804
rect 45388 55860 45444 55870
rect 45388 55766 45444 55804
rect 43372 55134 43374 55186
rect 43426 55134 43428 55186
rect 43372 55122 43428 55134
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 45500 54514 45556 54526
rect 45500 54462 45502 54514
rect 45554 54462 45556 54514
rect 44828 54402 44884 54414
rect 44828 54350 44830 54402
rect 44882 54350 44884 54402
rect 43036 54226 43092 54236
rect 43708 54292 43764 54302
rect 42588 53666 42644 53676
rect 42812 53730 42868 53742
rect 42812 53678 42814 53730
rect 42866 53678 42868 53730
rect 42140 53172 42196 53182
rect 42140 53078 42196 53116
rect 42588 53172 42644 53182
rect 42588 53078 42644 53116
rect 40796 52294 40852 52332
rect 40908 52386 41300 52388
rect 40908 52334 41246 52386
rect 41298 52334 41300 52386
rect 40908 52332 41300 52334
rect 40124 52162 40292 52164
rect 40124 52110 40126 52162
rect 40178 52110 40292 52162
rect 40124 52108 40292 52110
rect 40908 52162 40964 52332
rect 40908 52110 40910 52162
rect 40962 52110 40964 52162
rect 40124 52098 40180 52108
rect 40908 52098 40964 52110
rect 39788 51998 39790 52050
rect 39842 51998 39844 52050
rect 39788 51986 39844 51998
rect 39228 51326 39230 51378
rect 39282 51326 39284 51378
rect 39228 51314 39284 51326
rect 39452 51940 39508 51950
rect 39452 51378 39508 51884
rect 40796 51938 40852 51950
rect 40796 51886 40798 51938
rect 40850 51886 40852 51938
rect 40124 51828 40180 51838
rect 40012 51492 40068 51502
rect 40124 51492 40180 51772
rect 40012 51490 40180 51492
rect 40012 51438 40014 51490
rect 40066 51438 40180 51490
rect 40012 51436 40180 51438
rect 40012 51426 40068 51436
rect 39452 51326 39454 51378
rect 39506 51326 39508 51378
rect 39452 51314 39508 51326
rect 39788 51378 39844 51390
rect 39788 51326 39790 51378
rect 39842 51326 39844 51378
rect 39676 51268 39732 51278
rect 39676 51174 39732 51212
rect 39004 50988 39172 51044
rect 39004 50820 39060 50988
rect 39004 50482 39060 50764
rect 39228 50708 39284 50746
rect 39452 50708 39508 50718
rect 39788 50708 39844 51326
rect 39228 50642 39284 50652
rect 39340 50652 39452 50708
rect 39508 50652 39844 50708
rect 39116 50596 39172 50606
rect 39116 50502 39172 50540
rect 39004 50430 39006 50482
rect 39058 50430 39060 50482
rect 39004 50418 39060 50430
rect 39228 50484 39284 50494
rect 39116 50148 39172 50158
rect 39228 50148 39284 50428
rect 39340 50482 39396 50652
rect 39452 50614 39508 50652
rect 39900 50596 39956 50606
rect 39340 50430 39342 50482
rect 39394 50430 39396 50482
rect 39340 50418 39396 50430
rect 39788 50594 39956 50596
rect 39788 50542 39902 50594
rect 39954 50542 39956 50594
rect 39788 50540 39956 50542
rect 39564 50372 39620 50382
rect 39788 50372 39844 50540
rect 39900 50530 39956 50540
rect 40124 50482 40180 51436
rect 40796 51268 40852 51886
rect 41132 51940 41188 52332
rect 41244 52322 41300 52332
rect 41580 53058 41860 53060
rect 41580 53006 41806 53058
rect 41858 53006 41860 53058
rect 41580 53004 41860 53006
rect 41580 52276 41636 53004
rect 41804 52994 41860 53004
rect 41916 52948 41972 52958
rect 41356 52220 41636 52276
rect 41804 52276 41860 52286
rect 41244 52164 41300 52174
rect 41356 52164 41412 52220
rect 41804 52182 41860 52220
rect 41244 52162 41412 52164
rect 41244 52110 41246 52162
rect 41298 52110 41412 52162
rect 41244 52108 41412 52110
rect 41244 52098 41300 52108
rect 41580 52052 41636 52062
rect 41580 51958 41636 51996
rect 41132 51884 41524 51940
rect 41468 51378 41524 51884
rect 41468 51326 41470 51378
rect 41522 51326 41524 51378
rect 41468 51314 41524 51326
rect 41916 51716 41972 52892
rect 42476 52946 42532 52958
rect 42476 52894 42478 52946
rect 42530 52894 42532 52946
rect 41244 51268 41300 51278
rect 40796 51266 41300 51268
rect 40796 51214 41246 51266
rect 41298 51214 41300 51266
rect 40796 51212 41300 51214
rect 41244 51156 41300 51212
rect 41244 51090 41300 51100
rect 41804 51154 41860 51166
rect 41804 51102 41806 51154
rect 41858 51102 41860 51154
rect 41692 50932 41748 50942
rect 41580 50708 41636 50718
rect 40908 50596 40964 50606
rect 40124 50430 40126 50482
rect 40178 50430 40180 50482
rect 40124 50418 40180 50430
rect 40236 50484 40292 50494
rect 40684 50482 40740 50494
rect 40684 50430 40686 50482
rect 40738 50430 40740 50482
rect 40684 50428 40740 50430
rect 39564 50370 39844 50372
rect 39564 50318 39566 50370
rect 39618 50318 39844 50370
rect 39564 50316 39844 50318
rect 39564 50306 39620 50316
rect 39172 50092 39284 50148
rect 39116 50082 39172 50092
rect 39116 49922 39172 49934
rect 39116 49870 39118 49922
rect 39170 49870 39172 49922
rect 39116 49812 39172 49870
rect 39116 49746 39172 49756
rect 39228 49810 39284 50092
rect 39788 50034 39844 50316
rect 40012 50372 40068 50382
rect 40012 50278 40068 50316
rect 40236 50372 40740 50428
rect 39788 49982 39790 50034
rect 39842 49982 39844 50034
rect 39788 49970 39844 49982
rect 40012 50036 40068 50046
rect 39228 49758 39230 49810
rect 39282 49758 39284 49810
rect 39228 49746 39284 49758
rect 39900 49812 39956 49822
rect 39676 49586 39732 49598
rect 39676 49534 39678 49586
rect 39730 49534 39732 49586
rect 39004 49252 39060 49262
rect 39676 49252 39732 49534
rect 38892 49250 39732 49252
rect 38892 49198 39006 49250
rect 39058 49198 39732 49250
rect 38892 49196 39732 49198
rect 39788 49252 39844 49262
rect 39004 49186 39060 49196
rect 38332 48974 38334 49026
rect 38386 48974 38388 49026
rect 38332 48916 38388 48974
rect 39116 49028 39172 49038
rect 39116 48934 39172 48972
rect 39788 49028 39844 49196
rect 39788 48934 39844 48972
rect 38332 48850 38388 48860
rect 39452 48916 39508 48926
rect 39452 48822 39508 48860
rect 39900 48916 39956 49756
rect 40012 49810 40068 49980
rect 40012 49758 40014 49810
rect 40066 49758 40068 49810
rect 40012 49746 40068 49758
rect 40236 49138 40292 50372
rect 40908 50034 40964 50540
rect 40908 49982 40910 50034
rect 40962 49982 40964 50034
rect 40908 49970 40964 49982
rect 41356 50370 41412 50382
rect 41356 50318 41358 50370
rect 41410 50318 41412 50370
rect 41356 50036 41412 50318
rect 41356 49970 41412 49980
rect 41244 49810 41300 49822
rect 41244 49758 41246 49810
rect 41298 49758 41300 49810
rect 40236 49086 40238 49138
rect 40290 49086 40292 49138
rect 40236 49074 40292 49086
rect 40684 49700 40740 49710
rect 40684 49026 40740 49644
rect 41244 49700 41300 49758
rect 41244 49634 41300 49644
rect 40684 48974 40686 49026
rect 40738 48974 40740 49026
rect 40684 48962 40740 48974
rect 41356 49588 41412 49598
rect 41356 49026 41412 49532
rect 41356 48974 41358 49026
rect 41410 48974 41412 49026
rect 41356 48962 41412 48974
rect 39900 48850 39956 48860
rect 41580 48914 41636 50652
rect 41692 50594 41748 50876
rect 41692 50542 41694 50594
rect 41746 50542 41748 50594
rect 41692 50530 41748 50542
rect 41804 50428 41860 51102
rect 41916 50820 41972 51660
rect 42028 52164 42084 52174
rect 42028 51490 42084 52108
rect 42140 52050 42196 52062
rect 42140 51998 42142 52050
rect 42194 51998 42196 52050
rect 42140 51828 42196 51998
rect 42140 51762 42196 51772
rect 42028 51438 42030 51490
rect 42082 51438 42084 51490
rect 42028 51426 42084 51438
rect 42252 51380 42308 51390
rect 42476 51380 42532 52894
rect 42252 51378 42532 51380
rect 42252 51326 42254 51378
rect 42306 51326 42532 51378
rect 42252 51324 42532 51326
rect 42588 52722 42644 52734
rect 42588 52670 42590 52722
rect 42642 52670 42644 52722
rect 42252 51156 42308 51324
rect 42252 51090 42308 51100
rect 42364 50932 42420 50942
rect 41916 50764 42308 50820
rect 42252 50706 42308 50764
rect 42252 50654 42254 50706
rect 42306 50654 42308 50706
rect 42252 50642 42308 50654
rect 41692 50372 41860 50428
rect 41916 50596 41972 50606
rect 41692 49028 41748 50372
rect 41916 50034 41972 50540
rect 42140 50596 42196 50606
rect 41916 49982 41918 50034
rect 41970 49982 41972 50034
rect 41916 49970 41972 49982
rect 42028 50482 42084 50494
rect 42028 50430 42030 50482
rect 42082 50430 42084 50482
rect 42028 49812 42084 50430
rect 42028 49746 42084 49756
rect 42140 49812 42196 50540
rect 42364 50596 42420 50876
rect 42588 50820 42644 52670
rect 42700 52052 42756 52062
rect 42700 51492 42756 51996
rect 42812 51828 42868 53678
rect 43372 53620 43428 53630
rect 43036 53618 43428 53620
rect 43036 53566 43374 53618
rect 43426 53566 43428 53618
rect 43036 53564 43428 53566
rect 43036 53058 43092 53564
rect 43372 53554 43428 53564
rect 43708 53618 43764 54236
rect 44828 54292 44884 54350
rect 44828 54226 44884 54236
rect 43708 53566 43710 53618
rect 43762 53566 43764 53618
rect 43708 53554 43764 53566
rect 45052 53732 45108 53742
rect 43036 53006 43038 53058
rect 43090 53006 43092 53058
rect 43036 52994 43092 53006
rect 42812 51762 42868 51772
rect 43484 52946 43540 52958
rect 43484 52894 43486 52946
rect 43538 52894 43540 52946
rect 43484 51828 43540 52894
rect 43932 52948 43988 52958
rect 43484 51762 43540 51772
rect 43820 51940 43876 51950
rect 42700 51490 42868 51492
rect 42700 51438 42702 51490
rect 42754 51438 42868 51490
rect 42700 51436 42868 51438
rect 42700 51426 42756 51436
rect 42700 50820 42756 50830
rect 42588 50818 42756 50820
rect 42588 50766 42702 50818
rect 42754 50766 42756 50818
rect 42588 50764 42756 50766
rect 42700 50754 42756 50764
rect 42700 50596 42756 50606
rect 42364 50594 42700 50596
rect 42364 50542 42366 50594
rect 42418 50542 42700 50594
rect 42364 50540 42700 50542
rect 42364 50530 42420 50540
rect 42700 50530 42756 50540
rect 42812 50484 42868 51436
rect 42924 51490 42980 51502
rect 42924 51438 42926 51490
rect 42978 51438 42980 51490
rect 42924 50708 42980 51438
rect 43708 51490 43764 51502
rect 43708 51438 43710 51490
rect 43762 51438 43764 51490
rect 43596 51380 43652 51390
rect 42924 50642 42980 50652
rect 43036 51378 43652 51380
rect 43036 51326 43598 51378
rect 43650 51326 43652 51378
rect 43036 51324 43652 51326
rect 43036 50818 43092 51324
rect 43596 51314 43652 51324
rect 43708 51380 43764 51438
rect 43708 51314 43764 51324
rect 43036 50766 43038 50818
rect 43090 50766 43092 50818
rect 42924 50484 42980 50522
rect 42812 50428 42924 50484
rect 42924 50418 42980 50428
rect 42364 50372 42420 50382
rect 42140 49810 42308 49812
rect 42140 49758 42142 49810
rect 42194 49758 42308 49810
rect 42140 49756 42308 49758
rect 42140 49746 42196 49756
rect 41804 49586 41860 49598
rect 41804 49534 41806 49586
rect 41858 49534 41860 49586
rect 41804 49252 41860 49534
rect 41804 49186 41860 49196
rect 42028 49028 42084 49038
rect 41692 49026 42084 49028
rect 41692 48974 41694 49026
rect 41746 48974 42030 49026
rect 42082 48974 42084 49026
rect 41692 48972 42084 48974
rect 41692 48962 41748 48972
rect 42028 48962 42084 48972
rect 41580 48862 41582 48914
rect 41634 48862 41636 48914
rect 41580 48850 41636 48862
rect 42140 48916 42196 48926
rect 42252 48916 42308 49756
rect 42364 49026 42420 50316
rect 43036 50148 43092 50766
rect 43372 51156 43428 51166
rect 43372 50482 43428 51100
rect 43708 51156 43764 51166
rect 43820 51156 43876 51884
rect 43708 51154 43876 51156
rect 43708 51102 43710 51154
rect 43762 51102 43876 51154
rect 43708 51100 43876 51102
rect 43708 51090 43764 51100
rect 43596 50820 43652 50830
rect 43596 50596 43652 50764
rect 43372 50430 43374 50482
rect 43426 50430 43428 50482
rect 43372 50418 43428 50430
rect 43484 50594 43652 50596
rect 43484 50542 43598 50594
rect 43650 50542 43652 50594
rect 43484 50540 43652 50542
rect 43036 50082 43092 50092
rect 43484 50036 43540 50540
rect 43596 50530 43652 50540
rect 43932 50428 43988 52892
rect 45052 52946 45108 53676
rect 45500 53732 45556 54462
rect 45948 53844 46004 53854
rect 51548 53844 51604 53854
rect 45500 53666 45556 53676
rect 45724 53842 46004 53844
rect 45724 53790 45950 53842
rect 46002 53790 46004 53842
rect 45724 53788 46004 53790
rect 45724 53058 45780 53788
rect 45948 53778 46004 53788
rect 51436 53842 51604 53844
rect 51436 53790 51550 53842
rect 51602 53790 51604 53842
rect 51436 53788 51604 53790
rect 46956 53732 47012 53742
rect 46284 53620 46340 53630
rect 46284 53526 46340 53564
rect 46060 53508 46116 53518
rect 45724 53006 45726 53058
rect 45778 53006 45780 53058
rect 45724 52994 45780 53006
rect 45948 53506 46116 53508
rect 45948 53454 46062 53506
rect 46114 53454 46116 53506
rect 45948 53452 46116 53454
rect 45052 52894 45054 52946
rect 45106 52894 45108 52946
rect 45052 52882 45108 52894
rect 45948 52948 46004 53452
rect 46060 53442 46116 53452
rect 46004 52892 46228 52948
rect 45948 52882 46004 52892
rect 46172 52276 46228 52892
rect 46060 52274 46228 52276
rect 46060 52222 46174 52274
rect 46226 52222 46228 52274
rect 46060 52220 46228 52222
rect 45052 51380 45108 51390
rect 45052 50818 45108 51324
rect 45612 51268 45668 51278
rect 45052 50766 45054 50818
rect 45106 50766 45108 50818
rect 45052 50754 45108 50766
rect 45388 51212 45612 51268
rect 45388 50818 45444 51212
rect 45612 51174 45668 51212
rect 45836 51156 45892 51166
rect 45836 51062 45892 51100
rect 45388 50766 45390 50818
rect 45442 50766 45444 50818
rect 45388 50754 45444 50766
rect 46060 50594 46116 52220
rect 46172 52210 46228 52220
rect 46732 51940 46788 51950
rect 46396 51492 46452 51502
rect 46396 51378 46452 51436
rect 46396 51326 46398 51378
rect 46450 51326 46452 51378
rect 46396 51314 46452 51326
rect 46620 51266 46676 51278
rect 46620 51214 46622 51266
rect 46674 51214 46676 51266
rect 46172 51156 46228 51166
rect 46172 51154 46564 51156
rect 46172 51102 46174 51154
rect 46226 51102 46564 51154
rect 46172 51100 46564 51102
rect 46172 51090 46228 51100
rect 46060 50542 46062 50594
rect 46114 50542 46116 50594
rect 46060 50530 46116 50542
rect 46508 50596 46564 51100
rect 46620 50820 46676 51214
rect 46732 51156 46788 51884
rect 46732 51090 46788 51100
rect 46844 51378 46900 51390
rect 46844 51326 46846 51378
rect 46898 51326 46900 51378
rect 46620 50754 46676 50764
rect 46620 50596 46676 50606
rect 46508 50594 46676 50596
rect 46508 50542 46622 50594
rect 46674 50542 46676 50594
rect 46508 50540 46676 50542
rect 46620 50530 46676 50540
rect 46172 50484 46228 50522
rect 43260 49980 43540 50036
rect 43596 50372 43652 50382
rect 43932 50372 44100 50428
rect 46172 50418 46228 50428
rect 43596 50034 43652 50316
rect 43596 49982 43598 50034
rect 43650 49982 43652 50034
rect 43036 49922 43092 49934
rect 43036 49870 43038 49922
rect 43090 49870 43092 49922
rect 43036 49812 43092 49870
rect 43260 49922 43316 49980
rect 43596 49970 43652 49982
rect 43260 49870 43262 49922
rect 43314 49870 43316 49922
rect 43260 49858 43316 49870
rect 43036 49746 43092 49756
rect 43932 49812 43988 49822
rect 43932 49718 43988 49756
rect 42924 49700 42980 49710
rect 42924 49606 42980 49644
rect 43036 49252 43092 49262
rect 43036 49158 43092 49196
rect 42364 48974 42366 49026
rect 42418 48974 42420 49026
rect 42364 48962 42420 48974
rect 43372 49026 43428 49038
rect 43372 48974 43374 49026
rect 43426 48974 43428 49026
rect 42140 48914 42308 48916
rect 42140 48862 42142 48914
rect 42194 48862 42308 48914
rect 42140 48860 42308 48862
rect 42140 48850 42196 48860
rect 37996 48804 38052 48814
rect 37772 48748 37996 48804
rect 37996 48710 38052 48748
rect 43372 48468 43428 48974
rect 44044 49026 44100 50372
rect 45388 49810 45444 49822
rect 45388 49758 45390 49810
rect 45442 49758 45444 49810
rect 44492 49700 44548 49710
rect 44492 49606 44548 49644
rect 44940 49700 44996 49710
rect 44940 49606 44996 49644
rect 45388 49700 45444 49758
rect 44044 48974 44046 49026
rect 44098 48974 44100 49026
rect 44044 48962 44100 48974
rect 44828 49138 44884 49150
rect 44828 49086 44830 49138
rect 44882 49086 44884 49138
rect 44156 48914 44212 48926
rect 44156 48862 44158 48914
rect 44210 48862 44212 48914
rect 43372 48402 43428 48412
rect 43820 48692 43876 48702
rect 43260 48356 43316 48366
rect 43148 48354 43316 48356
rect 43148 48302 43262 48354
rect 43314 48302 43316 48354
rect 43148 48300 43316 48302
rect 41468 47458 41524 47470
rect 41468 47406 41470 47458
rect 41522 47406 41524 47458
rect 37100 47234 37156 47246
rect 37100 47182 37102 47234
rect 37154 47182 37156 47234
rect 37100 47012 37156 47182
rect 39228 47124 39284 47134
rect 37100 46946 37156 46956
rect 37772 47012 37828 47022
rect 37100 46562 37156 46574
rect 37100 46510 37102 46562
rect 37154 46510 37156 46562
rect 37100 46452 37156 46510
rect 37100 46386 37156 46396
rect 37548 45892 37604 45902
rect 37548 44994 37604 45836
rect 37548 44942 37550 44994
rect 37602 44942 37604 44994
rect 37548 44930 37604 44942
rect 36876 44594 36932 44604
rect 37772 44434 37828 46956
rect 39228 46562 39284 47068
rect 39676 46676 39732 46686
rect 40012 46676 40068 46686
rect 39732 46674 40068 46676
rect 39732 46622 40014 46674
rect 40066 46622 40068 46674
rect 39732 46620 40068 46622
rect 39676 46582 39732 46620
rect 40012 46610 40068 46620
rect 41020 46676 41076 46686
rect 41468 46676 41524 47406
rect 42140 47348 42196 47358
rect 42140 47254 42196 47292
rect 43148 47124 43204 48300
rect 43260 48290 43316 48300
rect 43372 48244 43428 48254
rect 43372 48150 43428 48188
rect 43820 48242 43876 48636
rect 44044 48356 44100 48366
rect 44044 48262 44100 48300
rect 43820 48190 43822 48242
rect 43874 48190 43876 48242
rect 43820 48178 43876 48190
rect 44156 48244 44212 48862
rect 44828 48692 44884 49086
rect 44828 48626 44884 48636
rect 43260 48020 43316 48030
rect 43260 47926 43316 47964
rect 44156 47572 44212 48188
rect 44492 48354 44548 48366
rect 44492 48302 44494 48354
rect 44546 48302 44548 48354
rect 44268 47572 44324 47582
rect 44156 47516 44268 47572
rect 44268 47478 44324 47516
rect 43260 47124 43316 47134
rect 43148 47068 43260 47124
rect 43260 47058 43316 47068
rect 44492 47124 44548 48302
rect 44604 48244 44660 48254
rect 44604 48242 45220 48244
rect 44604 48190 44606 48242
rect 44658 48190 45220 48242
rect 44604 48188 45220 48190
rect 44604 48178 44660 48188
rect 41020 46674 41524 46676
rect 41020 46622 41022 46674
rect 41074 46622 41524 46674
rect 41020 46620 41524 46622
rect 41020 46610 41076 46620
rect 39228 46510 39230 46562
rect 39282 46510 39284 46562
rect 39228 46498 39284 46510
rect 40236 46564 40292 46574
rect 40236 46470 40292 46508
rect 40348 46450 40404 46462
rect 40348 46398 40350 46450
rect 40402 46398 40404 46450
rect 39564 46002 39620 46014
rect 39564 45950 39566 46002
rect 39618 45950 39620 46002
rect 38332 45892 38388 45902
rect 38332 45106 38388 45836
rect 39228 45892 39284 45902
rect 39228 45798 39284 45836
rect 39564 45444 39620 45950
rect 40236 46004 40292 46014
rect 40348 46004 40404 46398
rect 40236 46002 40404 46004
rect 40236 45950 40238 46002
rect 40290 45950 40404 46002
rect 40236 45948 40404 45950
rect 40236 45938 40292 45948
rect 39900 45892 39956 45902
rect 39564 45378 39620 45388
rect 39788 45836 39900 45892
rect 39676 45332 39732 45342
rect 39788 45332 39844 45836
rect 39900 45798 39956 45836
rect 40460 45892 40516 45902
rect 40460 45798 40516 45836
rect 40908 45890 40964 45902
rect 41468 45892 41524 46620
rect 44492 46674 44548 47068
rect 44492 46622 44494 46674
rect 44546 46622 44548 46674
rect 44492 46610 44548 46622
rect 44716 48018 44772 48030
rect 44716 47966 44718 48018
rect 44770 47966 44772 48018
rect 44716 47572 44772 47966
rect 45164 47682 45220 48188
rect 45388 48242 45444 49644
rect 46844 49252 46900 51326
rect 46956 51380 47012 53676
rect 48748 53732 48804 53742
rect 48748 53638 48804 53676
rect 48860 53620 48916 53630
rect 49420 53620 49476 53630
rect 48860 52946 48916 53564
rect 49084 53618 49476 53620
rect 49084 53566 49422 53618
rect 49474 53566 49476 53618
rect 49084 53564 49476 53566
rect 49084 53170 49140 53564
rect 49420 53554 49476 53564
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 49084 53118 49086 53170
rect 49138 53118 49140 53170
rect 49084 53106 49140 53118
rect 48860 52894 48862 52946
rect 48914 52894 48916 52946
rect 47852 52834 47908 52846
rect 47852 52782 47854 52834
rect 47906 52782 47908 52834
rect 47404 52164 47460 52174
rect 47852 52164 47908 52782
rect 48860 52388 48916 52894
rect 49980 52948 50036 52958
rect 49196 52836 49252 52846
rect 49532 52836 49588 52846
rect 49196 52834 49588 52836
rect 49196 52782 49198 52834
rect 49250 52782 49534 52834
rect 49586 52782 49588 52834
rect 49196 52780 49588 52782
rect 49196 52770 49252 52780
rect 49532 52770 49588 52780
rect 49868 52834 49924 52846
rect 49868 52782 49870 52834
rect 49922 52782 49924 52834
rect 48916 52332 49028 52388
rect 48860 52322 48916 52332
rect 47404 52162 47908 52164
rect 47404 52110 47406 52162
rect 47458 52110 47854 52162
rect 47906 52110 47908 52162
rect 47404 52108 47908 52110
rect 47404 52098 47460 52108
rect 47852 52098 47908 52108
rect 47068 51940 47124 51950
rect 47068 51846 47124 51884
rect 47740 51940 47796 51950
rect 47740 51938 48132 51940
rect 47740 51886 47742 51938
rect 47794 51886 48132 51938
rect 47740 51884 48132 51886
rect 47740 51874 47796 51884
rect 47628 51492 47684 51502
rect 48076 51492 48132 51884
rect 47628 51490 47796 51492
rect 47628 51438 47630 51490
rect 47682 51438 47796 51490
rect 47628 51436 47796 51438
rect 47628 51426 47684 51436
rect 46956 50484 47012 51324
rect 47068 51378 47124 51390
rect 47068 51326 47070 51378
rect 47122 51326 47124 51378
rect 47068 51044 47124 51326
rect 47516 51378 47572 51390
rect 47516 51326 47518 51378
rect 47570 51326 47572 51378
rect 47516 51156 47572 51326
rect 47516 51090 47572 51100
rect 47628 51154 47684 51166
rect 47628 51102 47630 51154
rect 47682 51102 47684 51154
rect 47068 50978 47124 50988
rect 47068 50708 47124 50718
rect 47068 50614 47124 50652
rect 47516 50596 47572 50606
rect 47292 50484 47348 50522
rect 47516 50502 47572 50540
rect 46956 50428 47124 50484
rect 47068 50372 47236 50428
rect 47292 50418 47348 50428
rect 47180 49588 47236 50372
rect 47628 49924 47684 51102
rect 47740 50932 47796 51436
rect 47740 50866 47796 50876
rect 47964 51156 48020 51166
rect 47628 49858 47684 49868
rect 47740 50484 47796 50494
rect 47628 49698 47684 49710
rect 47628 49646 47630 49698
rect 47682 49646 47684 49698
rect 47628 49588 47684 49646
rect 47180 49532 47684 49588
rect 46844 49186 46900 49196
rect 47628 49026 47684 49532
rect 47628 48974 47630 49026
rect 47682 48974 47684 49026
rect 47628 48962 47684 48974
rect 46956 48916 47012 48926
rect 46620 48914 47012 48916
rect 46620 48862 46958 48914
rect 47010 48862 47012 48914
rect 46620 48860 47012 48862
rect 45388 48190 45390 48242
rect 45442 48190 45444 48242
rect 45388 48132 45444 48190
rect 45388 48066 45444 48076
rect 46060 48356 46116 48366
rect 45164 47630 45166 47682
rect 45218 47630 45220 47682
rect 45164 47618 45220 47630
rect 44716 46674 44772 47516
rect 45388 47572 45444 47582
rect 44940 47458 44996 47470
rect 44940 47406 44942 47458
rect 44994 47406 44996 47458
rect 44828 47348 44884 47358
rect 44828 47254 44884 47292
rect 44716 46622 44718 46674
rect 44770 46622 44772 46674
rect 44716 46610 44772 46622
rect 44940 46676 44996 47406
rect 45388 47460 45444 47516
rect 45836 47572 45892 47582
rect 45388 47458 45668 47460
rect 45388 47406 45390 47458
rect 45442 47406 45668 47458
rect 45388 47404 45668 47406
rect 45388 47394 45444 47404
rect 44940 46610 44996 46620
rect 41692 46564 41748 46574
rect 41692 46470 41748 46508
rect 43820 46562 43876 46574
rect 43820 46510 43822 46562
rect 43874 46510 43876 46562
rect 43820 46114 43876 46510
rect 45052 46450 45108 46462
rect 45052 46398 45054 46450
rect 45106 46398 45108 46450
rect 45052 46228 45108 46398
rect 45052 46162 45108 46172
rect 43820 46062 43822 46114
rect 43874 46062 43876 46114
rect 43820 46050 43876 46062
rect 44380 46114 44436 46126
rect 44380 46062 44382 46114
rect 44434 46062 44436 46114
rect 40908 45838 40910 45890
rect 40962 45838 40964 45890
rect 39676 45330 39844 45332
rect 39676 45278 39678 45330
rect 39730 45278 39844 45330
rect 39676 45276 39844 45278
rect 40348 45332 40404 45342
rect 39676 45266 39732 45276
rect 38332 45054 38334 45106
rect 38386 45054 38388 45106
rect 38332 45042 38388 45054
rect 38556 45218 38612 45230
rect 39564 45220 39620 45230
rect 40236 45220 40292 45230
rect 38556 45166 38558 45218
rect 38610 45166 38612 45218
rect 37772 44382 37774 44434
rect 37826 44382 37828 44434
rect 36092 44324 36148 44334
rect 36092 42868 36148 44268
rect 36988 43652 37044 43662
rect 36092 42866 36708 42868
rect 36092 42814 36094 42866
rect 36146 42814 36708 42866
rect 36092 42812 36708 42814
rect 36092 42802 36148 42812
rect 36204 42196 36260 42206
rect 36092 42082 36148 42094
rect 36092 42030 36094 42082
rect 36146 42030 36148 42082
rect 36092 41188 36148 42030
rect 36204 41858 36260 42140
rect 36204 41806 36206 41858
rect 36258 41806 36260 41858
rect 36204 41794 36260 41806
rect 36652 42194 36708 42812
rect 36988 42756 37044 43596
rect 37772 43652 37828 44382
rect 37772 43586 37828 43596
rect 37996 44324 38052 44334
rect 37996 43426 38052 44268
rect 38444 44212 38500 44222
rect 38444 44118 38500 44156
rect 38556 43876 38612 45166
rect 39340 45164 39564 45220
rect 39340 44434 39396 45164
rect 39564 45126 39620 45164
rect 39900 45218 40292 45220
rect 39900 45166 40238 45218
rect 40290 45166 40292 45218
rect 39900 45164 40292 45166
rect 39676 44884 39732 44894
rect 39676 44790 39732 44828
rect 39340 44382 39342 44434
rect 39394 44382 39396 44434
rect 39340 44370 39396 44382
rect 38780 44324 38836 44334
rect 38780 44230 38836 44268
rect 39788 44324 39844 44334
rect 39788 44230 39844 44268
rect 39116 44212 39172 44222
rect 38668 43876 38724 43886
rect 38556 43820 38668 43876
rect 38556 43650 38612 43662
rect 38556 43598 38558 43650
rect 38610 43598 38612 43650
rect 38444 43540 38500 43550
rect 38444 43446 38500 43484
rect 37996 43374 37998 43426
rect 38050 43374 38052 43426
rect 37996 43362 38052 43374
rect 38556 43316 38612 43598
rect 38556 43250 38612 43260
rect 36988 42754 37156 42756
rect 36988 42702 36990 42754
rect 37042 42702 37156 42754
rect 36988 42700 37156 42702
rect 36988 42690 37044 42700
rect 36652 42142 36654 42194
rect 36706 42142 36708 42194
rect 36204 41300 36260 41310
rect 36204 41206 36260 41244
rect 36092 41122 36148 41132
rect 36652 41076 36708 42142
rect 37100 42194 37156 42700
rect 37100 42142 37102 42194
rect 37154 42142 37156 42194
rect 36988 42084 37044 42094
rect 36988 41186 37044 42028
rect 37100 41300 37156 42142
rect 37772 42642 37828 42654
rect 37772 42590 37774 42642
rect 37826 42590 37828 42642
rect 37772 42196 37828 42590
rect 37772 42130 37828 42140
rect 38668 41970 38724 43820
rect 39116 43652 39172 44156
rect 39004 43650 39172 43652
rect 39004 43598 39118 43650
rect 39170 43598 39172 43650
rect 39004 43596 39172 43598
rect 38780 43538 38836 43550
rect 38780 43486 38782 43538
rect 38834 43486 38836 43538
rect 38780 42756 38836 43486
rect 38892 43540 38948 43550
rect 38892 43446 38948 43484
rect 38780 42690 38836 42700
rect 39004 42868 39060 43596
rect 39116 43586 39172 43596
rect 39228 44100 39284 44110
rect 39228 43650 39284 44044
rect 39900 43876 39956 45164
rect 40236 45154 40292 45164
rect 40348 45218 40404 45276
rect 40348 45166 40350 45218
rect 40402 45166 40404 45218
rect 40348 45154 40404 45166
rect 40796 44994 40852 45006
rect 40796 44942 40798 44994
rect 40850 44942 40852 44994
rect 40236 44882 40292 44894
rect 40236 44830 40238 44882
rect 40290 44830 40292 44882
rect 40124 44434 40180 44446
rect 40124 44382 40126 44434
rect 40178 44382 40180 44434
rect 40124 44100 40180 44382
rect 40124 44034 40180 44044
rect 39228 43598 39230 43650
rect 39282 43598 39284 43650
rect 39228 43586 39284 43598
rect 39564 43764 39620 43774
rect 39564 43650 39620 43708
rect 39788 43764 39844 43774
rect 39900 43764 39956 43820
rect 39788 43762 39956 43764
rect 39788 43710 39790 43762
rect 39842 43710 39956 43762
rect 39788 43708 39956 43710
rect 39788 43698 39844 43708
rect 39564 43598 39566 43650
rect 39618 43598 39620 43650
rect 39564 43586 39620 43598
rect 39900 43428 39956 43438
rect 39900 43334 39956 43372
rect 40236 43316 40292 44830
rect 40796 44436 40852 44942
rect 40684 44434 40852 44436
rect 40684 44382 40798 44434
rect 40850 44382 40852 44434
rect 40684 44380 40852 44382
rect 40348 43652 40404 43662
rect 40348 43558 40404 43596
rect 40236 43250 40292 43260
rect 38668 41918 38670 41970
rect 38722 41918 38724 41970
rect 38668 41906 38724 41918
rect 38892 41972 38948 41982
rect 39004 41972 39060 42812
rect 39900 42866 39956 42878
rect 39900 42814 39902 42866
rect 39954 42814 39956 42866
rect 39900 42644 39956 42814
rect 40348 42756 40404 42766
rect 40348 42662 40404 42700
rect 39900 42578 39956 42588
rect 40124 42532 40180 42542
rect 40124 42084 40180 42476
rect 38892 41970 39060 41972
rect 38892 41918 38894 41970
rect 38946 41918 39060 41970
rect 38892 41916 39060 41918
rect 39788 41972 39844 41982
rect 39788 41970 39956 41972
rect 39788 41918 39790 41970
rect 39842 41918 39956 41970
rect 39788 41916 39956 41918
rect 38892 41906 38948 41916
rect 39788 41906 39844 41916
rect 38332 41860 38388 41870
rect 38332 41412 38388 41804
rect 39900 41860 39956 41916
rect 40124 41970 40180 42028
rect 40124 41918 40126 41970
rect 40178 41918 40180 41970
rect 40124 41906 40180 41918
rect 39900 41794 39956 41804
rect 38332 41346 38388 41356
rect 39116 41746 39172 41758
rect 39116 41694 39118 41746
rect 39170 41694 39172 41746
rect 37156 41244 37380 41300
rect 37100 41234 37156 41244
rect 36988 41134 36990 41186
rect 37042 41134 37044 41186
rect 36988 41122 37044 41134
rect 36652 41010 36708 41020
rect 37212 41076 37268 41086
rect 37212 40982 37268 41020
rect 37100 40962 37156 40974
rect 37100 40910 37102 40962
rect 37154 40910 37156 40962
rect 37100 40740 37156 40910
rect 37100 40674 37156 40684
rect 37324 40404 37380 41244
rect 37100 40348 37324 40404
rect 35980 39218 36036 39228
rect 36428 39732 36484 39742
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34636 38276 34692 38286
rect 34636 38162 34692 38220
rect 34636 38110 34638 38162
rect 34690 38110 34692 38162
rect 33964 36484 34020 36494
rect 33964 36370 34020 36428
rect 33964 36318 33966 36370
rect 34018 36318 34020 36370
rect 33964 36306 34020 36318
rect 33740 35812 33796 35822
rect 33796 35756 33908 35812
rect 33740 35718 33796 35756
rect 33852 35364 33908 35756
rect 34076 35700 34132 35710
rect 34076 35698 34244 35700
rect 34076 35646 34078 35698
rect 34130 35646 34244 35698
rect 34076 35644 34244 35646
rect 34076 35634 34132 35644
rect 33852 34692 33908 35308
rect 33628 33954 33684 33964
rect 33740 34690 33908 34692
rect 33740 34638 33854 34690
rect 33906 34638 33908 34690
rect 33740 34636 33908 34638
rect 33516 33628 33684 33684
rect 33068 33236 33124 33246
rect 31948 33234 33124 33236
rect 31948 33182 33070 33234
rect 33122 33182 33124 33234
rect 31948 33180 33124 33182
rect 31948 32786 32004 33180
rect 31948 32734 31950 32786
rect 32002 32734 32004 32786
rect 31948 32722 32004 32734
rect 31276 32510 31278 32562
rect 31330 32510 31332 32562
rect 30828 32498 30884 32508
rect 30044 31666 30100 31948
rect 30380 31780 30436 31790
rect 30940 31780 30996 32508
rect 31276 32452 31332 32510
rect 31052 32396 31332 32452
rect 32396 32676 32452 32686
rect 32396 32450 32452 32620
rect 32396 32398 32398 32450
rect 32450 32398 32452 32450
rect 31052 31892 31108 32396
rect 32396 32386 32452 32398
rect 31052 31826 31108 31836
rect 30380 31778 30996 31780
rect 30380 31726 30382 31778
rect 30434 31726 30996 31778
rect 30380 31724 30996 31726
rect 30380 31714 30436 31724
rect 30044 31614 30046 31666
rect 30098 31614 30100 31666
rect 30044 31602 30100 31614
rect 30940 31668 30996 31724
rect 32172 31778 32228 31790
rect 32172 31726 32174 31778
rect 32226 31726 32228 31778
rect 31612 31668 31668 31678
rect 30940 31666 31668 31668
rect 30940 31614 31614 31666
rect 31666 31614 31668 31666
rect 30940 31612 31668 31614
rect 31612 31602 31668 31612
rect 29708 31126 29764 31164
rect 31052 31220 31108 31230
rect 30156 31106 30212 31118
rect 30156 31054 30158 31106
rect 30210 31054 30212 31106
rect 29708 30996 29764 31006
rect 30044 30996 30100 31006
rect 29764 30994 30100 30996
rect 29764 30942 30046 30994
rect 30098 30942 30100 30994
rect 29764 30940 30100 30942
rect 30156 30996 30212 31054
rect 30156 30940 30772 30996
rect 29708 30930 29764 30940
rect 30044 30930 30100 30940
rect 30716 30882 30772 30940
rect 30716 30830 30718 30882
rect 30770 30830 30772 30882
rect 30156 30772 30212 30782
rect 30156 30678 30212 30716
rect 30604 30770 30660 30782
rect 30604 30718 30606 30770
rect 30658 30718 30660 30770
rect 29596 30210 30100 30212
rect 29596 30158 29598 30210
rect 29650 30158 30100 30210
rect 29596 30156 30100 30158
rect 29596 30146 29652 30156
rect 29372 30100 29428 30110
rect 29260 29988 29316 29998
rect 28812 29986 29316 29988
rect 28812 29934 29262 29986
rect 29314 29934 29316 29986
rect 28812 29932 29316 29934
rect 28812 29538 28868 29932
rect 29260 29922 29316 29932
rect 28812 29486 28814 29538
rect 28866 29486 28868 29538
rect 28812 29474 28868 29486
rect 28252 28774 28308 28812
rect 28476 28924 28644 28980
rect 27916 28590 27918 28642
rect 27970 28590 27972 28642
rect 27916 28578 27972 28590
rect 28476 28530 28532 28924
rect 29148 28868 29204 28878
rect 29148 28774 29204 28812
rect 28588 28756 28644 28766
rect 28588 28754 28756 28756
rect 28588 28702 28590 28754
rect 28642 28702 28756 28754
rect 28588 28700 28756 28702
rect 28588 28690 28644 28700
rect 28476 28478 28478 28530
rect 28530 28478 28532 28530
rect 28476 28466 28532 28478
rect 28364 27858 28420 27870
rect 28364 27806 28366 27858
rect 28418 27806 28420 27858
rect 28364 27748 28420 27806
rect 28420 27692 28532 27748
rect 28364 27682 28420 27692
rect 28476 27186 28532 27692
rect 28476 27134 28478 27186
rect 28530 27134 28532 27186
rect 28476 26908 28532 27134
rect 28476 26852 28644 26908
rect 27804 25566 27806 25618
rect 27858 25566 27860 25618
rect 27804 25554 27860 25566
rect 28476 26292 28532 26302
rect 28476 24946 28532 26236
rect 28476 24894 28478 24946
rect 28530 24894 28532 24946
rect 28476 24882 28532 24894
rect 28588 25506 28644 26852
rect 28700 26292 28756 28700
rect 29372 28644 29428 30044
rect 30044 28754 30100 30156
rect 30604 30100 30660 30718
rect 30604 30034 30660 30044
rect 30716 29316 30772 30830
rect 31052 30210 31108 31164
rect 32172 30772 32228 31726
rect 32508 31780 32564 31790
rect 32508 31666 32564 31724
rect 32732 31778 32788 33180
rect 33068 33170 33124 33180
rect 33180 32676 33236 33404
rect 33516 33458 33572 33470
rect 33516 33406 33518 33458
rect 33570 33406 33572 33458
rect 32732 31726 32734 31778
rect 32786 31726 32788 31778
rect 32732 31714 32788 31726
rect 33068 32620 33236 32676
rect 33292 32676 33348 32686
rect 33068 31892 33124 32620
rect 33180 32452 33236 32462
rect 33292 32452 33348 32620
rect 33180 32450 33460 32452
rect 33180 32398 33182 32450
rect 33234 32398 33460 32450
rect 33180 32396 33460 32398
rect 33180 32386 33236 32396
rect 33404 32116 33460 32396
rect 33516 32340 33572 33406
rect 33628 32676 33684 33628
rect 33740 33460 33796 34636
rect 33852 34626 33908 34636
rect 33964 34690 34020 34702
rect 33964 34638 33966 34690
rect 34018 34638 34020 34690
rect 33964 34132 34020 34638
rect 34076 34692 34132 34702
rect 34076 34598 34132 34636
rect 33964 34066 34020 34076
rect 34188 34132 34244 35644
rect 34300 35476 34356 36540
rect 34300 35410 34356 35420
rect 34412 37604 34468 37614
rect 34412 35026 34468 37548
rect 34636 37044 34692 38110
rect 35084 37828 35140 37838
rect 35084 37268 35140 37772
rect 36204 37828 36260 37838
rect 36428 37828 36484 39676
rect 37100 39732 37156 40348
rect 37324 40338 37380 40348
rect 37548 41186 37604 41198
rect 37548 41134 37550 41186
rect 37602 41134 37604 41186
rect 37548 40964 37604 41134
rect 39116 41076 39172 41694
rect 39116 41010 39172 41020
rect 39340 41746 39396 41758
rect 39340 41694 39342 41746
rect 39394 41694 39396 41746
rect 39340 41636 39396 41694
rect 39452 41748 39508 41758
rect 39788 41748 39844 41758
rect 39452 41746 39620 41748
rect 39452 41694 39454 41746
rect 39506 41694 39620 41746
rect 39452 41692 39620 41694
rect 39452 41682 39508 41692
rect 38108 40964 38164 40974
rect 37548 40908 38108 40964
rect 37100 39618 37156 39676
rect 37100 39566 37102 39618
rect 37154 39566 37156 39618
rect 37100 39554 37156 39566
rect 37548 39172 37604 40908
rect 38108 40870 38164 40908
rect 38892 40964 38948 40974
rect 38892 40870 38948 40908
rect 39228 40962 39284 40974
rect 39228 40910 39230 40962
rect 39282 40910 39284 40962
rect 37884 40740 37940 40750
rect 37940 40684 38276 40740
rect 37884 40674 37940 40684
rect 38220 40514 38276 40684
rect 38444 40628 38500 40638
rect 38444 40534 38500 40572
rect 38220 40462 38222 40514
rect 38274 40462 38276 40514
rect 38220 40450 38276 40462
rect 39004 40404 39060 40414
rect 39004 40310 39060 40348
rect 39228 40404 39284 40910
rect 39340 40964 39396 41580
rect 39564 41186 39620 41692
rect 39564 41134 39566 41186
rect 39618 41134 39620 41186
rect 39564 41122 39620 41134
rect 39676 41746 39844 41748
rect 39676 41694 39790 41746
rect 39842 41694 39844 41746
rect 39676 41692 39844 41694
rect 39676 41074 39732 41692
rect 39788 41682 39844 41692
rect 39676 41022 39678 41074
rect 39730 41022 39732 41074
rect 39676 41010 39732 41022
rect 39788 41076 39844 41086
rect 39340 40898 39396 40908
rect 39788 40516 39844 41020
rect 39788 40422 39844 40460
rect 39900 40962 39956 40974
rect 39900 40910 39902 40962
rect 39954 40910 39956 40962
rect 39228 40338 39284 40348
rect 37884 40292 37940 40302
rect 37884 40198 37940 40236
rect 38332 40290 38388 40302
rect 38332 40238 38334 40290
rect 38386 40238 38388 40290
rect 38332 39956 38388 40238
rect 37772 39900 38388 39956
rect 39900 39956 39956 40910
rect 37772 39730 37828 39900
rect 39900 39890 39956 39900
rect 40012 40402 40068 40414
rect 40012 40350 40014 40402
rect 40066 40350 40068 40402
rect 37772 39678 37774 39730
rect 37826 39678 37828 39730
rect 37772 39666 37828 39678
rect 38892 39844 38948 39854
rect 37436 38946 37492 38958
rect 37436 38894 37438 38946
rect 37490 38894 37492 38946
rect 37324 38834 37380 38846
rect 37324 38782 37326 38834
rect 37378 38782 37380 38834
rect 37324 38668 37380 38782
rect 36876 38612 37380 38668
rect 36764 38388 36820 38398
rect 36652 38332 36764 38388
rect 36260 37772 36484 37828
rect 36540 37940 36596 37950
rect 36204 37734 36260 37772
rect 35084 37202 35140 37212
rect 35868 37604 35924 37614
rect 34636 35138 34692 36988
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35868 36370 35924 37548
rect 36428 37604 36484 37614
rect 36428 37490 36484 37548
rect 36428 37438 36430 37490
rect 36482 37438 36484 37490
rect 36428 37426 36484 37438
rect 36204 37380 36260 37390
rect 36204 37286 36260 37324
rect 36540 37266 36596 37884
rect 36540 37214 36542 37266
rect 36594 37214 36596 37266
rect 35980 37154 36036 37166
rect 35980 37102 35982 37154
rect 36034 37102 36036 37154
rect 35980 36484 36036 37102
rect 36540 36708 36596 37214
rect 36540 36642 36596 36652
rect 36652 37156 36708 38332
rect 36764 38322 36820 38332
rect 36876 37380 36932 38612
rect 37436 38388 37492 38894
rect 37548 38668 37604 39116
rect 37884 39116 38388 39172
rect 37660 39060 37716 39070
rect 37884 39060 37940 39116
rect 37660 39058 37940 39060
rect 37660 39006 37662 39058
rect 37714 39006 37940 39058
rect 37660 39004 37940 39006
rect 37660 38994 37716 39004
rect 37996 38946 38052 38958
rect 37996 38894 37998 38946
rect 38050 38894 38052 38946
rect 37884 38834 37940 38846
rect 37884 38782 37886 38834
rect 37938 38782 37940 38834
rect 37548 38612 37828 38668
rect 36988 38332 37492 38388
rect 36988 37492 37044 38332
rect 37212 38052 37268 38062
rect 37772 38052 37828 38612
rect 37884 38388 37940 38782
rect 37996 38668 38052 38894
rect 38220 38836 38276 38846
rect 38220 38742 38276 38780
rect 37996 38612 38276 38668
rect 38108 38388 38164 38398
rect 37884 38322 37940 38332
rect 37996 38332 38108 38388
rect 37772 37996 37940 38052
rect 37212 37958 37268 37996
rect 37324 37940 37380 37950
rect 37324 37846 37380 37884
rect 37100 37826 37156 37838
rect 37772 37828 37828 37838
rect 37100 37774 37102 37826
rect 37154 37774 37156 37826
rect 37100 37716 37156 37774
rect 37100 37650 37156 37660
rect 37548 37826 37828 37828
rect 37548 37774 37774 37826
rect 37826 37774 37828 37826
rect 37548 37772 37828 37774
rect 36988 37436 37156 37492
rect 36876 37314 36932 37324
rect 37100 37378 37156 37436
rect 37100 37326 37102 37378
rect 37154 37326 37156 37378
rect 36988 37266 37044 37278
rect 36988 37214 36990 37266
rect 37042 37214 37044 37266
rect 36988 37156 37044 37214
rect 36652 37100 37044 37156
rect 36092 36484 36148 36494
rect 35980 36428 36092 36484
rect 36092 36390 36148 36428
rect 35868 36318 35870 36370
rect 35922 36318 35924 36370
rect 35868 36306 35924 36318
rect 35756 36148 35812 36158
rect 34972 35364 35028 35374
rect 35028 35308 35140 35364
rect 34972 35298 35028 35308
rect 34636 35086 34638 35138
rect 34690 35086 34692 35138
rect 34636 35074 34692 35086
rect 35084 35138 35140 35308
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35084 35086 35086 35138
rect 35138 35086 35140 35138
rect 35084 35074 35140 35086
rect 34412 34974 34414 35026
rect 34466 34974 34468 35026
rect 34412 34962 34468 34974
rect 34860 35028 34916 35038
rect 34860 34934 34916 34972
rect 35756 34804 35812 36092
rect 36652 35812 36708 37100
rect 37100 37044 37156 37326
rect 37212 37380 37268 37390
rect 37548 37380 37604 37772
rect 37772 37762 37828 37772
rect 37268 37324 37604 37380
rect 37660 37380 37716 37390
rect 37212 37286 37268 37324
rect 37660 37286 37716 37324
rect 37100 36988 37604 37044
rect 37324 36820 37380 36830
rect 37212 36708 37268 36718
rect 37212 36614 37268 36652
rect 36988 36484 37044 36494
rect 36988 36390 37044 36428
rect 36652 35718 36708 35756
rect 37324 35698 37380 36764
rect 37548 36706 37604 36988
rect 37548 36654 37550 36706
rect 37602 36654 37604 36706
rect 37548 36642 37604 36654
rect 37324 35646 37326 35698
rect 37378 35646 37380 35698
rect 37324 35634 37380 35646
rect 37548 35700 37604 35710
rect 37548 35606 37604 35644
rect 37884 35252 37940 37996
rect 37996 38050 38052 38332
rect 38108 38322 38164 38332
rect 38220 38276 38276 38612
rect 38220 38210 38276 38220
rect 37996 37998 37998 38050
rect 38050 37998 38052 38050
rect 37996 37986 38052 37998
rect 38108 38164 38164 38174
rect 38108 38050 38164 38108
rect 38108 37998 38110 38050
rect 38162 37998 38164 38050
rect 38108 37986 38164 37998
rect 38220 38052 38276 38090
rect 38220 37986 38276 37996
rect 38220 37604 38276 37614
rect 37996 37380 38052 37390
rect 37996 37286 38052 37324
rect 38220 37266 38276 37548
rect 38220 37214 38222 37266
rect 38274 37214 38276 37266
rect 38220 35698 38276 37214
rect 38332 36482 38388 39116
rect 38556 38948 38612 38958
rect 38444 38946 38612 38948
rect 38444 38894 38558 38946
rect 38610 38894 38612 38946
rect 38444 38892 38612 38894
rect 38444 38388 38500 38892
rect 38556 38882 38612 38892
rect 38668 38836 38724 38846
rect 38668 38742 38724 38780
rect 38444 38050 38500 38332
rect 38444 37998 38446 38050
rect 38498 37998 38500 38050
rect 38444 37986 38500 37998
rect 38556 38610 38612 38622
rect 38556 38558 38558 38610
rect 38610 38558 38612 38610
rect 38556 36594 38612 38558
rect 38780 37938 38836 37950
rect 38780 37886 38782 37938
rect 38834 37886 38836 37938
rect 38668 37826 38724 37838
rect 38668 37774 38670 37826
rect 38722 37774 38724 37826
rect 38668 37156 38724 37774
rect 38668 37090 38724 37100
rect 38556 36542 38558 36594
rect 38610 36542 38612 36594
rect 38556 36530 38612 36542
rect 38332 36430 38334 36482
rect 38386 36430 38388 36482
rect 38332 36418 38388 36430
rect 38220 35646 38222 35698
rect 38274 35646 38276 35698
rect 37884 35196 38052 35252
rect 34188 34066 34244 34076
rect 34300 34692 34356 34702
rect 33852 34018 33908 34030
rect 33852 33966 33854 34018
rect 33906 33966 33908 34018
rect 33852 33684 33908 33966
rect 34300 33684 34356 34636
rect 35532 34690 35588 34702
rect 35532 34638 35534 34690
rect 35586 34638 35588 34690
rect 33852 33628 34132 33684
rect 33740 33404 34020 33460
rect 33740 32676 33796 32686
rect 33628 32674 33796 32676
rect 33628 32622 33742 32674
rect 33794 32622 33796 32674
rect 33628 32620 33796 32622
rect 33740 32610 33796 32620
rect 33964 32562 34020 33404
rect 34076 32786 34132 33628
rect 34076 32734 34078 32786
rect 34130 32734 34132 32786
rect 34076 32722 34132 32734
rect 34300 32674 34356 33628
rect 34300 32622 34302 32674
rect 34354 32622 34356 32674
rect 34300 32610 34356 32622
rect 34412 34020 34468 34030
rect 33964 32510 33966 32562
rect 34018 32510 34020 32562
rect 33964 32498 34020 32510
rect 33516 32274 33572 32284
rect 33404 32060 33684 32116
rect 32508 31614 32510 31666
rect 32562 31614 32564 31666
rect 32508 31602 32564 31614
rect 33068 30996 33124 31836
rect 33628 31890 33684 32060
rect 33628 31838 33630 31890
rect 33682 31838 33684 31890
rect 33180 31668 33236 31678
rect 33180 31666 33348 31668
rect 33180 31614 33182 31666
rect 33234 31614 33348 31666
rect 33180 31612 33348 31614
rect 33180 31602 33236 31612
rect 33068 30994 33236 30996
rect 33068 30942 33070 30994
rect 33122 30942 33236 30994
rect 33068 30940 33236 30942
rect 33068 30930 33124 30940
rect 32172 30706 32228 30716
rect 32172 30548 32228 30558
rect 31052 30158 31054 30210
rect 31106 30158 31108 30210
rect 31052 30146 31108 30158
rect 31948 30492 32172 30548
rect 31948 29650 32004 30492
rect 32172 30482 32228 30492
rect 31948 29598 31950 29650
rect 32002 29598 32004 29650
rect 31948 29586 32004 29598
rect 32284 29428 32340 29438
rect 32284 29334 32340 29372
rect 33068 29428 33124 29438
rect 30940 29316 30996 29326
rect 30716 29314 30996 29316
rect 30716 29262 30942 29314
rect 30994 29262 30996 29314
rect 30716 29260 30996 29262
rect 30940 29250 30996 29260
rect 32508 29316 32564 29326
rect 32508 29222 32564 29260
rect 33068 28980 33124 29372
rect 33068 28914 33124 28924
rect 30044 28702 30046 28754
rect 30098 28702 30100 28754
rect 30044 28690 30100 28702
rect 32172 28754 32228 28766
rect 33180 28756 33236 30940
rect 33292 29988 33348 31612
rect 33404 31666 33460 31678
rect 33404 31614 33406 31666
rect 33458 31614 33460 31666
rect 33404 30548 33460 31614
rect 33628 30548 33684 31838
rect 33852 31780 33908 31790
rect 33740 31778 33908 31780
rect 33740 31726 33854 31778
rect 33906 31726 33908 31778
rect 33740 31724 33908 31726
rect 33740 31556 33796 31724
rect 33852 31714 33908 31724
rect 34076 31666 34132 31678
rect 34076 31614 34078 31666
rect 34130 31614 34132 31666
rect 33964 31556 34020 31566
rect 33740 31490 33796 31500
rect 33852 31554 34020 31556
rect 33852 31502 33966 31554
rect 34018 31502 34020 31554
rect 33852 31500 34020 31502
rect 33852 31106 33908 31500
rect 33964 31490 34020 31500
rect 33852 31054 33854 31106
rect 33906 31054 33908 31106
rect 33852 31042 33908 31054
rect 33628 30492 33908 30548
rect 33404 30482 33460 30492
rect 33292 29932 33460 29988
rect 32172 28702 32174 28754
rect 32226 28702 32228 28754
rect 29484 28644 29540 28654
rect 29372 28642 29540 28644
rect 29372 28590 29486 28642
rect 29538 28590 29540 28642
rect 29372 28588 29540 28590
rect 29484 28578 29540 28588
rect 29260 28418 29316 28430
rect 29260 28366 29262 28418
rect 29314 28366 29316 28418
rect 28812 27858 28868 27870
rect 28812 27806 28814 27858
rect 28866 27806 28868 27858
rect 28812 27748 28868 27806
rect 28812 27682 28868 27692
rect 29260 26908 29316 28366
rect 31836 28082 31892 28094
rect 31836 28030 31838 28082
rect 31890 28030 31892 28082
rect 31836 27972 31892 28030
rect 31500 27916 31836 27972
rect 29596 27746 29652 27758
rect 29596 27694 29598 27746
rect 29650 27694 29652 27746
rect 29260 26852 29540 26908
rect 29036 26404 29092 26414
rect 29036 26402 29204 26404
rect 29036 26350 29038 26402
rect 29090 26350 29204 26402
rect 29036 26348 29204 26350
rect 29036 26338 29092 26348
rect 28700 26198 28756 26236
rect 28588 25454 28590 25506
rect 28642 25454 28644 25506
rect 28588 25396 28644 25454
rect 28140 24836 28196 24846
rect 28140 24834 28420 24836
rect 28140 24782 28142 24834
rect 28194 24782 28420 24834
rect 28140 24780 28420 24782
rect 28140 24770 28196 24780
rect 27804 23044 27860 23054
rect 27244 23042 27860 23044
rect 27244 22990 27806 23042
rect 27858 22990 27860 23042
rect 27244 22988 27860 22990
rect 27020 22260 27076 22270
rect 27020 22166 27076 22204
rect 26908 22082 26964 22092
rect 27132 21812 27188 21822
rect 27244 21812 27300 22988
rect 27804 22978 27860 22988
rect 27692 22372 27748 22382
rect 27692 22278 27748 22316
rect 28252 22258 28308 22270
rect 28252 22206 28254 22258
rect 28306 22206 28308 22258
rect 27132 21810 27300 21812
rect 27132 21758 27134 21810
rect 27186 21758 27300 21810
rect 27132 21756 27300 21758
rect 27356 22146 27412 22158
rect 27356 22094 27358 22146
rect 27410 22094 27412 22146
rect 27132 21746 27188 21756
rect 26908 21586 26964 21598
rect 26908 21534 26910 21586
rect 26962 21534 26964 21586
rect 26908 21476 26964 21534
rect 27356 21476 27412 22094
rect 27580 22148 27636 22158
rect 26908 21420 27412 21476
rect 27468 21700 27524 21710
rect 26348 21196 26852 21252
rect 26348 20914 26404 21196
rect 26348 20862 26350 20914
rect 26402 20862 26404 20914
rect 26348 20850 26404 20862
rect 27468 20914 27524 21644
rect 27468 20862 27470 20914
rect 27522 20862 27524 20914
rect 27468 20850 27524 20862
rect 27020 20690 27076 20702
rect 27020 20638 27022 20690
rect 27074 20638 27076 20690
rect 26684 20580 26740 20590
rect 26236 20178 26292 20188
rect 26460 20578 26740 20580
rect 26460 20526 26686 20578
rect 26738 20526 26740 20578
rect 26460 20524 26740 20526
rect 26124 20066 26180 20076
rect 26348 20132 26404 20142
rect 26460 20132 26516 20524
rect 26684 20514 26740 20524
rect 26348 20130 26516 20132
rect 26348 20078 26350 20130
rect 26402 20078 26516 20130
rect 26348 20076 26516 20078
rect 27020 20132 27076 20638
rect 27132 20356 27188 20366
rect 27188 20300 27300 20356
rect 27132 20290 27188 20300
rect 26348 20066 26404 20076
rect 27020 20066 27076 20076
rect 25900 18050 25956 18060
rect 26012 19234 26068 19246
rect 26012 19182 26014 19234
rect 26066 19182 26068 19234
rect 25788 17838 25790 17890
rect 25842 17838 25844 17890
rect 25788 17826 25844 17838
rect 26012 17892 26068 19182
rect 26460 19234 26516 19246
rect 26460 19182 26462 19234
rect 26514 19182 26516 19234
rect 26348 19012 26404 19022
rect 26348 18674 26404 18956
rect 26460 18900 26516 19182
rect 26460 18834 26516 18844
rect 26796 19122 26852 19134
rect 26796 19070 26798 19122
rect 26850 19070 26852 19122
rect 26348 18622 26350 18674
rect 26402 18622 26404 18674
rect 26348 18610 26404 18622
rect 26012 17826 26068 17836
rect 26460 18452 26516 18462
rect 25676 17554 25732 17566
rect 25676 17502 25678 17554
rect 25730 17502 25732 17554
rect 25676 16884 25732 17502
rect 25788 17444 25844 17454
rect 25788 17442 26180 17444
rect 25788 17390 25790 17442
rect 25842 17390 26180 17442
rect 25788 17388 26180 17390
rect 25788 17378 25844 17388
rect 26012 16996 26068 17006
rect 26124 16996 26180 17388
rect 26460 17108 26516 18396
rect 26796 18338 26852 19070
rect 27020 19012 27076 19022
rect 27020 18918 27076 18956
rect 26796 18286 26798 18338
rect 26850 18286 26852 18338
rect 26796 18116 26852 18286
rect 27244 18562 27300 20300
rect 27580 19348 27636 22092
rect 28252 20356 28308 22206
rect 28364 21812 28420 24780
rect 28588 23154 28644 25340
rect 28588 23102 28590 23154
rect 28642 23102 28644 23154
rect 28588 23044 28644 23102
rect 28588 22978 28644 22988
rect 28924 25060 28980 25070
rect 28924 24610 28980 25004
rect 28924 24558 28926 24610
rect 28978 24558 28980 24610
rect 28476 22370 28532 22382
rect 28476 22318 28478 22370
rect 28530 22318 28532 22370
rect 28476 22260 28532 22318
rect 28476 22194 28532 22204
rect 28364 21756 28644 21812
rect 28588 21252 28644 21756
rect 28588 20916 28644 21196
rect 28588 20822 28644 20860
rect 28700 21364 28756 21374
rect 28252 20290 28308 20300
rect 27580 19282 27636 19292
rect 28476 19906 28532 19918
rect 28476 19854 28478 19906
rect 28530 19854 28532 19906
rect 28476 19796 28532 19854
rect 27804 18788 27860 18798
rect 27244 18510 27246 18562
rect 27298 18510 27300 18562
rect 27244 18228 27300 18510
rect 27692 18676 27748 18686
rect 27692 18562 27748 18620
rect 27692 18510 27694 18562
rect 27746 18510 27748 18562
rect 27692 18452 27748 18510
rect 27692 18386 27748 18396
rect 27580 18228 27636 18238
rect 27244 18162 27300 18172
rect 27468 18226 27636 18228
rect 27468 18174 27582 18226
rect 27634 18174 27636 18226
rect 27468 18172 27636 18174
rect 26796 18050 26852 18060
rect 27132 17780 27188 17790
rect 26908 17778 27188 17780
rect 26908 17726 27134 17778
rect 27186 17726 27188 17778
rect 26908 17724 27188 17726
rect 26572 17668 26628 17678
rect 26572 17574 26628 17612
rect 26908 17220 26964 17724
rect 27132 17714 27188 17724
rect 27020 17442 27076 17454
rect 27020 17390 27022 17442
rect 27074 17390 27076 17442
rect 27020 17332 27076 17390
rect 27244 17442 27300 17454
rect 27244 17390 27246 17442
rect 27298 17390 27300 17442
rect 27132 17332 27188 17342
rect 27020 17276 27132 17332
rect 27132 17266 27188 17276
rect 26460 17014 26516 17052
rect 26684 17164 26964 17220
rect 27244 17220 27300 17390
rect 26124 16940 26292 16996
rect 26012 16902 26068 16940
rect 25676 16818 25732 16828
rect 25788 16882 25844 16894
rect 25788 16830 25790 16882
rect 25842 16830 25844 16882
rect 25564 16658 25620 16670
rect 25564 16606 25566 16658
rect 25618 16606 25620 16658
rect 25564 16436 25620 16606
rect 25676 16436 25732 16446
rect 25564 16380 25676 16436
rect 25676 16370 25732 16380
rect 25452 16268 25620 16324
rect 25060 16044 25172 16100
rect 25452 16100 25508 16110
rect 25004 16034 25060 16044
rect 24556 15922 24612 15932
rect 25340 15988 25396 15998
rect 24780 15876 24836 15886
rect 24668 15820 24780 15876
rect 24220 15486 24222 15538
rect 24274 15486 24276 15538
rect 24220 15474 24276 15486
rect 24444 15540 24500 15550
rect 24668 15540 24724 15820
rect 24780 15810 24836 15820
rect 25004 15874 25060 15886
rect 25340 15876 25396 15932
rect 25004 15822 25006 15874
rect 25058 15822 25060 15874
rect 24444 15538 24724 15540
rect 24444 15486 24446 15538
rect 24498 15486 24724 15538
rect 24444 15484 24724 15486
rect 24892 15764 24948 15774
rect 24444 15474 24500 15484
rect 24556 15316 24612 15326
rect 24556 15222 24612 15260
rect 24668 15314 24724 15326
rect 24668 15262 24670 15314
rect 24722 15262 24724 15314
rect 24668 15148 24724 15262
rect 24556 15092 24724 15148
rect 24220 14642 24276 14654
rect 24220 14590 24222 14642
rect 24274 14590 24276 14642
rect 24220 14532 24276 14590
rect 24220 14466 24276 14476
rect 24108 13794 24164 13804
rect 24220 14196 24276 14206
rect 24108 13524 24164 13534
rect 23772 12562 23828 12572
rect 23884 12850 23940 12862
rect 23884 12798 23886 12850
rect 23938 12798 23940 12850
rect 23884 12404 23940 12798
rect 23884 12338 23940 12348
rect 24108 12290 24164 13468
rect 24220 12962 24276 14140
rect 24444 13636 24500 13674
rect 24444 13570 24500 13580
rect 24444 13412 24500 13422
rect 24444 13076 24500 13356
rect 24220 12910 24222 12962
rect 24274 12910 24276 12962
rect 24220 12898 24276 12910
rect 24332 12964 24388 12974
rect 24332 12870 24388 12908
rect 24444 12962 24500 13020
rect 24444 12910 24446 12962
rect 24498 12910 24500 12962
rect 24444 12898 24500 12910
rect 24556 12740 24612 15092
rect 24668 14756 24724 14766
rect 24668 14644 24724 14700
rect 24668 14642 24836 14644
rect 24668 14590 24670 14642
rect 24722 14590 24836 14642
rect 24668 14588 24836 14590
rect 24668 14578 24724 14588
rect 24668 12740 24724 12750
rect 24556 12738 24724 12740
rect 24556 12686 24670 12738
rect 24722 12686 24724 12738
rect 24556 12684 24724 12686
rect 24668 12674 24724 12684
rect 24108 12238 24110 12290
rect 24162 12238 24164 12290
rect 24108 12226 24164 12238
rect 24444 12290 24500 12302
rect 24444 12238 24446 12290
rect 24498 12238 24500 12290
rect 23772 11954 23828 11966
rect 23772 11902 23774 11954
rect 23826 11902 23828 11954
rect 23772 8484 23828 11902
rect 23996 11732 24052 11742
rect 23996 11394 24052 11676
rect 24332 11620 24388 11630
rect 24332 11506 24388 11564
rect 24332 11454 24334 11506
rect 24386 11454 24388 11506
rect 24332 11442 24388 11454
rect 23996 11342 23998 11394
rect 24050 11342 24052 11394
rect 23996 11330 24052 11342
rect 24332 10722 24388 10734
rect 24332 10670 24334 10722
rect 24386 10670 24388 10722
rect 24332 9828 24388 10670
rect 23772 8418 23828 8428
rect 23884 8930 23940 8942
rect 23884 8878 23886 8930
rect 23938 8878 23940 8930
rect 23660 8372 23716 8382
rect 23660 8260 23716 8316
rect 23660 8258 23828 8260
rect 23660 8206 23662 8258
rect 23714 8206 23828 8258
rect 23660 8204 23828 8206
rect 23660 8194 23716 8204
rect 23548 7196 23716 7252
rect 23100 6850 23156 6860
rect 23548 6916 23604 6926
rect 23548 6822 23604 6860
rect 22764 6804 22820 6814
rect 22764 6710 22820 6748
rect 23212 6692 23268 6702
rect 23660 6692 23716 7196
rect 23212 6690 23716 6692
rect 23212 6638 23214 6690
rect 23266 6638 23716 6690
rect 23212 6636 23716 6638
rect 23212 6626 23268 6636
rect 21868 5906 22148 5908
rect 21868 5854 21870 5906
rect 21922 5854 22148 5906
rect 21868 5852 22148 5854
rect 22204 6466 22260 6478
rect 22204 6414 22206 6466
rect 22258 6414 22260 6466
rect 21868 5842 21924 5852
rect 21532 5684 21588 5694
rect 20524 5682 21588 5684
rect 20524 5630 21534 5682
rect 21586 5630 21588 5682
rect 20524 5628 21588 5630
rect 19852 5236 19908 5246
rect 19628 5180 19852 5236
rect 19852 5142 19908 5180
rect 16604 5070 16606 5122
rect 16658 5070 16660 5122
rect 16604 5058 16660 5070
rect 20524 5122 20580 5628
rect 21532 5618 21588 5628
rect 21532 5348 21588 5358
rect 20524 5070 20526 5122
rect 20578 5070 20580 5122
rect 20524 5058 20580 5070
rect 20860 5236 20916 5246
rect 20748 4898 20804 4910
rect 20748 4846 20750 4898
rect 20802 4846 20804 4898
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 15484 4174 15486 4226
rect 15538 4174 15540 4226
rect 15484 4162 15540 4174
rect 20748 4116 20804 4846
rect 20860 4338 20916 5180
rect 21532 5122 21588 5292
rect 22092 5236 22148 5246
rect 22204 5236 22260 6414
rect 22652 6244 22708 6254
rect 22540 6188 22652 6244
rect 22540 6018 22596 6188
rect 22652 6178 22708 6188
rect 22540 5966 22542 6018
rect 22594 5966 22596 6018
rect 22540 5954 22596 5966
rect 22652 6020 22708 6030
rect 22652 5906 22708 5964
rect 22652 5854 22654 5906
rect 22706 5854 22708 5906
rect 22652 5842 22708 5854
rect 23548 5908 23604 5918
rect 23772 5908 23828 8204
rect 23884 8148 23940 8878
rect 24332 8820 24388 9772
rect 24332 8754 24388 8764
rect 24444 8484 24500 12238
rect 24780 12180 24836 14588
rect 24892 14532 24948 15708
rect 25004 15540 25060 15822
rect 25004 15474 25060 15484
rect 25116 15874 25396 15876
rect 25116 15822 25342 15874
rect 25394 15822 25396 15874
rect 25116 15820 25396 15822
rect 25004 14532 25060 14542
rect 24892 14530 25060 14532
rect 24892 14478 25006 14530
rect 25058 14478 25060 14530
rect 24892 14476 25060 14478
rect 25004 14466 25060 14476
rect 25116 14196 25172 15820
rect 25340 15810 25396 15820
rect 25340 15540 25396 15550
rect 25452 15540 25508 16044
rect 25340 15538 25508 15540
rect 25340 15486 25342 15538
rect 25394 15486 25508 15538
rect 25340 15484 25508 15486
rect 25564 15538 25620 16268
rect 25676 16100 25732 16110
rect 25676 16006 25732 16044
rect 25564 15486 25566 15538
rect 25618 15486 25620 15538
rect 25340 15474 25396 15484
rect 25564 15474 25620 15486
rect 25676 15764 25732 15774
rect 25676 15428 25732 15708
rect 25788 15652 25844 16830
rect 26124 16772 26180 16782
rect 26124 16212 26180 16716
rect 26124 16146 26180 16156
rect 26236 16210 26292 16940
rect 26684 16324 26740 17164
rect 27244 17154 27300 17164
rect 27356 17444 27412 17454
rect 27132 17108 27188 17118
rect 27020 17106 27188 17108
rect 27020 17054 27134 17106
rect 27186 17054 27188 17106
rect 27020 17052 27188 17054
rect 26908 16884 26964 16894
rect 26908 16790 26964 16828
rect 26684 16258 26740 16268
rect 26796 16660 26852 16670
rect 26236 16158 26238 16210
rect 26290 16158 26292 16210
rect 26236 16146 26292 16158
rect 26684 16100 26740 16110
rect 26684 16006 26740 16044
rect 26124 15874 26180 15886
rect 26124 15822 26126 15874
rect 26178 15822 26180 15874
rect 26124 15652 26180 15822
rect 26348 15876 26404 15886
rect 26684 15876 26740 15886
rect 26348 15874 26628 15876
rect 26348 15822 26350 15874
rect 26402 15822 26628 15874
rect 26348 15820 26628 15822
rect 26348 15810 26404 15820
rect 25844 15596 25956 15652
rect 25788 15586 25844 15596
rect 25788 15428 25844 15438
rect 25676 15426 25844 15428
rect 25676 15374 25790 15426
rect 25842 15374 25844 15426
rect 25676 15372 25844 15374
rect 25228 15316 25284 15326
rect 25228 15222 25284 15260
rect 25452 15204 25508 15214
rect 25116 14130 25172 14140
rect 25228 15092 25284 15102
rect 25116 12964 25172 12974
rect 25116 12870 25172 12908
rect 25004 12852 25060 12862
rect 25004 12758 25060 12796
rect 24556 11508 24612 11518
rect 24556 11414 24612 11452
rect 24668 10836 24724 10846
rect 24668 10610 24724 10780
rect 24668 10558 24670 10610
rect 24722 10558 24724 10610
rect 24556 10052 24612 10062
rect 24556 9044 24612 9996
rect 24668 9940 24724 10558
rect 24668 9874 24724 9884
rect 24556 8950 24612 8988
rect 24332 8428 24500 8484
rect 23996 8260 24052 8270
rect 23996 8166 24052 8204
rect 23884 8082 23940 8092
rect 24220 7812 24276 7822
rect 23996 7700 24052 7710
rect 23996 7474 24052 7644
rect 23996 7422 23998 7474
rect 24050 7422 24052 7474
rect 23996 7410 24052 7422
rect 24108 7698 24164 7710
rect 24108 7646 24110 7698
rect 24162 7646 24164 7698
rect 23996 6692 24052 6702
rect 23996 6598 24052 6636
rect 24108 6580 24164 7646
rect 24220 7474 24276 7756
rect 24220 7422 24222 7474
rect 24274 7422 24276 7474
rect 24220 6804 24276 7422
rect 24332 6804 24388 8428
rect 24668 8260 24724 8270
rect 24444 8148 24500 8186
rect 24668 8166 24724 8204
rect 24444 8082 24500 8092
rect 24668 7700 24724 7710
rect 24780 7700 24836 12124
rect 25228 12292 25284 15036
rect 25340 13972 25396 13982
rect 25340 13878 25396 13916
rect 25340 12964 25396 12974
rect 25452 12964 25508 15148
rect 25788 15148 25844 15372
rect 25900 15428 25956 15596
rect 26124 15586 26180 15596
rect 25900 15362 25956 15372
rect 26460 15428 26516 15438
rect 26348 15316 26404 15326
rect 26348 15222 26404 15260
rect 25788 15092 25956 15148
rect 25564 14418 25620 14430
rect 25564 14366 25566 14418
rect 25618 14366 25620 14418
rect 25564 14084 25620 14366
rect 25564 13524 25620 14028
rect 25564 13458 25620 13468
rect 25564 13186 25620 13198
rect 25564 13134 25566 13186
rect 25618 13134 25620 13186
rect 25564 13076 25620 13134
rect 25564 13010 25620 13020
rect 25340 12962 25508 12964
rect 25340 12910 25342 12962
rect 25394 12910 25508 12962
rect 25340 12908 25508 12910
rect 25676 12964 25732 12974
rect 25340 12852 25396 12908
rect 25676 12870 25732 12908
rect 25340 12786 25396 12796
rect 25788 12404 25844 12414
rect 25900 12404 25956 15092
rect 26348 14756 26404 14766
rect 26124 14644 26180 14654
rect 26124 14532 26180 14588
rect 26124 14530 26292 14532
rect 26124 14478 26126 14530
rect 26178 14478 26292 14530
rect 26124 14476 26292 14478
rect 26124 14466 26180 14476
rect 26012 13746 26068 13758
rect 26012 13694 26014 13746
rect 26066 13694 26068 13746
rect 26012 13412 26068 13694
rect 26012 13346 26068 13356
rect 26236 13300 26292 14476
rect 26348 14530 26404 14700
rect 26348 14478 26350 14530
rect 26402 14478 26404 14530
rect 26348 14466 26404 14478
rect 26460 13746 26516 15372
rect 26572 13970 26628 15820
rect 26684 15782 26740 15820
rect 26684 15652 26740 15662
rect 26684 15538 26740 15596
rect 26684 15486 26686 15538
rect 26738 15486 26740 15538
rect 26684 15474 26740 15486
rect 26684 15314 26740 15326
rect 26684 15262 26686 15314
rect 26738 15262 26740 15314
rect 26684 15204 26740 15262
rect 26796 15316 26852 16604
rect 27020 16324 27076 17052
rect 27132 17042 27188 17052
rect 27356 16994 27412 17388
rect 27356 16942 27358 16994
rect 27410 16942 27412 16994
rect 27356 16930 27412 16942
rect 27132 16772 27188 16782
rect 27468 16772 27524 18172
rect 27580 18162 27636 18172
rect 27804 18004 27860 18732
rect 27916 18564 27972 18574
rect 28476 18564 28532 19740
rect 27916 18562 28532 18564
rect 27916 18510 27918 18562
rect 27970 18510 28532 18562
rect 27916 18508 28532 18510
rect 27916 18498 27972 18508
rect 27580 17948 27860 18004
rect 27580 17890 27636 17948
rect 27580 17838 27582 17890
rect 27634 17838 27636 17890
rect 27580 17826 27636 17838
rect 27916 17780 27972 17790
rect 27916 17778 28196 17780
rect 27916 17726 27918 17778
rect 27970 17726 28196 17778
rect 27916 17724 28196 17726
rect 27916 17714 27972 17724
rect 27916 17556 27972 17566
rect 27972 17500 28084 17556
rect 27916 17490 27972 17500
rect 27804 17444 27860 17454
rect 27580 17388 27804 17444
rect 27580 17108 27636 17388
rect 27804 17350 27860 17388
rect 27916 17108 27972 17118
rect 27580 17042 27636 17052
rect 27804 17106 27972 17108
rect 27804 17054 27918 17106
rect 27970 17054 27972 17106
rect 27804 17052 27972 17054
rect 27580 16884 27636 16894
rect 27580 16790 27636 16828
rect 27132 16770 27524 16772
rect 27132 16718 27134 16770
rect 27186 16718 27524 16770
rect 27132 16716 27524 16718
rect 27132 16706 27188 16716
rect 26796 15250 26852 15260
rect 26908 16268 27076 16324
rect 26684 15138 26740 15148
rect 26908 15090 26964 16268
rect 27020 16100 27076 16138
rect 27020 16034 27076 16044
rect 27244 16098 27300 16110
rect 27244 16046 27246 16098
rect 27298 16046 27300 16098
rect 27244 15988 27300 16046
rect 27804 16100 27860 17052
rect 27916 17042 27972 17052
rect 28028 16884 28084 17500
rect 27804 16034 27860 16044
rect 27916 16882 28084 16884
rect 27916 16830 28030 16882
rect 28082 16830 28084 16882
rect 27916 16828 28084 16830
rect 27916 16098 27972 16828
rect 28028 16818 28084 16828
rect 28140 16658 28196 17724
rect 28140 16606 28142 16658
rect 28194 16606 28196 16658
rect 28140 16594 28196 16606
rect 28252 17332 28308 17342
rect 28140 16324 28196 16334
rect 28140 16230 28196 16268
rect 27916 16046 27918 16098
rect 27970 16046 27972 16098
rect 27356 15988 27412 15998
rect 27244 15932 27356 15988
rect 27356 15922 27412 15932
rect 27468 15986 27524 15998
rect 27468 15934 27470 15986
rect 27522 15934 27524 15986
rect 27468 15652 27524 15934
rect 27468 15586 27524 15596
rect 27916 15540 27972 16046
rect 27580 15484 27972 15540
rect 28028 15988 28084 15998
rect 27132 15428 27188 15438
rect 27132 15314 27188 15372
rect 27468 15428 27524 15438
rect 27468 15334 27524 15372
rect 27132 15262 27134 15314
rect 27186 15262 27188 15314
rect 27132 15250 27188 15262
rect 26908 15038 26910 15090
rect 26962 15038 26964 15090
rect 26908 15026 26964 15038
rect 27580 14980 27636 15484
rect 28028 15426 28084 15932
rect 28028 15374 28030 15426
rect 28082 15374 28084 15426
rect 27244 14924 27636 14980
rect 27804 15314 27860 15326
rect 27804 15262 27806 15314
rect 27858 15262 27860 15314
rect 26796 14756 26852 14766
rect 26796 14662 26852 14700
rect 26572 13918 26574 13970
rect 26626 13918 26628 13970
rect 26572 13906 26628 13918
rect 27132 13972 27188 14010
rect 27132 13906 27188 13916
rect 26460 13694 26462 13746
rect 26514 13694 26516 13746
rect 26460 13682 26516 13694
rect 26796 13748 26852 13758
rect 26796 13654 26852 13692
rect 27132 13748 27188 13758
rect 27132 13654 27188 13692
rect 26348 13524 26404 13534
rect 26348 13430 26404 13468
rect 26908 13524 26964 13534
rect 26236 13244 26404 13300
rect 26236 13076 26292 13086
rect 26236 12982 26292 13020
rect 26124 12850 26180 12862
rect 26124 12798 26126 12850
rect 26178 12798 26180 12850
rect 26124 12740 26180 12798
rect 26124 12674 26180 12684
rect 25788 12402 25956 12404
rect 25788 12350 25790 12402
rect 25842 12350 25956 12402
rect 25788 12348 25956 12350
rect 25788 12338 25844 12348
rect 26348 12292 26404 13244
rect 26908 13074 26964 13468
rect 27244 13412 27300 14924
rect 27804 14868 27860 15262
rect 27356 14812 27860 14868
rect 27356 14754 27412 14812
rect 27356 14702 27358 14754
rect 27410 14702 27412 14754
rect 27356 14690 27412 14702
rect 27692 14532 27748 14542
rect 27692 14438 27748 14476
rect 28028 13972 28084 15374
rect 28140 15874 28196 15886
rect 28140 15822 28142 15874
rect 28194 15822 28196 15874
rect 28140 15316 28196 15822
rect 28252 15538 28308 17276
rect 28700 16994 28756 21308
rect 28924 20356 28980 24558
rect 29148 24724 29204 26348
rect 29484 26290 29540 26852
rect 29596 26852 29652 27694
rect 31500 27186 31556 27916
rect 31836 27906 31892 27916
rect 32172 28082 32228 28702
rect 32844 28700 33236 28756
rect 33292 28868 33348 28878
rect 32172 28030 32174 28082
rect 32226 28030 32228 28082
rect 31500 27134 31502 27186
rect 31554 27134 31556 27186
rect 31500 27122 31556 27134
rect 32172 27186 32228 28030
rect 32284 28642 32340 28654
rect 32284 28590 32286 28642
rect 32338 28590 32340 28642
rect 32284 27972 32340 28590
rect 32284 27906 32340 27916
rect 32396 28420 32452 28430
rect 32396 28082 32452 28364
rect 32396 28030 32398 28082
rect 32450 28030 32452 28082
rect 32172 27134 32174 27186
rect 32226 27134 32228 27186
rect 32172 27122 32228 27134
rect 31612 27076 31668 27086
rect 31612 26982 31668 27020
rect 32284 27076 32340 27086
rect 32284 26982 32340 27020
rect 29596 26786 29652 26796
rect 29708 26404 29764 26414
rect 32396 26404 32452 28030
rect 32508 27860 32564 27870
rect 32508 27766 32564 27804
rect 32844 27860 32900 28700
rect 33292 28642 33348 28812
rect 33404 28754 33460 29932
rect 33740 29652 33796 29662
rect 33740 29426 33796 29596
rect 33740 29374 33742 29426
rect 33794 29374 33796 29426
rect 33740 29362 33796 29374
rect 33516 29316 33572 29326
rect 33572 29260 33684 29316
rect 33516 29250 33572 29260
rect 33404 28702 33406 28754
rect 33458 28702 33460 28754
rect 33404 28690 33460 28702
rect 33292 28590 33294 28642
rect 33346 28590 33348 28642
rect 33292 28578 33348 28590
rect 33516 28644 33572 28654
rect 32956 28532 33012 28542
rect 32956 28438 33012 28476
rect 33180 27860 33236 27870
rect 32844 27858 33236 27860
rect 32844 27806 33182 27858
rect 33234 27806 33236 27858
rect 32844 27804 33236 27806
rect 32844 26908 32900 27804
rect 33180 27794 33236 27804
rect 33516 27636 33572 28588
rect 32956 27580 33572 27636
rect 33628 28642 33684 29260
rect 33852 28980 33908 30492
rect 34076 29652 34132 31614
rect 34076 29586 34132 29596
rect 34300 31668 34356 31678
rect 33964 29428 34020 29438
rect 33964 29334 34020 29372
rect 34300 29316 34356 31612
rect 34412 30100 34468 33964
rect 34748 33908 34804 33918
rect 34748 33234 34804 33852
rect 35084 33908 35140 33918
rect 34972 33684 35028 33694
rect 35084 33684 35140 33852
rect 35028 33628 35140 33684
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34972 33618 35028 33628
rect 35084 33346 35140 33628
rect 35084 33294 35086 33346
rect 35138 33294 35140 33346
rect 35084 33282 35140 33294
rect 34748 33182 34750 33234
rect 34802 33182 34804 33234
rect 34748 33170 34804 33182
rect 35420 33236 35476 33246
rect 35420 33142 35476 33180
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35532 32004 35588 34638
rect 35756 33348 35812 34748
rect 36428 35028 36484 35038
rect 36316 34692 36372 34702
rect 36092 34690 36372 34692
rect 36092 34638 36318 34690
rect 36370 34638 36372 34690
rect 36092 34636 36372 34638
rect 35980 34018 36036 34030
rect 35980 33966 35982 34018
rect 36034 33966 36036 34018
rect 35980 33796 36036 33966
rect 35980 33730 36036 33740
rect 35644 33346 35812 33348
rect 35644 33294 35758 33346
rect 35810 33294 35812 33346
rect 35644 33292 35812 33294
rect 35644 32786 35700 33292
rect 35756 33282 35812 33292
rect 35644 32734 35646 32786
rect 35698 32734 35700 32786
rect 35644 32722 35700 32734
rect 35532 31938 35588 31948
rect 36092 31892 36148 34636
rect 36316 34626 36372 34636
rect 36428 34354 36484 34972
rect 37884 35028 37940 35038
rect 37884 34802 37940 34972
rect 37884 34750 37886 34802
rect 37938 34750 37940 34802
rect 37884 34738 37940 34750
rect 37100 34692 37156 34702
rect 37100 34690 37268 34692
rect 37100 34638 37102 34690
rect 37154 34638 37268 34690
rect 37100 34636 37268 34638
rect 37100 34626 37156 34636
rect 36428 34302 36430 34354
rect 36482 34302 36484 34354
rect 36428 34290 36484 34302
rect 36540 34244 36596 34254
rect 36540 34150 36596 34188
rect 37100 34130 37156 34142
rect 37100 34078 37102 34130
rect 37154 34078 37156 34130
rect 36428 33908 36484 33918
rect 36428 33814 36484 33852
rect 37100 33572 37156 34078
rect 36988 33516 37156 33572
rect 37212 34018 37268 34636
rect 37212 33966 37214 34018
rect 37266 33966 37268 34018
rect 36316 33348 36372 33358
rect 36988 33348 37044 33516
rect 36316 33346 36932 33348
rect 36316 33294 36318 33346
rect 36370 33294 36932 33346
rect 36316 33292 36932 33294
rect 36316 33282 36372 33292
rect 36204 33236 36260 33246
rect 36204 33142 36260 33180
rect 36428 33124 36484 33134
rect 36428 33030 36484 33068
rect 36428 32788 36484 32798
rect 36204 31892 36260 31902
rect 36092 31836 36204 31892
rect 36260 31836 36372 31892
rect 36204 31798 36260 31836
rect 35644 31780 35700 31790
rect 34524 31556 34580 31566
rect 34524 31462 34580 31500
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 30212 35252 30222
rect 34636 30100 34692 30110
rect 34412 30098 34636 30100
rect 34412 30046 34414 30098
rect 34466 30046 34636 30098
rect 34412 30044 34636 30046
rect 34412 30034 34468 30044
rect 34524 29538 34580 29550
rect 34524 29486 34526 29538
rect 34578 29486 34580 29538
rect 34412 29316 34468 29326
rect 34300 29314 34468 29316
rect 34300 29262 34414 29314
rect 34466 29262 34468 29314
rect 34300 29260 34468 29262
rect 34412 29250 34468 29260
rect 34524 29316 34580 29486
rect 34524 29250 34580 29260
rect 34636 29204 34692 30044
rect 35196 29652 35252 30156
rect 35196 29558 35252 29596
rect 34748 29428 34804 29438
rect 34972 29428 35028 29438
rect 34748 29426 35028 29428
rect 34748 29374 34750 29426
rect 34802 29374 34974 29426
rect 35026 29374 35028 29426
rect 34748 29372 35028 29374
rect 34748 29362 34804 29372
rect 34972 29362 35028 29372
rect 35308 29428 35364 29438
rect 35308 29204 35364 29372
rect 34636 29148 34916 29204
rect 33852 28924 34244 28980
rect 33628 28590 33630 28642
rect 33682 28590 33684 28642
rect 32956 27186 33012 27580
rect 33628 27524 33684 28590
rect 33852 28756 33908 28766
rect 33852 28642 33908 28700
rect 33852 28590 33854 28642
rect 33906 28590 33908 28642
rect 33852 28578 33908 28590
rect 34076 28644 34132 28654
rect 34076 28550 34132 28588
rect 33740 28532 33796 28542
rect 33740 27636 33796 28476
rect 33964 27748 34020 27758
rect 33964 27746 34132 27748
rect 33964 27694 33966 27746
rect 34018 27694 34132 27746
rect 33964 27692 34132 27694
rect 33964 27682 34020 27692
rect 33740 27580 33908 27636
rect 33628 27458 33684 27468
rect 33740 27300 33796 27310
rect 33740 27206 33796 27244
rect 32956 27134 32958 27186
rect 33010 27134 33012 27186
rect 32956 27122 33012 27134
rect 33292 27076 33348 27114
rect 33516 27076 33572 27086
rect 33292 27010 33348 27020
rect 33404 27074 33684 27076
rect 33404 27022 33518 27074
rect 33570 27022 33684 27074
rect 33404 27020 33684 27022
rect 33404 26908 33460 27020
rect 33516 27010 33572 27020
rect 32732 26852 32900 26908
rect 33180 26852 33236 26862
rect 29708 26402 29876 26404
rect 29708 26350 29710 26402
rect 29762 26350 29876 26402
rect 29708 26348 29876 26350
rect 29708 26338 29764 26348
rect 29484 26238 29486 26290
rect 29538 26238 29540 26290
rect 29372 25396 29428 25406
rect 29372 25302 29428 25340
rect 29372 24948 29428 24958
rect 29484 24948 29540 26238
rect 29708 25506 29764 25518
rect 29708 25454 29710 25506
rect 29762 25454 29764 25506
rect 29596 25396 29652 25406
rect 29708 25396 29764 25454
rect 29652 25340 29764 25396
rect 29596 25330 29652 25340
rect 29372 24946 29540 24948
rect 29372 24894 29374 24946
rect 29426 24894 29540 24946
rect 29372 24892 29540 24894
rect 29372 24882 29428 24892
rect 29148 24276 29204 24668
rect 29148 24210 29204 24220
rect 29148 24052 29204 24062
rect 29148 24050 29652 24052
rect 29148 23998 29150 24050
rect 29202 23998 29652 24050
rect 29148 23996 29652 23998
rect 29148 23986 29204 23996
rect 29372 23828 29428 23838
rect 29372 23378 29428 23772
rect 29372 23326 29374 23378
rect 29426 23326 29428 23378
rect 29372 23314 29428 23326
rect 29148 23156 29204 23166
rect 29148 23154 29316 23156
rect 29148 23102 29150 23154
rect 29202 23102 29316 23154
rect 29148 23100 29316 23102
rect 29148 23090 29204 23100
rect 29260 22594 29316 23100
rect 29596 22596 29652 23996
rect 29820 22596 29876 26348
rect 32396 26402 32676 26404
rect 32396 26350 32398 26402
rect 32450 26350 32676 26402
rect 32396 26348 32676 26350
rect 32396 26338 32452 26348
rect 31612 26292 31668 26302
rect 31612 26198 31668 26236
rect 32060 26292 32116 26302
rect 32060 26198 32116 26236
rect 30492 26180 30548 26190
rect 30492 25618 30548 26124
rect 32508 26068 32564 26078
rect 32508 25974 32564 26012
rect 30492 25566 30494 25618
rect 30546 25566 30548 25618
rect 30492 25554 30548 25566
rect 32620 25618 32676 26348
rect 32620 25566 32622 25618
rect 32674 25566 32676 25618
rect 32620 25554 32676 25566
rect 32620 25396 32676 25406
rect 32060 25284 32116 25294
rect 32060 24834 32116 25228
rect 32508 24948 32564 24958
rect 32508 24854 32564 24892
rect 32620 24946 32676 25340
rect 32620 24894 32622 24946
rect 32674 24894 32676 24946
rect 32620 24882 32676 24894
rect 32060 24782 32062 24834
rect 32114 24782 32116 24834
rect 32060 24770 32116 24782
rect 32284 24722 32340 24734
rect 32284 24670 32286 24722
rect 32338 24670 32340 24722
rect 32284 24612 32340 24670
rect 32284 24546 32340 24556
rect 29260 22542 29262 22594
rect 29314 22542 29316 22594
rect 29260 22530 29316 22542
rect 29372 22594 29652 22596
rect 29372 22542 29598 22594
rect 29650 22542 29652 22594
rect 29372 22540 29652 22542
rect 29372 22372 29428 22540
rect 29596 22530 29652 22540
rect 29708 22540 29876 22596
rect 30156 24276 30212 24286
rect 29148 22316 29428 22372
rect 29148 21698 29204 22316
rect 29148 21646 29150 21698
rect 29202 21646 29204 21698
rect 29148 21634 29204 21646
rect 29708 21812 29764 22540
rect 29820 22260 29876 22270
rect 29820 22166 29876 22204
rect 29036 21364 29092 21374
rect 29036 21270 29092 21308
rect 29708 21028 29764 21756
rect 30044 21700 30100 21710
rect 29708 20962 29764 20972
rect 29932 21644 30044 21700
rect 29148 20916 29204 20926
rect 29148 20802 29204 20860
rect 29148 20750 29150 20802
rect 29202 20750 29204 20802
rect 29148 20738 29204 20750
rect 29484 20578 29540 20590
rect 29484 20526 29486 20578
rect 29538 20526 29540 20578
rect 29484 20356 29540 20526
rect 28924 20300 29204 20356
rect 28924 20132 28980 20142
rect 28924 20038 28980 20076
rect 28924 18676 28980 18686
rect 28924 18338 28980 18620
rect 28924 18286 28926 18338
rect 28978 18286 28980 18338
rect 28924 18274 28980 18286
rect 28700 16942 28702 16994
rect 28754 16942 28756 16994
rect 28700 16930 28756 16942
rect 28252 15486 28254 15538
rect 28306 15486 28308 15538
rect 28252 15474 28308 15486
rect 28364 16882 28420 16894
rect 28364 16830 28366 16882
rect 28418 16830 28420 16882
rect 28364 15986 28420 16830
rect 28364 15934 28366 15986
rect 28418 15934 28420 15986
rect 28364 15540 28420 15934
rect 28364 15474 28420 15484
rect 28588 15986 28644 15998
rect 28588 15934 28590 15986
rect 28642 15934 28644 15986
rect 28252 15316 28308 15326
rect 28140 15314 28308 15316
rect 28140 15262 28254 15314
rect 28306 15262 28308 15314
rect 28140 15260 28308 15262
rect 28252 15250 28308 15260
rect 28364 15316 28420 15326
rect 28364 15222 28420 15260
rect 28588 15148 28644 15934
rect 28588 15092 28756 15148
rect 28364 14530 28420 14542
rect 28364 14478 28366 14530
rect 28418 14478 28420 14530
rect 28364 14084 28420 14478
rect 28364 14018 28420 14028
rect 28476 14418 28532 14430
rect 28476 14366 28478 14418
rect 28530 14366 28532 14418
rect 27692 13916 28084 13972
rect 27692 13858 27748 13916
rect 27692 13806 27694 13858
rect 27746 13806 27748 13858
rect 27692 13794 27748 13806
rect 27916 13748 27972 13758
rect 27916 13654 27972 13692
rect 27468 13636 27524 13646
rect 27468 13542 27524 13580
rect 28476 13524 28532 14366
rect 28476 13458 28532 13468
rect 27356 13412 27412 13422
rect 27244 13356 27356 13412
rect 27356 13346 27412 13356
rect 26908 13022 26910 13074
rect 26962 13022 26964 13074
rect 26908 13010 26964 13022
rect 27244 13188 27300 13198
rect 25228 12236 25508 12292
rect 25228 10276 25284 12236
rect 25340 12066 25396 12078
rect 25340 12014 25342 12066
rect 25394 12014 25396 12066
rect 25340 11956 25396 12014
rect 25340 10836 25396 11900
rect 25452 11396 25508 12236
rect 26236 12236 26404 12292
rect 26460 12962 26516 12974
rect 26460 12910 26462 12962
rect 26514 12910 26516 12962
rect 25452 11302 25508 11340
rect 25900 11396 25956 11406
rect 26236 11396 26292 12236
rect 26348 12068 26404 12078
rect 26348 11844 26404 12012
rect 26460 11956 26516 12910
rect 27244 12964 27300 13132
rect 27356 13188 27412 13198
rect 27916 13188 27972 13198
rect 27356 13186 27972 13188
rect 27356 13134 27358 13186
rect 27410 13134 27918 13186
rect 27970 13134 27972 13186
rect 27356 13132 27972 13134
rect 27356 13122 27412 13132
rect 27916 13122 27972 13132
rect 27356 12964 27412 12974
rect 27244 12962 27412 12964
rect 27244 12910 27358 12962
rect 27410 12910 27412 12962
rect 27244 12908 27412 12910
rect 27356 12898 27412 12908
rect 27580 12964 27636 12974
rect 26796 12852 26852 12862
rect 26460 11890 26516 11900
rect 26572 12850 26852 12852
rect 26572 12798 26798 12850
rect 26850 12798 26852 12850
rect 26572 12796 26852 12798
rect 26348 11778 26404 11788
rect 26460 11396 26516 11406
rect 25900 11394 26068 11396
rect 25900 11342 25902 11394
rect 25954 11342 26068 11394
rect 25900 11340 26068 11342
rect 26236 11394 26516 11396
rect 26236 11342 26462 11394
rect 26514 11342 26516 11394
rect 26236 11340 26516 11342
rect 25900 11330 25956 11340
rect 25340 10780 25844 10836
rect 25676 10610 25732 10622
rect 25676 10558 25678 10610
rect 25730 10558 25732 10610
rect 25004 9940 25060 9950
rect 25004 9846 25060 9884
rect 25228 9604 25284 10220
rect 25228 9538 25284 9548
rect 25340 10500 25396 10510
rect 25676 10500 25732 10558
rect 25340 10498 25732 10500
rect 25340 10446 25342 10498
rect 25394 10446 25732 10498
rect 25340 10444 25732 10446
rect 24724 7644 24836 7700
rect 25228 9044 25284 9054
rect 25340 9044 25396 10444
rect 25788 10276 25844 10780
rect 26012 10388 26068 11340
rect 26460 11330 26516 11340
rect 26124 11172 26180 11182
rect 26124 11170 26516 11172
rect 26124 11118 26126 11170
rect 26178 11118 26516 11170
rect 26124 11116 26516 11118
rect 26124 11106 26180 11116
rect 26460 10722 26516 11116
rect 26460 10670 26462 10722
rect 26514 10670 26516 10722
rect 26460 10658 26516 10670
rect 26012 10332 26516 10388
rect 25788 10220 26180 10276
rect 26012 10052 26068 10062
rect 26012 9938 26068 9996
rect 26012 9886 26014 9938
rect 26066 9886 26068 9938
rect 26012 9874 26068 9886
rect 25564 9604 25620 9614
rect 25564 9492 25620 9548
rect 25564 9436 25956 9492
rect 25788 9156 25844 9166
rect 25284 8988 25396 9044
rect 25452 9154 25844 9156
rect 25452 9102 25790 9154
rect 25842 9102 25844 9154
rect 25452 9100 25844 9102
rect 25228 8370 25284 8988
rect 25340 8484 25396 8494
rect 25452 8484 25508 9100
rect 25788 9090 25844 9100
rect 25900 9156 25956 9436
rect 25900 9090 25956 9100
rect 26012 9268 26068 9278
rect 26012 9042 26068 9212
rect 26012 8990 26014 9042
rect 26066 8990 26068 9042
rect 25564 8932 25620 8942
rect 26012 8932 26068 8990
rect 25564 8930 26068 8932
rect 25564 8878 25566 8930
rect 25618 8878 26068 8930
rect 25564 8876 26068 8878
rect 25564 8708 25620 8876
rect 25564 8642 25620 8652
rect 25396 8428 25508 8484
rect 25340 8418 25396 8428
rect 25228 8318 25230 8370
rect 25282 8318 25284 8370
rect 25228 8260 25284 8318
rect 25676 8260 25732 8270
rect 25228 8258 25732 8260
rect 25228 8206 25678 8258
rect 25730 8206 25732 8258
rect 25228 8204 25732 8206
rect 25228 7700 25284 8204
rect 25676 8194 25732 8204
rect 25340 7700 25396 7710
rect 25228 7698 25396 7700
rect 25228 7646 25342 7698
rect 25394 7646 25396 7698
rect 25228 7644 25396 7646
rect 24668 7606 24724 7644
rect 25340 7634 25396 7644
rect 24892 6804 24948 6814
rect 24332 6748 24500 6804
rect 24220 6738 24276 6748
rect 24108 6524 24276 6580
rect 23548 5906 23828 5908
rect 23548 5854 23550 5906
rect 23602 5854 23828 5906
rect 23548 5852 23828 5854
rect 23884 6244 23940 6254
rect 23548 5842 23604 5852
rect 23212 5682 23268 5694
rect 23212 5630 23214 5682
rect 23266 5630 23268 5682
rect 23212 5348 23268 5630
rect 23212 5282 23268 5292
rect 22148 5180 22260 5236
rect 21532 5070 21534 5122
rect 21586 5070 21588 5122
rect 21532 5058 21588 5070
rect 21756 5124 21812 5134
rect 21756 5010 21812 5068
rect 22092 5122 22148 5180
rect 22092 5070 22094 5122
rect 22146 5070 22148 5122
rect 22092 5058 22148 5070
rect 22876 5124 22932 5134
rect 22876 5030 22932 5068
rect 21756 4958 21758 5010
rect 21810 4958 21812 5010
rect 21756 4946 21812 4958
rect 20860 4286 20862 4338
rect 20914 4286 20916 4338
rect 20860 4274 20916 4286
rect 21644 4226 21700 4238
rect 21644 4174 21646 4226
rect 21698 4174 21700 4226
rect 21644 4116 21700 4174
rect 23772 4228 23828 4238
rect 23884 4228 23940 6188
rect 24220 6020 24276 6524
rect 24332 6578 24388 6590
rect 24332 6526 24334 6578
rect 24386 6526 24388 6578
rect 24332 6244 24388 6526
rect 24332 6178 24388 6188
rect 24220 5906 24276 5964
rect 24332 6020 24388 6030
rect 24444 6020 24500 6748
rect 24892 6710 24948 6748
rect 26124 6692 26180 10220
rect 26460 10050 26516 10332
rect 26460 9998 26462 10050
rect 26514 9998 26516 10050
rect 26460 9986 26516 9998
rect 26124 6626 26180 6636
rect 26236 9492 26292 9502
rect 26236 6132 26292 9436
rect 26572 9492 26628 12796
rect 26796 12786 26852 12796
rect 27020 12850 27076 12862
rect 27020 12798 27022 12850
rect 27074 12798 27076 12850
rect 27020 12628 27076 12798
rect 27020 12562 27076 12572
rect 27020 12180 27076 12190
rect 27020 12086 27076 12124
rect 26908 12068 26964 12078
rect 26908 11788 26964 12012
rect 26796 11732 26964 11788
rect 27468 12066 27524 12078
rect 27468 12014 27470 12066
rect 27522 12014 27524 12066
rect 26684 11396 26740 11406
rect 26684 11302 26740 11340
rect 26796 10052 26852 11732
rect 27468 11396 27524 12014
rect 27580 11618 27636 12908
rect 28028 12964 28084 12974
rect 28028 12850 28084 12908
rect 28028 12798 28030 12850
rect 28082 12798 28084 12850
rect 28028 12786 28084 12798
rect 28252 12850 28308 12862
rect 28252 12798 28254 12850
rect 28306 12798 28308 12850
rect 27916 12180 27972 12190
rect 27916 12086 27972 12124
rect 27580 11566 27582 11618
rect 27634 11566 27636 11618
rect 27580 11554 27636 11566
rect 27468 11330 27524 11340
rect 27244 11284 27300 11294
rect 27244 11282 27412 11284
rect 27244 11230 27246 11282
rect 27298 11230 27412 11282
rect 27244 11228 27412 11230
rect 27244 11218 27300 11228
rect 26852 9996 27076 10052
rect 26796 9986 26852 9996
rect 26572 9426 26628 9436
rect 26796 9826 26852 9838
rect 26796 9774 26798 9826
rect 26850 9774 26852 9826
rect 26796 9380 26852 9774
rect 26796 9324 26964 9380
rect 26460 9044 26516 9054
rect 26684 9044 26740 9054
rect 26516 9042 26740 9044
rect 26516 8990 26686 9042
rect 26738 8990 26740 9042
rect 26516 8988 26740 8990
rect 26460 8978 26516 8988
rect 26684 8978 26740 8988
rect 26908 8932 26964 9324
rect 27020 9042 27076 9996
rect 27020 8990 27022 9042
rect 27074 8990 27076 9042
rect 27020 8978 27076 8990
rect 27356 9826 27412 11228
rect 27356 9774 27358 9826
rect 27410 9774 27412 9826
rect 26908 8866 26964 8876
rect 27244 8930 27300 8942
rect 27244 8878 27246 8930
rect 27298 8878 27300 8930
rect 26460 8708 26516 8718
rect 26460 8370 26516 8652
rect 26684 8708 26740 8718
rect 26740 8652 26852 8708
rect 26684 8642 26740 8652
rect 26460 8318 26462 8370
rect 26514 8318 26516 8370
rect 26460 8306 26516 8318
rect 26572 8484 26628 8494
rect 26348 6132 26404 6142
rect 26236 6130 26404 6132
rect 26236 6078 26350 6130
rect 26402 6078 26404 6130
rect 26236 6076 26404 6078
rect 26348 6066 26404 6076
rect 24332 6018 25060 6020
rect 24332 5966 24334 6018
rect 24386 5966 25060 6018
rect 24332 5964 25060 5966
rect 24332 5954 24388 5964
rect 24220 5854 24222 5906
rect 24274 5854 24276 5906
rect 24220 5842 24276 5854
rect 25004 5234 25060 5964
rect 25004 5182 25006 5234
rect 25058 5182 25060 5234
rect 25004 5170 25060 5182
rect 25340 5794 25396 5806
rect 25340 5742 25342 5794
rect 25394 5742 25396 5794
rect 25340 5122 25396 5742
rect 25340 5070 25342 5122
rect 25394 5070 25396 5122
rect 24220 5012 24276 5022
rect 24220 4562 24276 4956
rect 25340 5012 25396 5070
rect 25788 5794 25844 5806
rect 25788 5742 25790 5794
rect 25842 5742 25844 5794
rect 25788 5012 25844 5742
rect 26236 5796 26292 5806
rect 26236 5702 26292 5740
rect 25396 4956 25844 5012
rect 26124 5010 26180 5022
rect 26124 4958 26126 5010
rect 26178 4958 26180 5010
rect 25340 4946 25396 4956
rect 24220 4510 24222 4562
rect 24274 4510 24276 4562
rect 24220 4498 24276 4510
rect 25676 4564 25732 4956
rect 25676 4470 25732 4508
rect 26012 4564 26068 4574
rect 26124 4564 26180 4958
rect 26012 4562 26180 4564
rect 26012 4510 26014 4562
rect 26066 4510 26180 4562
rect 26012 4508 26180 4510
rect 26012 4498 26068 4508
rect 23772 4226 23940 4228
rect 23772 4174 23774 4226
rect 23826 4174 23940 4226
rect 23772 4172 23940 4174
rect 26236 4338 26292 4350
rect 26236 4286 26238 4338
rect 26290 4286 26292 4338
rect 23772 4162 23828 4172
rect 20748 4060 21700 4116
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 26236 3778 26292 4286
rect 26236 3726 26238 3778
rect 26290 3726 26292 3778
rect 26236 3714 26292 3726
rect 26572 3778 26628 8428
rect 26796 7698 26852 8652
rect 26796 7646 26798 7698
rect 26850 7646 26852 7698
rect 26796 7634 26852 7646
rect 27132 8372 27188 8382
rect 27132 7474 27188 8316
rect 27132 7422 27134 7474
rect 27186 7422 27188 7474
rect 26908 6578 26964 6590
rect 26908 6526 26910 6578
rect 26962 6526 26964 6578
rect 26796 6132 26852 6142
rect 26908 6132 26964 6526
rect 26796 6130 26964 6132
rect 26796 6078 26798 6130
rect 26850 6078 26964 6130
rect 26796 6076 26964 6078
rect 26796 6066 26852 6076
rect 27132 5906 27188 7422
rect 27244 6692 27300 8878
rect 27356 7586 27412 9774
rect 27692 11282 27748 11294
rect 27692 11230 27694 11282
rect 27746 11230 27748 11282
rect 27692 10500 27748 11230
rect 28252 10724 28308 12798
rect 28252 10658 28308 10668
rect 27580 9716 27636 9726
rect 27692 9716 27748 10444
rect 28588 10500 28644 10510
rect 28588 10406 28644 10444
rect 27580 9714 27748 9716
rect 27580 9662 27582 9714
rect 27634 9662 27748 9714
rect 27580 9660 27748 9662
rect 27580 9650 27636 9660
rect 28588 9268 28644 9278
rect 28700 9268 28756 15092
rect 29148 14868 29204 20300
rect 29484 20290 29540 20300
rect 29820 20356 29876 20366
rect 29932 20356 29988 21644
rect 30044 21606 30100 21644
rect 29876 20300 29988 20356
rect 29484 20130 29540 20142
rect 29484 20078 29486 20130
rect 29538 20078 29540 20130
rect 29484 20020 29540 20078
rect 29540 19964 29764 20020
rect 29484 19954 29540 19964
rect 29260 19796 29316 19806
rect 29260 19702 29316 19740
rect 29708 19234 29764 19964
rect 29708 19182 29710 19234
rect 29762 19182 29764 19234
rect 29708 19170 29764 19182
rect 29820 19122 29876 20300
rect 30044 20244 30100 20254
rect 30044 20130 30100 20188
rect 30044 20078 30046 20130
rect 30098 20078 30100 20130
rect 30044 20066 30100 20078
rect 30156 19908 30212 24220
rect 32508 24052 32564 24062
rect 32732 24052 32788 26852
rect 33180 26758 33236 26796
rect 33292 26852 33460 26908
rect 33628 26964 33684 27020
rect 33628 26898 33684 26908
rect 33516 26852 33572 26862
rect 33068 26290 33124 26302
rect 33068 26238 33070 26290
rect 33122 26238 33124 26290
rect 33068 26068 33124 26238
rect 33292 26290 33348 26852
rect 33292 26238 33294 26290
rect 33346 26238 33348 26290
rect 33292 26226 33348 26238
rect 33516 26292 33572 26796
rect 33516 26198 33572 26236
rect 33628 26516 33684 26526
rect 33628 26290 33684 26460
rect 33628 26238 33630 26290
rect 33682 26238 33684 26290
rect 33180 26180 33236 26190
rect 33180 26086 33236 26124
rect 33068 25732 33124 26012
rect 33068 25676 33348 25732
rect 33068 25506 33124 25518
rect 33068 25454 33070 25506
rect 33122 25454 33124 25506
rect 33068 25284 33124 25454
rect 33068 24836 33124 25228
rect 33068 24834 33236 24836
rect 33068 24782 33070 24834
rect 33122 24782 33236 24834
rect 33068 24780 33236 24782
rect 33068 24770 33124 24780
rect 32060 24050 32788 24052
rect 32060 23998 32510 24050
rect 32562 23998 32788 24050
rect 32060 23996 32788 23998
rect 32060 23938 32116 23996
rect 32508 23986 32564 23996
rect 32060 23886 32062 23938
rect 32114 23886 32116 23938
rect 32060 23874 32116 23886
rect 31276 23828 31332 23838
rect 31276 23734 31332 23772
rect 30716 23044 30772 23054
rect 30380 22258 30436 22270
rect 30380 22206 30382 22258
rect 30434 22206 30436 22258
rect 30380 21700 30436 22206
rect 30492 21812 30548 21822
rect 30492 21718 30548 21756
rect 30380 21634 30436 21644
rect 30716 20804 30772 22988
rect 32732 22484 32788 23996
rect 33180 23938 33236 24780
rect 33292 24724 33348 25676
rect 33628 25396 33684 26238
rect 33628 25330 33684 25340
rect 33852 25394 33908 27580
rect 33964 27524 34020 27534
rect 33964 27074 34020 27468
rect 33964 27022 33966 27074
rect 34018 27022 34020 27074
rect 33964 25618 34020 27022
rect 34076 26852 34132 27692
rect 34188 27300 34244 28924
rect 34748 28756 34804 28766
rect 34412 28642 34468 28654
rect 34412 28590 34414 28642
rect 34466 28590 34468 28642
rect 34188 27234 34244 27244
rect 34300 28418 34356 28430
rect 34300 28366 34302 28418
rect 34354 28366 34356 28418
rect 34300 27074 34356 28366
rect 34300 27022 34302 27074
rect 34354 27022 34356 27074
rect 34300 27010 34356 27022
rect 34076 26786 34132 26796
rect 34412 26516 34468 28590
rect 34748 28642 34804 28700
rect 34748 28590 34750 28642
rect 34802 28590 34804 28642
rect 34748 27074 34804 28590
rect 34748 27022 34750 27074
rect 34802 27022 34804 27074
rect 34748 27010 34804 27022
rect 34524 26964 34580 27002
rect 34524 26852 34804 26908
rect 34412 26450 34468 26460
rect 34524 26404 34580 26414
rect 34524 26402 34692 26404
rect 34524 26350 34526 26402
rect 34578 26350 34692 26402
rect 34524 26348 34692 26350
rect 34524 26338 34580 26348
rect 34076 26292 34132 26302
rect 34076 26290 34244 26292
rect 34076 26238 34078 26290
rect 34130 26238 34244 26290
rect 34076 26236 34244 26238
rect 34076 26226 34132 26236
rect 33964 25566 33966 25618
rect 34018 25566 34020 25618
rect 33964 25554 34020 25566
rect 33852 25342 33854 25394
rect 33906 25342 33908 25394
rect 33852 25330 33908 25342
rect 33292 24658 33348 24668
rect 33852 25172 33908 25182
rect 33852 24722 33908 25116
rect 33852 24670 33854 24722
rect 33906 24670 33908 24722
rect 33852 24658 33908 24670
rect 34076 24724 34132 24734
rect 34076 24630 34132 24668
rect 33180 23886 33182 23938
rect 33234 23886 33236 23938
rect 33180 23874 33236 23886
rect 33516 24612 33572 24622
rect 33404 23826 33460 23838
rect 33404 23774 33406 23826
rect 33458 23774 33460 23826
rect 33404 23156 33460 23774
rect 33516 23828 33572 24556
rect 33628 24052 33684 24062
rect 34076 24052 34132 24062
rect 33628 24050 34132 24052
rect 33628 23998 33630 24050
rect 33682 23998 34078 24050
rect 34130 23998 34132 24050
rect 33628 23996 34132 23998
rect 33628 23986 33684 23996
rect 34076 23986 34132 23996
rect 34188 24050 34244 26236
rect 34412 26290 34468 26302
rect 34412 26238 34414 26290
rect 34466 26238 34468 26290
rect 34188 23998 34190 24050
rect 34242 23998 34244 24050
rect 34188 23986 34244 23998
rect 34300 25060 34356 25070
rect 33740 23828 33796 23838
rect 34300 23828 34356 25004
rect 34412 24836 34468 26238
rect 34524 26068 34580 26078
rect 34524 25974 34580 26012
rect 34636 25394 34692 26348
rect 34636 25342 34638 25394
rect 34690 25342 34692 25394
rect 34636 24948 34692 25342
rect 34468 24780 34580 24836
rect 34412 24770 34468 24780
rect 33516 23826 33796 23828
rect 33516 23774 33742 23826
rect 33794 23774 33796 23826
rect 33516 23772 33796 23774
rect 33740 23604 33796 23772
rect 33964 23826 34356 23828
rect 33964 23774 34302 23826
rect 34354 23774 34356 23826
rect 33964 23772 34356 23774
rect 33852 23604 33908 23614
rect 33740 23548 33852 23604
rect 33852 23538 33908 23548
rect 33964 23378 34020 23772
rect 34300 23762 34356 23772
rect 33964 23326 33966 23378
rect 34018 23326 34020 23378
rect 33964 23314 34020 23326
rect 34300 23380 34356 23390
rect 34300 23286 34356 23324
rect 34524 23378 34580 24780
rect 34524 23326 34526 23378
rect 34578 23326 34580 23378
rect 34524 23314 34580 23326
rect 34188 23268 34244 23278
rect 34188 23174 34244 23212
rect 33516 23156 33572 23166
rect 33404 23100 33516 23156
rect 33516 23090 33572 23100
rect 34636 23044 34692 24892
rect 34748 23716 34804 26852
rect 34748 23650 34804 23660
rect 34748 23266 34804 23278
rect 34748 23214 34750 23266
rect 34802 23214 34804 23266
rect 34748 23156 34804 23214
rect 34748 23090 34804 23100
rect 34636 22978 34692 22988
rect 32732 22418 32788 22428
rect 34188 22484 34244 22494
rect 34188 22390 34244 22428
rect 33292 22370 33348 22382
rect 33292 22318 33294 22370
rect 33346 22318 33348 22370
rect 33292 21924 33348 22318
rect 34860 21924 34916 29148
rect 35084 29148 35364 29204
rect 35084 28754 35140 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35084 28702 35086 28754
rect 35138 28702 35140 28754
rect 35084 28690 35140 28702
rect 35532 28530 35588 28542
rect 35532 28478 35534 28530
rect 35586 28478 35588 28530
rect 35084 28418 35140 28430
rect 35084 28366 35086 28418
rect 35138 28366 35140 28418
rect 35084 27972 35140 28366
rect 35308 28420 35364 28430
rect 35308 28326 35364 28364
rect 35084 27906 35140 27916
rect 35532 27860 35588 28478
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35532 26908 35588 27804
rect 35644 27074 35700 31724
rect 35980 30882 36036 30894
rect 35980 30830 35982 30882
rect 36034 30830 36036 30882
rect 35756 30212 35812 30222
rect 35756 30118 35812 30156
rect 35868 30212 35924 30222
rect 35980 30212 36036 30830
rect 35868 30210 36036 30212
rect 35868 30158 35870 30210
rect 35922 30158 36036 30210
rect 35868 30156 36036 30158
rect 35868 30146 35924 30156
rect 36316 28754 36372 31836
rect 36428 30994 36484 32732
rect 36876 32674 36932 33292
rect 36876 32622 36878 32674
rect 36930 32622 36932 32674
rect 36876 32610 36932 32622
rect 36988 32564 37044 33292
rect 37100 33346 37156 33358
rect 37100 33294 37102 33346
rect 37154 33294 37156 33346
rect 37100 33124 37156 33294
rect 37100 32788 37156 33068
rect 37100 32722 37156 32732
rect 37212 33236 37268 33966
rect 37772 33236 37828 33246
rect 37100 32564 37156 32574
rect 36988 32562 37156 32564
rect 36988 32510 37102 32562
rect 37154 32510 37156 32562
rect 36988 32508 37156 32510
rect 37212 32564 37268 33180
rect 37324 33234 37828 33236
rect 37324 33182 37774 33234
rect 37826 33182 37828 33234
rect 37324 33180 37828 33182
rect 37324 32786 37380 33180
rect 37772 33170 37828 33180
rect 37324 32734 37326 32786
rect 37378 32734 37380 32786
rect 37324 32722 37380 32734
rect 37436 32564 37492 32574
rect 37212 32562 37492 32564
rect 37212 32510 37438 32562
rect 37490 32510 37492 32562
rect 37212 32508 37492 32510
rect 37100 32498 37156 32508
rect 37436 32498 37492 32508
rect 36428 30942 36430 30994
rect 36482 30942 36484 30994
rect 36428 30930 36484 30942
rect 36652 32340 36708 32350
rect 36316 28702 36318 28754
rect 36370 28702 36372 28754
rect 36316 28690 36372 28702
rect 36428 28420 36484 28430
rect 36092 27860 36148 27870
rect 36092 27746 36148 27804
rect 36428 27858 36484 28364
rect 36540 27972 36596 27982
rect 36540 27878 36596 27916
rect 36428 27806 36430 27858
rect 36482 27806 36484 27858
rect 36428 27794 36484 27806
rect 36092 27694 36094 27746
rect 36146 27694 36148 27746
rect 36092 27682 36148 27694
rect 35644 27022 35646 27074
rect 35698 27022 35700 27074
rect 35644 27010 35700 27022
rect 35980 27074 36036 27086
rect 35980 27022 35982 27074
rect 36034 27022 36036 27074
rect 35084 26852 35588 26908
rect 35980 26908 36036 27022
rect 36428 27076 36484 27086
rect 36204 26964 36260 27002
rect 36428 26982 36484 27020
rect 35644 26852 35700 26862
rect 35980 26852 36148 26908
rect 36204 26898 36260 26908
rect 35084 25508 35140 26852
rect 35644 26758 35700 26796
rect 36092 26514 36148 26852
rect 36092 26462 36094 26514
rect 36146 26462 36148 26514
rect 36092 26450 36148 26462
rect 35308 26292 35364 26302
rect 35308 26198 35364 26236
rect 35532 26290 35588 26302
rect 35532 26238 35534 26290
rect 35586 26238 35588 26290
rect 35532 26068 35588 26238
rect 35980 26292 36036 26302
rect 35980 26198 36036 26236
rect 36204 26290 36260 26302
rect 36204 26238 36206 26290
rect 36258 26238 36260 26290
rect 35756 26180 35812 26190
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34972 25452 35140 25508
rect 34972 25172 35028 25452
rect 35532 25396 35588 26012
rect 34972 25106 35028 25116
rect 35084 25340 35588 25396
rect 35644 26178 35812 26180
rect 35644 26126 35758 26178
rect 35810 26126 35812 26178
rect 35644 26124 35812 26126
rect 35084 23940 35140 25340
rect 35644 25060 35700 26124
rect 35756 26114 35812 26124
rect 35532 25004 35700 25060
rect 36204 25506 36260 26238
rect 36204 25454 36206 25506
rect 36258 25454 36260 25506
rect 35420 24836 35476 24846
rect 35420 24742 35476 24780
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35420 24164 35476 24174
rect 35420 24070 35476 24108
rect 35532 24052 35588 25004
rect 36204 24948 36260 25454
rect 36540 26290 36596 26302
rect 36540 26238 36542 26290
rect 36594 26238 36596 26290
rect 36204 24892 36484 24948
rect 35644 24834 35700 24846
rect 35644 24782 35646 24834
rect 35698 24782 35700 24834
rect 35644 24164 35700 24782
rect 36204 24722 36260 24734
rect 36204 24670 36206 24722
rect 36258 24670 36260 24722
rect 35756 24500 35812 24510
rect 35756 24498 36148 24500
rect 35756 24446 35758 24498
rect 35810 24446 36148 24498
rect 35756 24444 36148 24446
rect 35756 24434 35812 24444
rect 35644 24108 35812 24164
rect 35196 23940 35252 23950
rect 35084 23938 35252 23940
rect 35084 23886 35198 23938
rect 35250 23886 35252 23938
rect 35084 23884 35252 23886
rect 35196 23874 35252 23884
rect 34972 23826 35028 23838
rect 34972 23774 34974 23826
rect 35026 23774 35028 23826
rect 34972 22596 35028 23774
rect 35084 23154 35140 23166
rect 35084 23102 35086 23154
rect 35138 23102 35140 23154
rect 35084 23044 35140 23102
rect 35532 23156 35588 23996
rect 35644 23938 35700 23950
rect 35644 23886 35646 23938
rect 35698 23886 35700 23938
rect 35644 23716 35700 23886
rect 35644 23650 35700 23660
rect 35644 23156 35700 23166
rect 35532 23154 35700 23156
rect 35532 23102 35646 23154
rect 35698 23102 35700 23154
rect 35532 23100 35700 23102
rect 35644 23090 35700 23100
rect 35756 23156 35812 24108
rect 35868 23828 35924 23838
rect 35868 23734 35924 23772
rect 35756 23090 35812 23100
rect 35980 23714 36036 23726
rect 35980 23662 35982 23714
rect 36034 23662 36036 23714
rect 35084 22978 35140 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34972 22530 35028 22540
rect 35532 22484 35588 22494
rect 34972 21924 35028 21934
rect 34860 21868 34972 21924
rect 31948 21698 32004 21710
rect 31948 21646 31950 21698
rect 32002 21646 32004 21698
rect 31836 20916 31892 20926
rect 31948 20916 32004 21646
rect 32284 21588 32340 21598
rect 33180 21588 33236 21598
rect 32284 21586 33236 21588
rect 32284 21534 32286 21586
rect 32338 21534 33182 21586
rect 33234 21534 33236 21586
rect 32284 21532 33236 21534
rect 32284 21522 32340 21532
rect 33180 21522 33236 21532
rect 31836 20914 32004 20916
rect 31836 20862 31838 20914
rect 31890 20862 32004 20914
rect 31836 20860 32004 20862
rect 32396 21364 32452 21374
rect 31836 20850 31892 20860
rect 31052 20804 31108 20814
rect 30716 20802 31108 20804
rect 30716 20750 30718 20802
rect 30770 20750 31054 20802
rect 31106 20750 31108 20802
rect 30716 20748 31108 20750
rect 30716 20738 30772 20748
rect 31052 20738 31108 20748
rect 30828 20132 30884 20142
rect 30828 20130 31108 20132
rect 30828 20078 30830 20130
rect 30882 20078 31108 20130
rect 30828 20076 31108 20078
rect 30828 20066 30884 20076
rect 30604 20020 30660 20030
rect 30604 20018 30772 20020
rect 30604 19966 30606 20018
rect 30658 19966 30772 20018
rect 30604 19964 30772 19966
rect 30604 19954 30660 19964
rect 29820 19070 29822 19122
rect 29874 19070 29876 19122
rect 29820 19058 29876 19070
rect 29932 19852 30212 19908
rect 29820 17666 29876 17678
rect 29820 17614 29822 17666
rect 29874 17614 29876 17666
rect 29820 17444 29876 17614
rect 29820 16884 29876 17388
rect 29596 16548 29652 16558
rect 29596 16322 29652 16492
rect 29596 16270 29598 16322
rect 29650 16270 29652 16322
rect 29596 16258 29652 16270
rect 29820 15986 29876 16828
rect 29820 15934 29822 15986
rect 29874 15934 29876 15986
rect 29820 15922 29876 15934
rect 29260 15874 29316 15886
rect 29260 15822 29262 15874
rect 29314 15822 29316 15874
rect 29260 15428 29316 15822
rect 29260 15362 29316 15372
rect 29932 15148 29988 19852
rect 30716 19458 30772 19964
rect 30716 19406 30718 19458
rect 30770 19406 30772 19458
rect 30716 19394 30772 19406
rect 30380 19236 30436 19246
rect 30156 19234 30436 19236
rect 30156 19182 30382 19234
rect 30434 19182 30436 19234
rect 30156 19180 30436 19182
rect 30156 18676 30212 19180
rect 30380 19170 30436 19180
rect 30156 17890 30212 18620
rect 31052 18562 31108 20076
rect 31052 18510 31054 18562
rect 31106 18510 31108 18562
rect 31052 18498 31108 18510
rect 31836 19234 31892 19246
rect 31836 19182 31838 19234
rect 31890 19182 31892 19234
rect 31836 18450 31892 19182
rect 31836 18398 31838 18450
rect 31890 18398 31892 18450
rect 31836 18340 31892 18398
rect 31836 18274 31892 18284
rect 32284 18340 32340 18350
rect 32284 18246 32340 18284
rect 30156 17838 30158 17890
rect 30210 17838 30212 17890
rect 30156 17826 30212 17838
rect 30044 17442 30100 17454
rect 30044 17390 30046 17442
rect 30098 17390 30100 17442
rect 30044 16324 30100 17390
rect 30828 16994 30884 17006
rect 30828 16942 30830 16994
rect 30882 16942 30884 16994
rect 30604 16884 30660 16894
rect 30604 16882 30772 16884
rect 30604 16830 30606 16882
rect 30658 16830 30772 16882
rect 30604 16828 30772 16830
rect 30604 16818 30660 16828
rect 30044 16258 30100 16268
rect 30380 16212 30436 16222
rect 30380 15986 30436 16156
rect 30380 15934 30382 15986
rect 30434 15934 30436 15986
rect 30380 15922 30436 15934
rect 30716 15540 30772 16828
rect 30828 16436 30884 16942
rect 31276 16996 31332 17006
rect 31276 16902 31332 16940
rect 31948 16994 32004 17006
rect 31948 16942 31950 16994
rect 32002 16942 32004 16994
rect 31948 16884 32004 16942
rect 32396 16994 32452 21308
rect 33068 20132 33124 20142
rect 32508 20130 33124 20132
rect 32508 20078 33070 20130
rect 33122 20078 33124 20130
rect 32508 20076 33124 20078
rect 32508 19346 32564 20076
rect 33068 20066 33124 20076
rect 32508 19294 32510 19346
rect 32562 19294 32564 19346
rect 32508 19282 32564 19294
rect 33292 18564 33348 21868
rect 34972 21858 35028 21868
rect 35532 21812 35588 22428
rect 35980 22260 36036 23662
rect 36092 22594 36148 24444
rect 36204 23828 36260 24670
rect 36316 24164 36372 24174
rect 36316 24050 36372 24108
rect 36316 23998 36318 24050
rect 36370 23998 36372 24050
rect 36316 23986 36372 23998
rect 36204 23762 36260 23772
rect 36428 23604 36484 24892
rect 36540 23940 36596 26238
rect 36652 24164 36708 32284
rect 37996 32228 38052 35196
rect 38108 35026 38164 35038
rect 38108 34974 38110 35026
rect 38162 34974 38164 35026
rect 38108 34244 38164 34974
rect 38108 34178 38164 34188
rect 38220 33906 38276 35646
rect 38332 35812 38388 35822
rect 38332 35586 38388 35756
rect 38332 35534 38334 35586
rect 38386 35534 38388 35586
rect 38332 35522 38388 35534
rect 38780 35700 38836 37886
rect 38892 37492 38948 39788
rect 39900 39732 39956 39742
rect 40012 39732 40068 40350
rect 39900 39730 40068 39732
rect 39900 39678 39902 39730
rect 39954 39678 40068 39730
rect 39900 39676 40068 39678
rect 40236 40068 40292 40078
rect 39900 39620 39956 39676
rect 39900 39554 39956 39564
rect 39228 38722 39284 38734
rect 39228 38670 39230 38722
rect 39282 38670 39284 38722
rect 39228 38668 39284 38670
rect 39228 38612 39732 38668
rect 39676 38050 39732 38612
rect 39676 37998 39678 38050
rect 39730 37998 39732 38050
rect 39340 37940 39396 37950
rect 38892 37426 38948 37436
rect 39004 37938 39396 37940
rect 39004 37886 39342 37938
rect 39394 37886 39396 37938
rect 39004 37884 39396 37886
rect 39004 36594 39060 37884
rect 39340 37874 39396 37884
rect 39004 36542 39006 36594
rect 39058 36542 39060 36594
rect 39004 36530 39060 36542
rect 39452 37826 39508 37838
rect 39452 37774 39454 37826
rect 39506 37774 39508 37826
rect 39452 36596 39508 37774
rect 39452 36530 39508 36540
rect 39564 36482 39620 36494
rect 39564 36430 39566 36482
rect 39618 36430 39620 36482
rect 38780 35252 38836 35644
rect 39116 35700 39172 35710
rect 39452 35700 39508 35710
rect 39116 35698 39508 35700
rect 39116 35646 39118 35698
rect 39170 35646 39454 35698
rect 39506 35646 39508 35698
rect 39116 35644 39508 35646
rect 39116 35634 39172 35644
rect 39452 35634 39508 35644
rect 38780 35186 38836 35196
rect 39340 34916 39396 34926
rect 39564 34916 39620 36430
rect 39676 36484 39732 37998
rect 39788 37604 39844 37614
rect 39788 37266 39844 37548
rect 40236 37490 40292 40012
rect 40236 37438 40238 37490
rect 40290 37438 40292 37490
rect 40236 37426 40292 37438
rect 40684 39508 40740 44380
rect 40796 44370 40852 44380
rect 40796 43538 40852 43550
rect 40796 43486 40798 43538
rect 40850 43486 40852 43538
rect 40796 43316 40852 43486
rect 40908 43540 40964 45838
rect 41244 45836 41468 45892
rect 41020 45106 41076 45118
rect 41020 45054 41022 45106
rect 41074 45054 41076 45106
rect 41020 44994 41076 45054
rect 41020 44942 41022 44994
rect 41074 44942 41076 44994
rect 41020 44930 41076 44942
rect 41244 44322 41300 45836
rect 41468 45826 41524 45836
rect 44044 45892 44100 45902
rect 44044 45798 44100 45836
rect 44380 45332 44436 46062
rect 41468 45220 41524 45230
rect 41468 45126 41524 45164
rect 42364 45220 42420 45230
rect 42364 45126 42420 45164
rect 41580 45108 41636 45118
rect 41580 45014 41636 45052
rect 41692 45108 41748 45118
rect 41916 45108 41972 45118
rect 41692 45106 41972 45108
rect 41692 45054 41694 45106
rect 41746 45054 41918 45106
rect 41970 45054 41972 45106
rect 41692 45052 41972 45054
rect 41244 44270 41246 44322
rect 41298 44270 41300 44322
rect 41244 44258 41300 44270
rect 41356 43764 41412 43774
rect 41692 43764 41748 45052
rect 41916 45042 41972 45052
rect 42476 45108 42532 45118
rect 44380 45108 44436 45276
rect 44492 45892 44548 45902
rect 44492 45330 44548 45836
rect 44940 45892 44996 45902
rect 44940 45798 44996 45836
rect 45612 45778 45668 47404
rect 45836 47458 45892 47516
rect 45836 47406 45838 47458
rect 45890 47406 45892 47458
rect 45836 47394 45892 47406
rect 46060 47460 46116 48300
rect 46396 48132 46452 48142
rect 46396 47682 46452 48076
rect 46396 47630 46398 47682
rect 46450 47630 46452 47682
rect 46396 47618 46452 47630
rect 46508 47908 46564 47918
rect 46060 47366 46116 47404
rect 46508 47458 46564 47852
rect 46508 47406 46510 47458
rect 46562 47406 46564 47458
rect 46508 47394 46564 47406
rect 46620 47234 46676 48860
rect 46956 48850 47012 48860
rect 47740 48692 47796 50428
rect 47964 50484 48020 51100
rect 48076 50596 48132 51436
rect 48860 51378 48916 51390
rect 48860 51326 48862 51378
rect 48914 51326 48916 51378
rect 48860 51268 48916 51326
rect 48860 51202 48916 51212
rect 48188 51044 48244 51054
rect 48188 50706 48244 50988
rect 48188 50654 48190 50706
rect 48242 50654 48244 50706
rect 48188 50642 48244 50654
rect 48076 50502 48132 50540
rect 48300 50596 48356 50606
rect 48300 50502 48356 50540
rect 47964 50418 48020 50428
rect 48524 50482 48580 50494
rect 48524 50430 48526 50482
rect 48578 50430 48580 50482
rect 48524 50260 48580 50430
rect 48972 50428 49028 52332
rect 49868 52386 49924 52782
rect 49868 52334 49870 52386
rect 49922 52334 49924 52386
rect 49868 52322 49924 52334
rect 49420 52276 49476 52286
rect 49420 52182 49476 52220
rect 49980 52276 50036 52892
rect 51436 52948 51492 53788
rect 51548 53778 51604 53788
rect 50540 52388 50596 52398
rect 49980 52210 50036 52220
rect 50316 52386 50596 52388
rect 50316 52334 50542 52386
rect 50594 52334 50596 52386
rect 50316 52332 50596 52334
rect 49756 52164 49812 52174
rect 49196 52052 49252 52062
rect 49084 51996 49196 52052
rect 49084 51602 49140 51996
rect 49196 51986 49252 51996
rect 49420 52052 49476 52062
rect 49756 52052 49812 52108
rect 49980 52052 50036 52062
rect 49084 51550 49086 51602
rect 49138 51550 49140 51602
rect 49084 51538 49140 51550
rect 49308 51938 49364 51950
rect 49308 51886 49310 51938
rect 49362 51886 49364 51938
rect 49308 50596 49364 51886
rect 49420 51490 49476 51996
rect 49420 51438 49422 51490
rect 49474 51438 49476 51490
rect 49420 51426 49476 51438
rect 49532 52050 49812 52052
rect 49532 51998 49758 52050
rect 49810 51998 49812 52050
rect 49532 51996 49812 51998
rect 49308 50502 49364 50540
rect 49420 50932 49476 50942
rect 49420 50482 49476 50876
rect 49420 50430 49422 50482
rect 49474 50430 49476 50482
rect 48972 50372 49252 50428
rect 49420 50418 49476 50430
rect 48580 50204 49028 50260
rect 48524 50194 48580 50204
rect 48748 49924 48804 49934
rect 48748 49830 48804 49868
rect 48972 49810 49028 50204
rect 48972 49758 48974 49810
rect 49026 49758 49028 49810
rect 48972 49746 49028 49758
rect 49084 49812 49140 49822
rect 49084 49698 49140 49756
rect 49084 49646 49086 49698
rect 49138 49646 49140 49698
rect 49084 49634 49140 49646
rect 49196 49476 49252 50372
rect 48972 49420 49252 49476
rect 48972 49028 49028 49420
rect 49084 49252 49140 49262
rect 49140 49196 49252 49252
rect 49084 49158 49140 49196
rect 48972 48972 49140 49028
rect 46956 48356 47012 48366
rect 46620 47182 46622 47234
rect 46674 47182 46676 47234
rect 46620 47170 46676 47182
rect 46732 48300 46956 48356
rect 46060 47124 46116 47134
rect 45836 46676 45892 46686
rect 45836 46582 45892 46620
rect 46060 46674 46116 47068
rect 46060 46622 46062 46674
rect 46114 46622 46116 46674
rect 46060 46610 46116 46622
rect 46172 46564 46228 46574
rect 46172 46470 46228 46508
rect 46620 46564 46676 46574
rect 46620 46470 46676 46508
rect 45724 46452 45780 46462
rect 45724 46358 45780 46396
rect 45836 46228 45892 46238
rect 45836 45890 45892 46172
rect 45836 45838 45838 45890
rect 45890 45838 45892 45890
rect 45836 45826 45892 45838
rect 46620 45892 46676 45902
rect 46732 45892 46788 48300
rect 46956 48262 47012 48300
rect 47292 48020 47348 48030
rect 47180 47460 47236 47470
rect 47180 46786 47236 47404
rect 47292 47458 47348 47964
rect 47292 47406 47294 47458
rect 47346 47406 47348 47458
rect 47292 47394 47348 47406
rect 47628 47460 47684 47470
rect 47740 47460 47796 48636
rect 48748 48802 48804 48814
rect 48748 48750 48750 48802
rect 48802 48750 48804 48802
rect 47964 48244 48020 48254
rect 47964 47570 48020 48188
rect 48636 48244 48692 48254
rect 48748 48244 48804 48750
rect 48692 48188 48804 48244
rect 48972 48242 49028 48254
rect 48972 48190 48974 48242
rect 49026 48190 49028 48242
rect 48636 48150 48692 48188
rect 47964 47518 47966 47570
rect 48018 47518 48020 47570
rect 47964 47506 48020 47518
rect 48188 48130 48244 48142
rect 48188 48078 48190 48130
rect 48242 48078 48244 48130
rect 48188 48020 48244 48078
rect 48860 48132 48916 48142
rect 48860 48038 48916 48076
rect 47628 47458 47796 47460
rect 47628 47406 47630 47458
rect 47682 47406 47796 47458
rect 47628 47404 47796 47406
rect 47628 47394 47684 47404
rect 47180 46734 47182 46786
rect 47234 46734 47236 46786
rect 47180 46722 47236 46734
rect 47404 46788 47460 46798
rect 47068 46674 47124 46686
rect 47068 46622 47070 46674
rect 47122 46622 47124 46674
rect 47068 46228 47124 46622
rect 47404 46674 47460 46732
rect 47404 46622 47406 46674
rect 47458 46622 47460 46674
rect 47404 46610 47460 46622
rect 47068 46162 47124 46172
rect 47292 46452 47348 46462
rect 47292 46002 47348 46396
rect 47292 45950 47294 46002
rect 47346 45950 47348 46002
rect 47292 45938 47348 45950
rect 46676 45836 46788 45892
rect 46620 45798 46676 45836
rect 48188 45780 48244 47964
rect 48972 47684 49028 48190
rect 49084 47908 49140 48972
rect 49196 48468 49252 49196
rect 49532 49140 49588 51996
rect 49756 51986 49812 51996
rect 49868 51996 49980 52052
rect 49868 51938 49924 51996
rect 49980 51986 50036 51996
rect 50204 52052 50260 52062
rect 49868 51886 49870 51938
rect 49922 51886 49924 51938
rect 49868 51874 49924 51886
rect 49868 51492 49924 51502
rect 49756 51436 49868 51492
rect 49756 51378 49812 51436
rect 49868 51426 49924 51436
rect 49756 51326 49758 51378
rect 49810 51326 49812 51378
rect 49756 51314 49812 51326
rect 49980 51378 50036 51390
rect 49980 51326 49982 51378
rect 50034 51326 50036 51378
rect 49868 51266 49924 51278
rect 49868 51214 49870 51266
rect 49922 51214 49924 51266
rect 49868 51156 49924 51214
rect 49868 51090 49924 51100
rect 49868 50820 49924 50830
rect 49980 50820 50036 51326
rect 50204 51156 50260 51996
rect 49644 50818 50036 50820
rect 49644 50766 49870 50818
rect 49922 50766 50036 50818
rect 49644 50764 50036 50766
rect 50092 51100 50260 51156
rect 50316 51156 50372 52332
rect 50540 52322 50596 52332
rect 50652 52388 50708 52398
rect 50540 52164 50596 52174
rect 50652 52164 50708 52332
rect 50540 52162 50708 52164
rect 50540 52110 50542 52162
rect 50594 52110 50708 52162
rect 50540 52108 50708 52110
rect 50764 52164 50820 52174
rect 50540 52098 50596 52108
rect 50764 52070 50820 52108
rect 51100 52050 51156 52062
rect 51100 51998 51102 52050
rect 51154 51998 51156 52050
rect 50988 51940 51044 51950
rect 50988 51846 51044 51884
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 51100 51716 51156 51998
rect 51436 52050 51492 52892
rect 51884 52276 51940 52286
rect 51884 52162 51940 52220
rect 51884 52110 51886 52162
rect 51938 52110 51940 52162
rect 51884 52098 51940 52110
rect 51436 51998 51438 52050
rect 51490 51998 51492 52050
rect 51436 51986 51492 51998
rect 51324 51940 51380 51950
rect 50556 51706 50820 51716
rect 50876 51660 51156 51716
rect 51212 51938 51380 51940
rect 51212 51886 51326 51938
rect 51378 51886 51380 51938
rect 51212 51884 51380 51886
rect 50876 51492 50932 51660
rect 51212 51604 51268 51884
rect 51324 51874 51380 51884
rect 51660 51940 51716 51950
rect 52444 51940 52500 51950
rect 51660 51938 51828 51940
rect 51660 51886 51662 51938
rect 51714 51886 51828 51938
rect 51660 51884 51828 51886
rect 51660 51874 51716 51884
rect 49644 50594 49700 50764
rect 49868 50754 49924 50764
rect 49644 50542 49646 50594
rect 49698 50542 49700 50594
rect 49644 50530 49700 50542
rect 49980 50484 50036 50494
rect 49868 49810 49924 49822
rect 49868 49758 49870 49810
rect 49922 49758 49924 49810
rect 49868 49476 49924 49758
rect 49980 49698 50036 50428
rect 50092 50482 50148 51100
rect 50316 51090 50372 51100
rect 50764 51378 50820 51390
rect 50764 51326 50766 51378
rect 50818 51326 50820 51378
rect 50204 50706 50260 50718
rect 50204 50654 50206 50706
rect 50258 50654 50260 50706
rect 50204 50596 50260 50654
rect 50764 50708 50820 51326
rect 50764 50642 50820 50652
rect 50540 50596 50596 50606
rect 50204 50594 50596 50596
rect 50204 50542 50542 50594
rect 50594 50542 50596 50594
rect 50204 50540 50596 50542
rect 50540 50530 50596 50540
rect 50876 50594 50932 51436
rect 50988 51548 51268 51604
rect 50988 51266 51044 51548
rect 51660 51380 51716 51390
rect 51660 51286 51716 51324
rect 51324 51268 51380 51278
rect 50988 51214 50990 51266
rect 51042 51214 51044 51266
rect 50988 51202 51044 51214
rect 51100 51266 51380 51268
rect 51100 51214 51326 51266
rect 51378 51214 51380 51266
rect 51100 51212 51380 51214
rect 51100 50818 51156 51212
rect 51324 51202 51380 51212
rect 51772 51268 51828 51884
rect 52444 51490 52500 51884
rect 52444 51438 52446 51490
rect 52498 51438 52500 51490
rect 52444 51426 52500 51438
rect 51772 51202 51828 51212
rect 52668 51380 52724 51390
rect 51100 50766 51102 50818
rect 51154 50766 51156 50818
rect 51100 50754 51156 50766
rect 50876 50542 50878 50594
rect 50930 50542 50932 50594
rect 50092 50430 50094 50482
rect 50146 50430 50148 50482
rect 50092 50418 50148 50430
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 49980 49646 49982 49698
rect 50034 49646 50036 49698
rect 49980 49634 50036 49646
rect 49532 49074 49588 49084
rect 49644 49420 49924 49476
rect 49308 48916 49364 48926
rect 49644 48916 49700 49420
rect 49308 48914 49700 48916
rect 49308 48862 49310 48914
rect 49362 48862 49700 48914
rect 49308 48860 49700 48862
rect 49756 49252 49812 49262
rect 49756 48914 49812 49196
rect 50540 49252 50596 49262
rect 50876 49252 50932 50542
rect 51212 50594 51268 50606
rect 51212 50542 51214 50594
rect 51266 50542 51268 50594
rect 50596 49196 50932 49252
rect 50988 49698 51044 49710
rect 50988 49646 50990 49698
rect 51042 49646 51044 49698
rect 50540 49158 50596 49196
rect 49868 49140 49924 49150
rect 50988 49140 51044 49646
rect 51212 49252 51268 50542
rect 52668 50594 52724 51324
rect 54572 51268 54628 51278
rect 54572 51174 54628 51212
rect 55580 50708 55636 50718
rect 55580 50614 55636 50652
rect 52668 50542 52670 50594
rect 52722 50542 52724 50594
rect 52668 50530 52724 50542
rect 51324 50484 51380 50494
rect 51324 50370 51380 50428
rect 53452 50484 53508 50494
rect 53452 50390 53508 50428
rect 51324 50318 51326 50370
rect 51378 50318 51380 50370
rect 51324 50306 51380 50318
rect 51212 49196 51716 49252
rect 49868 49028 49924 49084
rect 50876 49084 51380 49140
rect 49980 49028 50036 49038
rect 49868 49026 50260 49028
rect 49868 48974 49982 49026
rect 50034 48974 50260 49026
rect 49868 48972 50260 48974
rect 49980 48962 50036 48972
rect 49756 48862 49758 48914
rect 49810 48862 49812 48914
rect 49308 48850 49364 48860
rect 49196 48412 49364 48468
rect 49084 47842 49140 47852
rect 49196 48242 49252 48254
rect 49196 48190 49198 48242
rect 49250 48190 49252 48242
rect 48524 47628 49028 47684
rect 48524 47572 48580 47628
rect 49196 47572 49252 48190
rect 48300 47460 48356 47470
rect 48300 47366 48356 47404
rect 48524 47458 48580 47516
rect 48972 47516 49252 47572
rect 48524 47406 48526 47458
rect 48578 47406 48580 47458
rect 48524 47394 48580 47406
rect 48748 47460 48804 47470
rect 48972 47460 49028 47516
rect 48748 47458 49028 47460
rect 48748 47406 48750 47458
rect 48802 47406 49028 47458
rect 48748 47404 49028 47406
rect 48748 47348 48804 47404
rect 48748 47282 48804 47292
rect 49084 47348 49140 47358
rect 49308 47348 49364 48412
rect 49084 47346 49364 47348
rect 49084 47294 49086 47346
rect 49138 47294 49364 47346
rect 49084 47292 49364 47294
rect 48636 47234 48692 47246
rect 48636 47182 48638 47234
rect 48690 47182 48692 47234
rect 48636 47124 48692 47182
rect 48636 47058 48692 47068
rect 49084 46788 49140 47292
rect 49140 46732 49252 46788
rect 49084 46722 49140 46732
rect 48860 46564 48916 46574
rect 48860 46470 48916 46508
rect 49196 45892 49252 46732
rect 49308 46676 49364 46686
rect 49420 46676 49476 48860
rect 49756 48850 49812 48862
rect 49644 48468 49700 48478
rect 49644 47684 49700 48412
rect 50092 48354 50148 48366
rect 50092 48302 50094 48354
rect 50146 48302 50148 48354
rect 49756 48242 49812 48254
rect 49756 48190 49758 48242
rect 49810 48190 49812 48242
rect 49756 48020 49812 48190
rect 49756 47954 49812 47964
rect 50092 47908 50148 48302
rect 50092 47842 50148 47852
rect 49644 47570 49700 47628
rect 50204 47682 50260 48972
rect 50652 49026 50708 49038
rect 50652 48974 50654 49026
rect 50706 48974 50708 49026
rect 50652 48804 50708 48974
rect 50876 49026 50932 49084
rect 50876 48974 50878 49026
rect 50930 48974 50932 49026
rect 50876 48962 50932 48974
rect 50988 48916 51044 48926
rect 50988 48914 51268 48916
rect 50988 48862 50990 48914
rect 51042 48862 51268 48914
rect 50988 48860 51268 48862
rect 50988 48850 51044 48860
rect 50652 48748 50932 48804
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50652 48468 50708 48478
rect 50540 48356 50596 48366
rect 50540 48244 50596 48300
rect 50204 47630 50206 47682
rect 50258 47630 50260 47682
rect 50204 47618 50260 47630
rect 50428 48242 50596 48244
rect 50428 48190 50542 48242
rect 50594 48190 50596 48242
rect 50428 48188 50596 48190
rect 49644 47518 49646 47570
rect 49698 47518 49700 47570
rect 49644 47506 49700 47518
rect 49868 47460 49924 47470
rect 49868 47366 49924 47404
rect 50316 47460 50372 47470
rect 49308 46674 49476 46676
rect 49308 46622 49310 46674
rect 49362 46622 49476 46674
rect 49308 46620 49476 46622
rect 49756 46676 49812 46686
rect 50092 46676 50148 46686
rect 49756 46674 50148 46676
rect 49756 46622 49758 46674
rect 49810 46622 50094 46674
rect 50146 46622 50148 46674
rect 49756 46620 50148 46622
rect 49308 46116 49364 46620
rect 49756 46610 49812 46620
rect 50092 46610 50148 46620
rect 50316 46674 50372 47404
rect 50316 46622 50318 46674
rect 50370 46622 50372 46674
rect 50316 46610 50372 46622
rect 50428 46452 50484 48188
rect 50540 48178 50596 48188
rect 50652 48020 50708 48412
rect 50876 48132 50932 48748
rect 51212 48354 51268 48860
rect 51324 48468 51380 49084
rect 51324 48402 51380 48412
rect 51436 48802 51492 48814
rect 51436 48750 51438 48802
rect 51490 48750 51492 48802
rect 51212 48302 51214 48354
rect 51266 48302 51268 48354
rect 51212 48290 51268 48302
rect 51436 48356 51492 48750
rect 51436 48290 51492 48300
rect 51548 48132 51604 48142
rect 50876 48076 51380 48132
rect 50652 47460 50708 47964
rect 51324 47570 51380 48076
rect 51324 47518 51326 47570
rect 51378 47518 51380 47570
rect 51324 47506 51380 47518
rect 51548 47684 51604 48076
rect 51212 47460 51268 47470
rect 50652 47458 51156 47460
rect 50652 47406 50654 47458
rect 50706 47406 51156 47458
rect 50652 47404 51156 47406
rect 50652 47394 50708 47404
rect 50876 47236 50932 47246
rect 50876 47234 51044 47236
rect 50876 47182 50878 47234
rect 50930 47182 51044 47234
rect 50876 47180 51044 47182
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50876 46900 50932 47180
rect 50988 47012 51044 47180
rect 50988 46946 51044 46956
rect 50540 46844 50932 46900
rect 51100 46898 51156 47404
rect 51212 47366 51268 47404
rect 51548 47458 51604 47628
rect 51548 47406 51550 47458
rect 51602 47406 51604 47458
rect 51548 47394 51604 47406
rect 51660 47012 51716 49196
rect 53340 48132 53396 48142
rect 53340 48038 53396 48076
rect 51660 46946 51716 46956
rect 51100 46846 51102 46898
rect 51154 46846 51156 46898
rect 50540 46676 50596 46844
rect 51100 46834 51156 46846
rect 50540 46582 50596 46620
rect 49308 46050 49364 46060
rect 50092 46396 50484 46452
rect 50652 46450 50708 46462
rect 50652 46398 50654 46450
rect 50706 46398 50708 46450
rect 49420 46002 49476 46014
rect 49420 45950 49422 46002
rect 49474 45950 49476 46002
rect 49420 45892 49476 45950
rect 49196 45836 49476 45892
rect 45612 45726 45614 45778
rect 45666 45726 45668 45778
rect 45612 45714 45668 45726
rect 47628 45724 48244 45780
rect 44492 45278 44494 45330
rect 44546 45278 44548 45330
rect 44492 45266 44548 45278
rect 44380 45052 44548 45108
rect 42476 45014 42532 45052
rect 42140 44994 42196 45006
rect 42140 44942 42142 44994
rect 42194 44942 42196 44994
rect 42140 44548 42196 44942
rect 41916 44492 42196 44548
rect 42364 44884 42420 44894
rect 41916 44434 41972 44492
rect 41916 44382 41918 44434
rect 41970 44382 41972 44434
rect 41916 44370 41972 44382
rect 41356 43762 41748 43764
rect 41356 43710 41358 43762
rect 41410 43710 41748 43762
rect 41356 43708 41748 43710
rect 41804 44100 41860 44110
rect 41356 43698 41412 43708
rect 41804 43652 41860 44044
rect 42364 43764 42420 44828
rect 44156 44100 44212 44110
rect 44156 44006 44212 44044
rect 42028 43708 42420 43764
rect 41692 43596 41860 43652
rect 41916 43650 41972 43662
rect 41916 43598 41918 43650
rect 41970 43598 41972 43650
rect 41244 43540 41300 43550
rect 40908 43484 41244 43540
rect 41244 43446 41300 43484
rect 41468 43538 41524 43550
rect 41468 43486 41470 43538
rect 41522 43486 41524 43538
rect 41468 43428 41524 43486
rect 41468 43362 41524 43372
rect 40796 43250 40852 43260
rect 41132 42868 41188 42878
rect 41132 42754 41188 42812
rect 41132 42702 41134 42754
rect 41186 42702 41188 42754
rect 41132 42690 41188 42702
rect 41692 42754 41748 43596
rect 41692 42702 41694 42754
rect 41746 42702 41748 42754
rect 41692 42690 41748 42702
rect 41804 42644 41860 42654
rect 41916 42644 41972 43598
rect 42028 42868 42084 43708
rect 42364 43650 42420 43708
rect 42364 43598 42366 43650
rect 42418 43598 42420 43650
rect 42364 43586 42420 43598
rect 42140 43540 42196 43550
rect 42140 43446 42196 43484
rect 43260 43540 43316 43550
rect 42252 43426 42308 43438
rect 42252 43374 42254 43426
rect 42306 43374 42308 43426
rect 42140 42868 42196 42878
rect 42028 42866 42196 42868
rect 42028 42814 42142 42866
rect 42194 42814 42196 42866
rect 42028 42812 42196 42814
rect 42140 42802 42196 42812
rect 41804 42642 41972 42644
rect 41804 42590 41806 42642
rect 41858 42590 41972 42642
rect 41804 42588 41972 42590
rect 41804 42308 41860 42588
rect 41804 42242 41860 42252
rect 42252 42196 42308 43374
rect 42364 42756 42420 42766
rect 42364 42754 42868 42756
rect 42364 42702 42366 42754
rect 42418 42702 42868 42754
rect 42364 42700 42868 42702
rect 42364 42690 42420 42700
rect 42700 42530 42756 42542
rect 42700 42478 42702 42530
rect 42754 42478 42756 42530
rect 42700 42308 42756 42478
rect 42140 42140 42308 42196
rect 42364 42252 42756 42308
rect 42028 41188 42084 41198
rect 42028 41094 42084 41132
rect 41580 41076 41636 41086
rect 41580 40982 41636 41020
rect 41468 40962 41524 40974
rect 41468 40910 41470 40962
rect 41522 40910 41524 40962
rect 41468 40628 41524 40910
rect 41692 40964 41748 40974
rect 41692 40870 41748 40908
rect 41916 40628 41972 40638
rect 41468 40572 41916 40628
rect 41356 40404 41412 40414
rect 41356 40310 41412 40348
rect 41916 40402 41972 40572
rect 41916 40350 41918 40402
rect 41970 40350 41972 40402
rect 41916 40338 41972 40350
rect 42140 40404 42196 42140
rect 42252 41972 42308 41982
rect 42364 41972 42420 42252
rect 42812 42196 42868 42700
rect 42252 41970 42420 41972
rect 42252 41918 42254 41970
rect 42306 41918 42420 41970
rect 42252 41916 42420 41918
rect 42700 42140 42868 42196
rect 42252 41906 42308 41916
rect 42476 41074 42532 41086
rect 42476 41022 42478 41074
rect 42530 41022 42532 41074
rect 42476 40964 42532 41022
rect 42476 40898 42532 40908
rect 42252 40404 42308 40414
rect 42140 40402 42420 40404
rect 42140 40350 42254 40402
rect 42306 40350 42420 40402
rect 42140 40348 42420 40350
rect 42252 40338 42308 40348
rect 42028 40290 42084 40302
rect 42028 40238 42030 40290
rect 42082 40238 42084 40290
rect 41580 40180 41636 40190
rect 41468 39956 41524 39966
rect 41244 39620 41300 39630
rect 41244 39526 41300 39564
rect 39788 37214 39790 37266
rect 39842 37214 39844 37266
rect 39788 37202 39844 37214
rect 40348 36596 40404 36606
rect 40348 36502 40404 36540
rect 39676 35700 39732 36428
rect 40684 36148 40740 39452
rect 41468 38668 41524 39900
rect 41580 39058 41636 40124
rect 41916 39732 41972 39742
rect 41580 39006 41582 39058
rect 41634 39006 41636 39058
rect 41580 38994 41636 39006
rect 41692 39618 41748 39630
rect 41692 39566 41694 39618
rect 41746 39566 41748 39618
rect 41580 38836 41636 38874
rect 41580 38770 41636 38780
rect 41468 38612 41636 38668
rect 40908 37156 40964 37166
rect 40908 37062 40964 37100
rect 40684 36082 40740 36092
rect 39788 35700 39844 35710
rect 40236 35700 40292 35710
rect 39676 35698 40292 35700
rect 39676 35646 39790 35698
rect 39842 35646 40238 35698
rect 40290 35646 40292 35698
rect 39676 35644 40292 35646
rect 39788 35634 39844 35644
rect 40236 35634 40292 35644
rect 39788 35476 39844 35486
rect 40236 35476 40292 35486
rect 39788 35474 40068 35476
rect 39788 35422 39790 35474
rect 39842 35422 40068 35474
rect 39788 35420 40068 35422
rect 39788 35410 39844 35420
rect 40012 35026 40068 35420
rect 40012 34974 40014 35026
rect 40066 34974 40068 35026
rect 40012 34962 40068 34974
rect 39340 34914 39620 34916
rect 39340 34862 39342 34914
rect 39394 34862 39620 34914
rect 39340 34860 39620 34862
rect 39340 34850 39396 34860
rect 38780 34132 38836 34142
rect 38780 34038 38836 34076
rect 38220 33854 38222 33906
rect 38274 33854 38276 33906
rect 38220 33842 38276 33854
rect 39564 33124 39620 34860
rect 39900 34132 39956 34142
rect 39900 33458 39956 34076
rect 39900 33406 39902 33458
rect 39954 33406 39956 33458
rect 39900 33394 39956 33406
rect 39676 33124 39732 33134
rect 39564 33068 39676 33124
rect 39676 33058 39732 33068
rect 37996 32172 38388 32228
rect 37548 32004 37604 32014
rect 38108 32004 38164 32014
rect 37436 32002 38164 32004
rect 37436 31950 37550 32002
rect 37602 31950 38110 32002
rect 38162 31950 38164 32002
rect 37436 31948 38164 31950
rect 37324 31892 37380 31902
rect 37324 31778 37380 31836
rect 37324 31726 37326 31778
rect 37378 31726 37380 31778
rect 37324 31714 37380 31726
rect 36988 31668 37044 31678
rect 36988 31574 37044 31612
rect 37100 31554 37156 31566
rect 37100 31502 37102 31554
rect 37154 31502 37156 31554
rect 37100 31106 37156 31502
rect 37100 31054 37102 31106
rect 37154 31054 37156 31106
rect 37100 31042 37156 31054
rect 37436 30210 37492 31948
rect 37548 31938 37604 31948
rect 38108 31938 38164 31948
rect 37548 31780 37604 31790
rect 37548 31686 37604 31724
rect 38220 31668 38276 31678
rect 38220 31574 38276 31612
rect 37436 30158 37438 30210
rect 37490 30158 37492 30210
rect 37436 30146 37492 30158
rect 38220 30212 38276 30222
rect 38220 30118 38276 30156
rect 37660 30100 37716 30110
rect 37660 30098 37828 30100
rect 37660 30046 37662 30098
rect 37714 30046 37828 30098
rect 37660 30044 37828 30046
rect 37660 30034 37716 30044
rect 36988 29092 37044 29102
rect 36988 27076 37044 29036
rect 37660 29092 37716 29102
rect 37660 28754 37716 29036
rect 37660 28702 37662 28754
rect 37714 28702 37716 28754
rect 37660 28690 37716 28702
rect 37212 28644 37268 28654
rect 37212 27748 37268 28588
rect 36988 26514 37044 27020
rect 36988 26462 36990 26514
rect 37042 26462 37044 26514
rect 36988 26450 37044 26462
rect 37100 27692 37268 27748
rect 37324 27860 37380 27870
rect 37100 26292 37156 27692
rect 37324 27186 37380 27804
rect 37772 27300 37828 30044
rect 38108 29876 38164 29886
rect 38108 28754 38164 29820
rect 38108 28702 38110 28754
rect 38162 28702 38164 28754
rect 38108 28644 38164 28702
rect 38108 28578 38164 28588
rect 37772 27234 37828 27244
rect 37324 27134 37326 27186
rect 37378 27134 37380 27186
rect 37324 27122 37380 27134
rect 38332 27188 38388 32172
rect 38668 31892 38724 31902
rect 38668 31556 38724 31836
rect 39900 31892 39956 31902
rect 39228 31668 39284 31678
rect 38668 31554 38836 31556
rect 38668 31502 38670 31554
rect 38722 31502 38836 31554
rect 38668 31500 38836 31502
rect 38668 31490 38724 31500
rect 38668 30212 38724 30222
rect 38444 30210 38724 30212
rect 38444 30158 38670 30210
rect 38722 30158 38724 30210
rect 38444 30156 38724 30158
rect 38444 27970 38500 30156
rect 38668 30146 38724 30156
rect 38556 28754 38612 28766
rect 38556 28702 38558 28754
rect 38610 28702 38612 28754
rect 38556 28084 38612 28702
rect 38556 28018 38612 28028
rect 38444 27918 38446 27970
rect 38498 27918 38500 27970
rect 38444 27906 38500 27918
rect 38556 27860 38612 27870
rect 38556 27766 38612 27804
rect 38780 27412 38836 31500
rect 39228 30882 39284 31612
rect 39676 31666 39732 31678
rect 39676 31614 39678 31666
rect 39730 31614 39732 31666
rect 39228 30830 39230 30882
rect 39282 30830 39284 30882
rect 39228 30818 39284 30830
rect 39340 31554 39396 31566
rect 39340 31502 39342 31554
rect 39394 31502 39396 31554
rect 39004 30436 39060 30446
rect 39004 30342 39060 30380
rect 39228 30210 39284 30222
rect 39228 30158 39230 30210
rect 39282 30158 39284 30210
rect 39228 29876 39284 30158
rect 39228 29810 39284 29820
rect 39340 28644 39396 31502
rect 39676 31556 39732 31614
rect 39676 31490 39732 31500
rect 39900 31108 39956 31836
rect 40124 31780 40180 31790
rect 39900 31014 39956 31052
rect 40012 31666 40068 31678
rect 40012 31614 40014 31666
rect 40066 31614 40068 31666
rect 40012 31218 40068 31614
rect 40012 31166 40014 31218
rect 40066 31166 40068 31218
rect 40012 30772 40068 31166
rect 40124 31106 40180 31724
rect 40124 31054 40126 31106
rect 40178 31054 40180 31106
rect 40124 31042 40180 31054
rect 39788 30716 40068 30772
rect 40236 30772 40292 35420
rect 41020 35252 41076 35262
rect 41020 34242 41076 35196
rect 41020 34190 41022 34242
rect 41074 34190 41076 34242
rect 41020 34178 41076 34190
rect 40908 34132 40964 34142
rect 40908 34038 40964 34076
rect 41580 33236 41636 38612
rect 41692 37156 41748 39566
rect 41916 38946 41972 39676
rect 41916 38894 41918 38946
rect 41970 38894 41972 38946
rect 41916 38882 41972 38894
rect 42028 38836 42084 40238
rect 42028 38770 42084 38780
rect 42140 38948 42196 38958
rect 42140 38668 42196 38892
rect 42364 38724 42420 40348
rect 42588 40402 42644 40414
rect 42588 40350 42590 40402
rect 42642 40350 42644 40402
rect 42476 40290 42532 40302
rect 42476 40238 42478 40290
rect 42530 40238 42532 40290
rect 42476 39730 42532 40238
rect 42476 39678 42478 39730
rect 42530 39678 42532 39730
rect 42476 39666 42532 39678
rect 42588 39732 42644 40350
rect 42700 40180 42756 42140
rect 43036 41972 43092 41982
rect 43036 41298 43092 41916
rect 43036 41246 43038 41298
rect 43090 41246 43092 41298
rect 43036 41234 43092 41246
rect 43260 41970 43316 43484
rect 44380 42420 44436 42430
rect 43260 41918 43262 41970
rect 43314 41918 43316 41970
rect 42812 41186 42868 41198
rect 42812 41134 42814 41186
rect 42866 41134 42868 41186
rect 42812 40292 42868 41134
rect 43260 40964 43316 41918
rect 44044 41972 44100 41982
rect 44044 41878 44100 41916
rect 43372 41188 43428 41198
rect 43428 41132 43652 41188
rect 43372 41122 43428 41132
rect 43260 40908 43428 40964
rect 42924 40404 42980 40414
rect 43260 40404 43316 40414
rect 42924 40402 43316 40404
rect 42924 40350 42926 40402
rect 42978 40350 43262 40402
rect 43314 40350 43316 40402
rect 42924 40348 43316 40350
rect 42924 40338 42980 40348
rect 43260 40338 43316 40348
rect 42812 40226 42868 40236
rect 42700 40114 42756 40124
rect 43260 40068 43316 40078
rect 43372 40068 43428 40908
rect 43316 40012 43428 40068
rect 43596 40402 43652 41132
rect 43820 41186 43876 41198
rect 43820 41134 43822 41186
rect 43874 41134 43876 41186
rect 43708 40964 43764 40974
rect 43708 40870 43764 40908
rect 43596 40350 43598 40402
rect 43650 40350 43652 40402
rect 43260 40002 43316 40012
rect 42588 38834 42644 39676
rect 42588 38782 42590 38834
rect 42642 38782 42644 38834
rect 42588 38770 42644 38782
rect 42700 39618 42756 39630
rect 42700 39566 42702 39618
rect 42754 39566 42756 39618
rect 42700 38836 42756 39566
rect 42700 38770 42756 38780
rect 43372 38834 43428 38846
rect 43372 38782 43374 38834
rect 43426 38782 43428 38834
rect 42476 38724 42532 38734
rect 42364 38722 42532 38724
rect 42364 38670 42478 38722
rect 42530 38670 42532 38722
rect 42364 38668 42532 38670
rect 42140 38612 42308 38668
rect 42476 38658 42532 38668
rect 43372 38724 43428 38782
rect 43372 38658 43428 38668
rect 43596 38668 43652 40350
rect 43820 40516 43876 41134
rect 44268 41076 44324 41086
rect 44268 40982 44324 41020
rect 44156 40964 44212 40974
rect 44156 40870 44212 40908
rect 44380 40740 44436 42364
rect 44380 40626 44436 40684
rect 44380 40574 44382 40626
rect 44434 40574 44436 40626
rect 44380 40562 44436 40574
rect 43820 40402 43876 40460
rect 43820 40350 43822 40402
rect 43874 40350 43876 40402
rect 43820 40338 43876 40350
rect 44044 40292 44100 40302
rect 43708 39396 43764 39406
rect 43708 39302 43764 39340
rect 43932 38834 43988 38846
rect 43932 38782 43934 38834
rect 43986 38782 43988 38834
rect 43932 38724 43988 38782
rect 43596 38612 43764 38668
rect 43932 38658 43988 38668
rect 41692 37090 41748 37100
rect 42140 35252 42196 35262
rect 42140 35026 42196 35196
rect 42140 34974 42142 35026
rect 42194 34974 42196 35026
rect 42140 34962 42196 34974
rect 42028 34132 42084 34142
rect 42028 34038 42084 34076
rect 41692 34018 41748 34030
rect 41692 33966 41694 34018
rect 41746 33966 41748 34018
rect 41692 33684 41748 33966
rect 41692 33618 41748 33628
rect 42252 33460 42308 38612
rect 43708 38052 43764 38612
rect 44044 38164 44100 40236
rect 44268 39508 44324 39518
rect 44268 39414 44324 39452
rect 44156 38722 44212 38734
rect 44156 38670 44158 38722
rect 44210 38670 44212 38722
rect 44156 38612 44212 38670
rect 44156 38546 44212 38556
rect 44044 38108 44324 38164
rect 43708 38050 44100 38052
rect 43708 37998 43710 38050
rect 43762 37998 44100 38050
rect 43708 37996 44100 37998
rect 42476 37938 42532 37950
rect 42476 37886 42478 37938
rect 42530 37886 42532 37938
rect 42476 37156 42532 37886
rect 42812 37940 42868 37950
rect 42812 37846 42868 37884
rect 43708 37940 43764 37996
rect 43708 37874 43764 37884
rect 43484 37826 43540 37838
rect 43484 37774 43486 37826
rect 43538 37774 43540 37826
rect 43484 37492 43540 37774
rect 43484 37426 43540 37436
rect 43820 37826 43876 37838
rect 43820 37774 43822 37826
rect 43874 37774 43876 37826
rect 43820 37492 43876 37774
rect 43820 37426 43876 37436
rect 43932 37380 43988 37390
rect 43820 37268 43876 37278
rect 43932 37268 43988 37324
rect 43148 37266 43988 37268
rect 43148 37214 43822 37266
rect 43874 37214 43988 37266
rect 43148 37212 43988 37214
rect 42476 37090 42532 37100
rect 43036 37154 43092 37166
rect 43036 37102 43038 37154
rect 43090 37102 43092 37154
rect 42476 36708 42532 36718
rect 43036 36708 43092 37102
rect 42476 36594 42532 36652
rect 42476 36542 42478 36594
rect 42530 36542 42532 36594
rect 42476 36530 42532 36542
rect 42812 36652 43092 36708
rect 42812 36148 42868 36652
rect 42924 36260 42980 36270
rect 43148 36260 43204 37212
rect 43820 37202 43876 37212
rect 43484 37044 43540 37054
rect 42924 36258 43204 36260
rect 42924 36206 42926 36258
rect 42978 36206 43204 36258
rect 42924 36204 43204 36206
rect 42924 36194 42980 36204
rect 42812 36082 42868 36092
rect 42588 34692 42644 34702
rect 43148 34692 43204 36204
rect 42588 34690 43204 34692
rect 42588 34638 42590 34690
rect 42642 34638 43204 34690
rect 42588 34636 43204 34638
rect 42588 34626 42644 34636
rect 42588 34242 42644 34254
rect 42588 34190 42590 34242
rect 42642 34190 42644 34242
rect 42588 34132 42644 34190
rect 42588 34066 42644 34076
rect 43148 34130 43204 34636
rect 43372 36932 43428 36942
rect 43372 34468 43428 36876
rect 43484 36484 43540 36988
rect 43932 36932 43988 36942
rect 43932 36484 43988 36876
rect 43484 35922 43540 36428
rect 43820 36482 43988 36484
rect 43820 36430 43934 36482
rect 43986 36430 43988 36482
rect 43820 36428 43988 36430
rect 43484 35870 43486 35922
rect 43538 35870 43540 35922
rect 43484 35858 43540 35870
rect 43596 36258 43652 36270
rect 43596 36206 43598 36258
rect 43650 36206 43652 36258
rect 43484 34692 43540 34702
rect 43596 34692 43652 36206
rect 43820 35922 43876 36428
rect 43932 36418 43988 36428
rect 43820 35870 43822 35922
rect 43874 35870 43876 35922
rect 43820 35858 43876 35870
rect 43484 34690 43652 34692
rect 43484 34638 43486 34690
rect 43538 34638 43652 34690
rect 43484 34636 43652 34638
rect 43484 34626 43540 34636
rect 43372 34412 43540 34468
rect 43148 34078 43150 34130
rect 43202 34078 43204 34130
rect 43148 34066 43204 34078
rect 42028 33458 42308 33460
rect 42028 33406 42254 33458
rect 42306 33406 42308 33458
rect 42028 33404 42308 33406
rect 41580 33180 41860 33236
rect 40348 33124 40404 33134
rect 40348 31892 40404 33068
rect 41804 32562 41860 33180
rect 41804 32510 41806 32562
rect 41858 32510 41860 32562
rect 41580 32450 41636 32462
rect 41580 32398 41582 32450
rect 41634 32398 41636 32450
rect 41468 32228 41524 32238
rect 41356 32172 41468 32228
rect 40404 31836 40516 31892
rect 40348 31826 40404 31836
rect 39788 30210 39844 30716
rect 40236 30706 40292 30716
rect 40348 31556 40404 31566
rect 40348 30548 40404 31500
rect 39788 30158 39790 30210
rect 39842 30158 39844 30210
rect 39788 30146 39844 30158
rect 40124 30492 40404 30548
rect 39900 29540 39956 29550
rect 39900 29446 39956 29484
rect 40124 29426 40180 30492
rect 40460 30436 40516 31836
rect 40908 31556 40964 31566
rect 40908 31218 40964 31500
rect 40908 31166 40910 31218
rect 40962 31166 40964 31218
rect 40908 31154 40964 31166
rect 41356 30884 41412 32172
rect 41468 32162 41524 32172
rect 41468 31892 41524 31902
rect 41468 31778 41524 31836
rect 41468 31726 41470 31778
rect 41522 31726 41524 31778
rect 41468 31714 41524 31726
rect 41580 31108 41636 32398
rect 41804 31780 41860 32510
rect 41804 31714 41860 31724
rect 41916 31892 41972 31902
rect 41804 31556 41860 31566
rect 41804 31218 41860 31500
rect 41804 31166 41806 31218
rect 41858 31166 41860 31218
rect 41804 31154 41860 31166
rect 41580 31042 41636 31052
rect 41244 30882 41412 30884
rect 41244 30830 41358 30882
rect 41410 30830 41412 30882
rect 41244 30828 41412 30830
rect 41020 30772 41076 30782
rect 40348 30380 40516 30436
rect 40572 30660 40628 30670
rect 40236 30212 40292 30222
rect 40348 30212 40404 30380
rect 40572 30212 40628 30604
rect 40236 30210 40404 30212
rect 40236 30158 40238 30210
rect 40290 30158 40404 30210
rect 40236 30156 40404 30158
rect 40460 30156 40628 30212
rect 40236 30146 40292 30156
rect 40124 29374 40126 29426
rect 40178 29374 40180 29426
rect 40124 29362 40180 29374
rect 39340 28578 39396 28588
rect 40460 28420 40516 30156
rect 40572 29986 40628 29998
rect 40572 29934 40574 29986
rect 40626 29934 40628 29986
rect 40572 28644 40628 29934
rect 40572 28578 40628 28588
rect 41020 29650 41076 30716
rect 41020 29598 41022 29650
rect 41074 29598 41076 29650
rect 40684 28532 40740 28542
rect 40684 28530 40964 28532
rect 40684 28478 40686 28530
rect 40738 28478 40964 28530
rect 40684 28476 40964 28478
rect 40684 28466 40740 28476
rect 40460 28364 40628 28420
rect 40348 28084 40404 28094
rect 39676 27970 39732 27982
rect 39676 27918 39678 27970
rect 39730 27918 39732 27970
rect 38892 27412 38948 27422
rect 38780 27356 38892 27412
rect 38892 27346 38948 27356
rect 38332 27074 38388 27132
rect 39564 27300 39620 27310
rect 38332 27022 38334 27074
rect 38386 27022 38388 27074
rect 38332 27010 38388 27022
rect 38780 27076 38836 27086
rect 39228 27076 39284 27086
rect 38780 27074 39284 27076
rect 38780 27022 38782 27074
rect 38834 27022 39230 27074
rect 39282 27022 39284 27074
rect 38780 27020 39284 27022
rect 38780 27010 38836 27020
rect 39228 27010 39284 27020
rect 37212 26964 37268 26974
rect 37212 26850 37268 26908
rect 37212 26798 37214 26850
rect 37266 26798 37268 26850
rect 37212 26786 37268 26798
rect 37436 26964 37492 26974
rect 37100 26226 37156 26236
rect 37212 26180 37268 26190
rect 37212 26086 37268 26124
rect 37100 25506 37156 25518
rect 37100 25454 37102 25506
rect 37154 25454 37156 25506
rect 36988 25172 37044 25182
rect 36988 24946 37044 25116
rect 36988 24894 36990 24946
rect 37042 24894 37044 24946
rect 36988 24882 37044 24894
rect 36652 24098 36708 24108
rect 36540 23884 36708 23940
rect 36428 23266 36484 23548
rect 36428 23214 36430 23266
rect 36482 23214 36484 23266
rect 36428 23202 36484 23214
rect 36540 23268 36596 23278
rect 36540 23154 36596 23212
rect 36540 23102 36542 23154
rect 36594 23102 36596 23154
rect 36540 23090 36596 23102
rect 36652 23156 36708 23884
rect 36652 23090 36708 23100
rect 37100 23828 37156 25454
rect 37436 24834 37492 26908
rect 38668 26852 38724 26862
rect 38668 26758 38724 26796
rect 38892 26852 38948 26862
rect 38892 26758 38948 26796
rect 39340 26850 39396 26862
rect 39340 26798 39342 26850
rect 39394 26798 39396 26850
rect 39340 26402 39396 26798
rect 39340 26350 39342 26402
rect 39394 26350 39396 26402
rect 39340 26338 39396 26350
rect 39452 26850 39508 26862
rect 39452 26798 39454 26850
rect 39506 26798 39508 26850
rect 37996 25506 38052 25518
rect 37996 25454 37998 25506
rect 38050 25454 38052 25506
rect 37436 24782 37438 24834
rect 37490 24782 37492 24834
rect 37324 24052 37380 24062
rect 37324 23958 37380 23996
rect 36092 22542 36094 22594
rect 36146 22542 36148 22594
rect 36092 22530 36148 22542
rect 36204 22596 36260 22606
rect 36204 22482 36260 22540
rect 36204 22430 36206 22482
rect 36258 22430 36260 22482
rect 36204 22418 36260 22430
rect 36428 22596 36484 22606
rect 36428 22370 36484 22540
rect 37100 22482 37156 23772
rect 37212 23940 37268 23950
rect 37212 23268 37268 23884
rect 37436 23826 37492 24782
rect 37436 23774 37438 23826
rect 37490 23774 37492 23826
rect 37436 23762 37492 23774
rect 37772 25394 37828 25406
rect 37772 25342 37774 25394
rect 37826 25342 37828 25394
rect 37212 23202 37268 23212
rect 37772 23380 37828 25342
rect 37884 25172 37940 25182
rect 37884 23938 37940 25116
rect 37996 24724 38052 25454
rect 38220 25506 38276 25518
rect 38220 25454 38222 25506
rect 38274 25454 38276 25506
rect 38220 24836 38276 25454
rect 38220 24770 38276 24780
rect 38556 24836 38612 24846
rect 37996 24658 38052 24668
rect 37884 23886 37886 23938
rect 37938 23886 37940 23938
rect 37884 23874 37940 23886
rect 38332 23940 38388 23950
rect 38332 23846 38388 23884
rect 37772 23154 37828 23324
rect 38444 23716 38500 23726
rect 38444 23268 38500 23660
rect 38556 23380 38612 24780
rect 38892 24836 38948 24846
rect 38892 24742 38948 24780
rect 38556 23286 38612 23324
rect 38668 24612 38724 24622
rect 39452 24612 39508 26798
rect 39564 25730 39620 27244
rect 39564 25678 39566 25730
rect 39618 25678 39620 25730
rect 39564 25666 39620 25678
rect 38668 23492 38724 24556
rect 38332 23212 38500 23268
rect 38668 23268 38724 23436
rect 38892 24556 39508 24612
rect 38780 23268 38836 23278
rect 38668 23266 38836 23268
rect 38668 23214 38782 23266
rect 38834 23214 38836 23266
rect 38668 23212 38836 23214
rect 37772 23102 37774 23154
rect 37826 23102 37828 23154
rect 37772 23090 37828 23102
rect 38220 23156 38276 23166
rect 37436 22596 37492 22606
rect 37100 22430 37102 22482
rect 37154 22430 37156 22482
rect 37100 22418 37156 22430
rect 37324 22484 37380 22494
rect 37324 22390 37380 22428
rect 36428 22318 36430 22370
rect 36482 22318 36484 22370
rect 36428 22306 36484 22318
rect 35980 22204 36260 22260
rect 36204 21924 36260 22204
rect 36988 21924 37044 21934
rect 36204 21868 36708 21924
rect 35532 21810 35924 21812
rect 35532 21758 35534 21810
rect 35586 21758 35924 21810
rect 35532 21756 35924 21758
rect 35532 21746 35588 21756
rect 33740 21698 33796 21710
rect 33740 21646 33742 21698
rect 33794 21646 33796 21698
rect 33740 21588 33796 21646
rect 33740 21522 33796 21532
rect 34076 21698 34132 21710
rect 34076 21646 34078 21698
rect 34130 21646 34132 21698
rect 33516 21364 33572 21374
rect 33572 21308 34020 21364
rect 33516 21270 33572 21308
rect 33964 20914 34020 21308
rect 33964 20862 33966 20914
rect 34018 20862 34020 20914
rect 33964 20850 34020 20862
rect 34076 20244 34132 21646
rect 34748 21700 34804 21710
rect 34748 21698 35028 21700
rect 34748 21646 34750 21698
rect 34802 21646 35028 21698
rect 34748 21644 35028 21646
rect 34748 21634 34804 21644
rect 33292 18498 33348 18508
rect 33404 20018 33460 20030
rect 33404 19966 33406 20018
rect 33458 19966 33460 20018
rect 33180 18340 33236 18350
rect 33404 18340 33460 19966
rect 33180 18338 33460 18340
rect 33180 18286 33182 18338
rect 33234 18286 33460 18338
rect 33180 18284 33460 18286
rect 33516 19348 33572 19358
rect 33180 18274 33236 18284
rect 32396 16942 32398 16994
rect 32450 16942 32452 16994
rect 32396 16930 32452 16942
rect 32732 18228 32788 18238
rect 31948 16818 32004 16828
rect 31612 16660 31668 16670
rect 31612 16566 31668 16604
rect 30828 16370 30884 16380
rect 30828 16212 30884 16222
rect 30828 16118 30884 16156
rect 31836 16212 31892 16222
rect 30940 15540 30996 15550
rect 30716 15538 30996 15540
rect 30716 15486 30942 15538
rect 30994 15486 30996 15538
rect 30716 15484 30996 15486
rect 30940 15474 30996 15484
rect 31500 15426 31556 15438
rect 31500 15374 31502 15426
rect 31554 15374 31556 15426
rect 29820 15092 29988 15148
rect 31276 15316 31332 15326
rect 31276 15202 31332 15260
rect 31276 15150 31278 15202
rect 31330 15150 31332 15202
rect 31276 15138 31332 15150
rect 29148 14812 29316 14868
rect 29148 12852 29204 12862
rect 28588 9266 28756 9268
rect 28588 9214 28590 9266
rect 28642 9214 28756 9266
rect 28588 9212 28756 9214
rect 28812 12850 29204 12852
rect 28812 12798 29150 12850
rect 29202 12798 29204 12850
rect 28812 12796 29204 12798
rect 28588 9202 28644 9212
rect 27580 9156 27636 9166
rect 27580 9062 27636 9100
rect 27804 9044 27860 9054
rect 27804 8950 27860 8988
rect 28476 8930 28532 8942
rect 28476 8878 28478 8930
rect 28530 8878 28532 8930
rect 27356 7534 27358 7586
rect 27410 7534 27412 7586
rect 27356 7522 27412 7534
rect 27916 8372 27972 8382
rect 28476 8372 28532 8878
rect 28588 8372 28644 8382
rect 28476 8316 28588 8372
rect 27916 7586 27972 8316
rect 28588 8278 28644 8316
rect 28812 8036 28868 12796
rect 29148 12786 29204 12796
rect 29260 12404 29316 14812
rect 29596 13634 29652 13646
rect 29596 13582 29598 13634
rect 29650 13582 29652 13634
rect 29596 13524 29652 13582
rect 29596 13458 29652 13468
rect 29372 12964 29428 12974
rect 29372 12870 29428 12908
rect 29596 12962 29652 12974
rect 29596 12910 29598 12962
rect 29650 12910 29652 12962
rect 29596 12516 29652 12910
rect 29708 12964 29764 12974
rect 29708 12870 29764 12908
rect 29596 12460 29764 12516
rect 29148 12402 29652 12404
rect 29148 12350 29262 12402
rect 29314 12350 29652 12402
rect 29148 12348 29652 12350
rect 29148 9268 29204 12348
rect 29260 12338 29316 12348
rect 29596 12290 29652 12348
rect 29596 12238 29598 12290
rect 29650 12238 29652 12290
rect 29596 12226 29652 12238
rect 29596 11956 29652 11966
rect 29596 11394 29652 11900
rect 29596 11342 29598 11394
rect 29650 11342 29652 11394
rect 29596 11330 29652 11342
rect 29148 9202 29204 9212
rect 29260 11284 29316 11294
rect 29260 8930 29316 11228
rect 29372 11172 29428 11182
rect 29708 11172 29764 12460
rect 29372 11170 29764 11172
rect 29372 11118 29374 11170
rect 29426 11118 29764 11170
rect 29372 11116 29764 11118
rect 29372 11106 29428 11116
rect 29596 10836 29652 10846
rect 29820 10836 29876 15092
rect 31500 14756 31556 15374
rect 31836 15426 31892 16156
rect 32732 16100 32788 18172
rect 33516 18226 33572 19292
rect 33740 19012 33796 19022
rect 33740 18562 33796 18956
rect 33740 18510 33742 18562
rect 33794 18510 33796 18562
rect 33740 18498 33796 18510
rect 34076 18562 34132 20188
rect 34972 20130 35028 21644
rect 35084 21586 35140 21598
rect 35084 21534 35086 21586
rect 35138 21534 35140 21586
rect 35084 21026 35140 21534
rect 35644 21588 35700 21598
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20974 35086 21026
rect 35138 20974 35140 21026
rect 35084 20962 35140 20974
rect 34972 20078 34974 20130
rect 35026 20078 35028 20130
rect 34972 20066 35028 20078
rect 35420 20802 35476 20814
rect 35420 20750 35422 20802
rect 35474 20750 35476 20802
rect 34076 18510 34078 18562
rect 34130 18510 34132 18562
rect 34076 18498 34132 18510
rect 34300 20018 34356 20030
rect 34300 19966 34302 20018
rect 34354 19966 34356 20018
rect 33516 18174 33518 18226
rect 33570 18174 33572 18226
rect 32956 16436 33012 16446
rect 32956 16210 33012 16380
rect 32956 16158 32958 16210
rect 33010 16158 33012 16210
rect 32956 16146 33012 16158
rect 32732 16034 32788 16044
rect 31836 15374 31838 15426
rect 31890 15374 31892 15426
rect 31836 15362 31892 15374
rect 32508 15540 32564 15550
rect 30380 14530 30436 14542
rect 30380 14478 30382 14530
rect 30434 14478 30436 14530
rect 29932 13636 29988 13646
rect 29932 12738 29988 13580
rect 30380 13186 30436 14478
rect 30604 14308 30660 14318
rect 30604 14214 30660 14252
rect 30380 13134 30382 13186
rect 30434 13134 30436 13186
rect 30380 13122 30436 13134
rect 31276 13524 31332 13534
rect 29932 12686 29934 12738
rect 29986 12686 29988 12738
rect 29932 12674 29988 12686
rect 30716 12962 30772 12974
rect 30716 12910 30718 12962
rect 30770 12910 30772 12962
rect 29932 12404 29988 12414
rect 29932 12310 29988 12348
rect 30716 12404 30772 12910
rect 31276 12850 31332 13468
rect 31500 12962 31556 14700
rect 31612 14308 31668 14318
rect 31668 14252 31780 14308
rect 31612 14242 31668 14252
rect 31724 13858 31780 14252
rect 31724 13806 31726 13858
rect 31778 13806 31780 13858
rect 31724 13794 31780 13806
rect 32508 13748 32564 15484
rect 33404 15540 33460 15550
rect 33404 15446 33460 15484
rect 33180 13748 33236 13758
rect 32508 13746 32788 13748
rect 32508 13694 32510 13746
rect 32562 13694 32788 13746
rect 32508 13692 32788 13694
rect 32508 13682 32564 13692
rect 32732 13076 32788 13692
rect 33180 13654 33236 13692
rect 33516 13746 33572 18174
rect 33628 18340 33684 18350
rect 33628 16882 33684 18284
rect 34300 18340 34356 19966
rect 35420 19908 35476 20750
rect 35644 20690 35700 21532
rect 35868 21586 35924 21756
rect 36652 21698 36708 21868
rect 36652 21646 36654 21698
rect 36706 21646 36708 21698
rect 36652 21634 36708 21646
rect 35868 21534 35870 21586
rect 35922 21534 35924 21586
rect 35868 21522 35924 21534
rect 35644 20638 35646 20690
rect 35698 20638 35700 20690
rect 35644 20626 35700 20638
rect 35980 20690 36036 20702
rect 35980 20638 35982 20690
rect 36034 20638 36036 20690
rect 35980 20468 36036 20638
rect 35420 19796 35476 19852
rect 35084 19740 35476 19796
rect 35532 20412 36036 20468
rect 35532 20356 35588 20412
rect 34636 19348 34692 19358
rect 34636 19254 34692 19292
rect 34300 18274 34356 18284
rect 34860 18340 34916 18350
rect 34860 18246 34916 18284
rect 35084 18116 35140 19740
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35308 19234 35364 19246
rect 35308 19182 35310 19234
rect 35362 19182 35364 19234
rect 35308 19012 35364 19182
rect 35420 19124 35476 19134
rect 35532 19124 35588 20300
rect 36988 20132 37044 21868
rect 37212 20916 37268 20926
rect 37436 20916 37492 22540
rect 38220 22594 38276 23100
rect 38220 22542 38222 22594
rect 38274 22542 38276 22594
rect 38220 22530 38276 22542
rect 38332 22594 38388 23212
rect 38780 23202 38836 23212
rect 38892 22932 38948 24556
rect 39116 24388 39172 24398
rect 39004 23604 39060 23614
rect 39004 23154 39060 23548
rect 39004 23102 39006 23154
rect 39058 23102 39060 23154
rect 39004 23090 39060 23102
rect 38668 22876 38948 22932
rect 38332 22542 38334 22594
rect 38386 22542 38388 22594
rect 38332 22530 38388 22542
rect 38556 22596 38612 22606
rect 38556 22502 38612 22540
rect 38668 22594 38724 22876
rect 38668 22542 38670 22594
rect 38722 22542 38724 22594
rect 38668 22530 38724 22542
rect 39116 22596 39172 24332
rect 39676 23828 39732 27918
rect 40012 27412 40068 27422
rect 40012 27186 40068 27356
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 40012 27076 40068 27134
rect 40012 27010 40068 27020
rect 40348 27076 40404 28028
rect 40460 27188 40516 27198
rect 40460 27094 40516 27132
rect 40124 26292 40180 26302
rect 40124 26198 40180 26236
rect 39900 26180 39956 26190
rect 39900 25508 39956 26124
rect 40124 25620 40180 25630
rect 40348 25620 40404 27020
rect 40180 25564 40404 25620
rect 40124 25526 40180 25564
rect 39900 25414 39956 25452
rect 40012 25506 40068 25518
rect 40012 25454 40014 25506
rect 40066 25454 40068 25506
rect 40012 24948 40068 25454
rect 40012 24892 40180 24948
rect 40124 24836 40180 24892
rect 40124 24780 40292 24836
rect 40012 24724 40068 24734
rect 40068 24668 40180 24724
rect 40012 24630 40068 24668
rect 40012 23938 40068 23950
rect 40012 23886 40014 23938
rect 40066 23886 40068 23938
rect 39900 23828 39956 23838
rect 39676 23826 39956 23828
rect 39676 23774 39902 23826
rect 39954 23774 39956 23826
rect 39676 23772 39956 23774
rect 39564 23604 39620 23614
rect 39452 23548 39564 23604
rect 39452 23154 39508 23548
rect 39564 23538 39620 23548
rect 39452 23102 39454 23154
rect 39506 23102 39508 23154
rect 39452 23090 39508 23102
rect 39564 23380 39620 23390
rect 38892 22484 38948 22494
rect 37772 22146 37828 22158
rect 37772 22094 37774 22146
rect 37826 22094 37828 22146
rect 37772 21924 37828 22094
rect 37772 21858 37828 21868
rect 38892 21810 38948 22428
rect 39116 22482 39172 22540
rect 39116 22430 39118 22482
rect 39170 22430 39172 22482
rect 39116 22418 39172 22430
rect 39564 22372 39620 23324
rect 39788 23380 39844 23390
rect 39676 23268 39732 23278
rect 39676 23174 39732 23212
rect 39788 23266 39844 23324
rect 39788 23214 39790 23266
rect 39842 23214 39844 23266
rect 39788 23202 39844 23214
rect 39900 22484 39956 23772
rect 39900 22418 39956 22428
rect 40012 23492 40068 23886
rect 39788 22372 39844 22382
rect 39564 22370 39844 22372
rect 39564 22318 39790 22370
rect 39842 22318 39844 22370
rect 39564 22316 39844 22318
rect 39788 22306 39844 22316
rect 40012 22372 40068 23436
rect 40124 22484 40180 24668
rect 40236 23604 40292 24780
rect 40236 23538 40292 23548
rect 40124 22390 40180 22428
rect 40236 23154 40292 23166
rect 40236 23102 40238 23154
rect 40290 23102 40292 23154
rect 40012 22306 40068 22316
rect 40236 22260 40292 23102
rect 40460 22930 40516 22942
rect 40460 22878 40462 22930
rect 40514 22878 40516 22930
rect 40460 22484 40516 22878
rect 40572 22708 40628 28364
rect 40908 27746 40964 28476
rect 41020 28082 41076 29598
rect 41132 30210 41188 30222
rect 41132 30158 41134 30210
rect 41186 30158 41188 30210
rect 41132 28980 41188 30158
rect 41132 28914 41188 28924
rect 41020 28030 41022 28082
rect 41074 28030 41076 28082
rect 41020 28018 41076 28030
rect 41244 27860 41300 30828
rect 41356 30818 41412 30828
rect 41692 30772 41748 30782
rect 41692 30210 41748 30716
rect 41692 30158 41694 30210
rect 41746 30158 41748 30210
rect 41692 30146 41748 30158
rect 41692 29316 41748 29326
rect 41468 28756 41524 28766
rect 41468 28642 41524 28700
rect 41468 28590 41470 28642
rect 41522 28590 41524 28642
rect 41468 28578 41524 28590
rect 40908 27694 40910 27746
rect 40962 27694 40964 27746
rect 40908 27682 40964 27694
rect 41020 27804 41300 27860
rect 41692 27858 41748 29260
rect 41916 28756 41972 31836
rect 42028 30436 42084 33404
rect 42252 33394 42308 33404
rect 42812 33124 42868 33134
rect 43260 33124 43316 33134
rect 42812 33122 43316 33124
rect 42812 33070 42814 33122
rect 42866 33070 43262 33122
rect 43314 33070 43316 33122
rect 42812 33068 43316 33070
rect 42812 33058 42868 33068
rect 42140 32788 42196 32798
rect 42140 32786 43204 32788
rect 42140 32734 42142 32786
rect 42194 32734 43204 32786
rect 42140 32732 43204 32734
rect 42140 32722 42196 32732
rect 42924 32564 42980 32574
rect 42812 32452 42868 32462
rect 42140 31668 42196 31678
rect 42140 31666 42532 31668
rect 42140 31614 42142 31666
rect 42194 31614 42532 31666
rect 42140 31612 42532 31614
rect 42140 31602 42196 31612
rect 42140 31108 42196 31118
rect 42140 31106 42308 31108
rect 42140 31054 42142 31106
rect 42194 31054 42308 31106
rect 42140 31052 42308 31054
rect 42140 31042 42196 31052
rect 42028 30380 42196 30436
rect 41916 28662 41972 28700
rect 42028 30212 42084 30222
rect 41692 27806 41694 27858
rect 41746 27806 41748 27858
rect 41020 26404 41076 27804
rect 41244 27636 41300 27646
rect 41244 27542 41300 27580
rect 41692 27188 41748 27806
rect 41356 27132 41748 27188
rect 41804 27636 41860 27646
rect 41804 27186 41860 27580
rect 42028 27524 42084 30156
rect 42028 27458 42084 27468
rect 42140 27300 42196 30380
rect 42252 29428 42308 31052
rect 42476 30882 42532 31612
rect 42476 30830 42478 30882
rect 42530 30830 42532 30882
rect 42476 30818 42532 30830
rect 42588 31106 42644 31118
rect 42588 31054 42590 31106
rect 42642 31054 42644 31106
rect 42588 30772 42644 31054
rect 42812 31106 42868 32396
rect 42812 31054 42814 31106
rect 42866 31054 42868 31106
rect 42812 31042 42868 31054
rect 42924 32450 42980 32508
rect 42924 32398 42926 32450
rect 42978 32398 42980 32450
rect 42588 30706 42644 30716
rect 42924 30436 42980 32398
rect 42476 30380 42980 30436
rect 43148 31218 43204 32732
rect 43260 31332 43316 33068
rect 43372 32788 43428 32798
rect 43372 32694 43428 32732
rect 43484 32564 43540 34412
rect 43596 33796 43652 34636
rect 43596 33730 43652 33740
rect 43708 35252 43764 35262
rect 43708 32900 43764 35196
rect 43820 35140 43876 35150
rect 44044 35140 44100 37996
rect 44156 37378 44212 37390
rect 44156 37326 44158 37378
rect 44210 37326 44212 37378
rect 44156 36708 44212 37326
rect 44156 36642 44212 36652
rect 44268 36484 44324 38108
rect 44380 37826 44436 37838
rect 44380 37774 44382 37826
rect 44434 37774 44436 37826
rect 44380 37380 44436 37774
rect 44492 37828 44548 45052
rect 44828 44660 44884 44670
rect 44828 44434 44884 44604
rect 44828 44382 44830 44434
rect 44882 44382 44884 44434
rect 44828 43652 44884 44382
rect 46956 44212 47012 44222
rect 46172 44210 47012 44212
rect 46172 44158 46958 44210
rect 47010 44158 47012 44210
rect 46172 44156 47012 44158
rect 46172 43762 46228 44156
rect 46956 44146 47012 44156
rect 46172 43710 46174 43762
rect 46226 43710 46228 43762
rect 46172 43698 46228 43710
rect 44828 43538 44884 43596
rect 46844 43652 46900 43662
rect 46844 43558 46900 43596
rect 44828 43486 44830 43538
rect 44882 43486 44884 43538
rect 44828 43474 44884 43486
rect 45276 43538 45332 43550
rect 45276 43486 45278 43538
rect 45330 43486 45332 43538
rect 45276 42980 45332 43486
rect 45388 43428 45444 43438
rect 45388 43334 45444 43372
rect 46172 43428 46228 43438
rect 46172 43334 46228 43372
rect 47292 43426 47348 43438
rect 47292 43374 47294 43426
rect 47346 43374 47348 43426
rect 45836 43316 45892 43326
rect 45276 42886 45332 42924
rect 45724 43314 45892 43316
rect 45724 43262 45838 43314
rect 45890 43262 45892 43314
rect 45724 43260 45892 43262
rect 45388 42532 45444 42542
rect 45724 42532 45780 43260
rect 45836 43250 45892 43260
rect 46060 43316 46116 43326
rect 45836 42978 45892 42990
rect 45836 42926 45838 42978
rect 45890 42926 45892 42978
rect 45836 42866 45892 42926
rect 45836 42814 45838 42866
rect 45890 42814 45892 42866
rect 45836 42802 45892 42814
rect 45388 42530 45780 42532
rect 45388 42478 45390 42530
rect 45442 42478 45780 42530
rect 45388 42476 45780 42478
rect 45388 42466 45444 42476
rect 45388 41970 45444 41982
rect 45388 41918 45390 41970
rect 45442 41918 45444 41970
rect 44828 41300 44884 41310
rect 44828 41298 45108 41300
rect 44828 41246 44830 41298
rect 44882 41246 45108 41298
rect 44828 41244 45108 41246
rect 44828 41234 44884 41244
rect 44828 40852 44884 40862
rect 44884 40796 44996 40852
rect 44828 40786 44884 40796
rect 44940 40402 44996 40796
rect 45052 40628 45108 41244
rect 45276 40628 45332 40638
rect 45108 40626 45332 40628
rect 45108 40574 45278 40626
rect 45330 40574 45332 40626
rect 45108 40572 45332 40574
rect 45052 40534 45108 40572
rect 45276 40562 45332 40572
rect 44940 40350 44942 40402
rect 44994 40350 44996 40402
rect 44940 40338 44996 40350
rect 45052 40292 45108 40302
rect 44828 39618 44884 39630
rect 44828 39566 44830 39618
rect 44882 39566 44884 39618
rect 44828 39508 44884 39566
rect 44828 39442 44884 39452
rect 44604 39396 44660 39406
rect 44604 38836 44660 39340
rect 45052 39396 45108 40236
rect 45388 40180 45444 41918
rect 45388 40114 45444 40124
rect 45500 39844 45556 42476
rect 45612 42308 45668 42318
rect 45612 41858 45668 42252
rect 46060 41972 46116 43260
rect 47292 43316 47348 43374
rect 47292 43250 47348 43260
rect 47628 43092 47684 45724
rect 49868 45668 49924 45678
rect 50092 45668 50148 46396
rect 50652 45668 50708 46398
rect 51548 46116 51604 46126
rect 51548 46022 51604 46060
rect 49868 45666 50148 45668
rect 49868 45614 49870 45666
rect 49922 45614 50148 45666
rect 49868 45612 50148 45614
rect 50204 45612 50708 45668
rect 51660 45778 51716 45790
rect 51660 45726 51662 45778
rect 51714 45726 51716 45778
rect 49420 45108 49476 45118
rect 49868 45108 49924 45612
rect 50204 45218 50260 45612
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50204 45166 50206 45218
rect 50258 45166 50260 45218
rect 50204 45154 50260 45166
rect 49420 45106 49924 45108
rect 49420 45054 49422 45106
rect 49474 45054 49924 45106
rect 49420 45052 49924 45054
rect 49084 44996 49140 45006
rect 49420 44996 49476 45052
rect 49084 44994 49476 44996
rect 49084 44942 49086 44994
rect 49138 44942 49476 44994
rect 49084 44940 49476 44942
rect 51660 44996 51716 45726
rect 47740 44322 47796 44334
rect 47740 44270 47742 44322
rect 47794 44270 47796 44322
rect 47740 44100 47796 44270
rect 48188 44100 48244 44110
rect 47740 44044 48188 44100
rect 47292 43036 47684 43092
rect 46620 42868 46676 42878
rect 46284 42756 46340 42766
rect 46284 42662 46340 42700
rect 46620 42642 46676 42812
rect 46620 42590 46622 42642
rect 46674 42590 46676 42642
rect 46620 42084 46676 42590
rect 46844 42754 46900 42766
rect 46844 42702 46846 42754
rect 46898 42702 46900 42754
rect 46844 42644 46900 42702
rect 46844 42578 46900 42588
rect 46620 42018 46676 42028
rect 45612 41806 45614 41858
rect 45666 41806 45668 41858
rect 45612 41794 45668 41806
rect 45836 41916 46116 41972
rect 45612 40514 45668 40526
rect 45612 40462 45614 40514
rect 45666 40462 45668 40514
rect 45612 40292 45668 40462
rect 45836 40404 45892 41916
rect 46060 41748 46116 41758
rect 46060 41654 46116 41692
rect 46956 41076 47012 41086
rect 46060 41074 47012 41076
rect 46060 41022 46958 41074
rect 47010 41022 47012 41074
rect 46060 41020 47012 41022
rect 45948 40740 46004 40750
rect 45948 40626 46004 40684
rect 45948 40574 45950 40626
rect 46002 40574 46004 40626
rect 45948 40562 46004 40574
rect 45836 40348 46004 40404
rect 45612 40226 45668 40236
rect 45052 39330 45108 39340
rect 45164 39788 45556 39844
rect 44604 38742 44660 38780
rect 45052 38834 45108 38846
rect 45052 38782 45054 38834
rect 45106 38782 45108 38834
rect 44828 38612 44884 38622
rect 44716 38052 44772 38062
rect 44828 38052 44884 38556
rect 44716 38050 44884 38052
rect 44716 37998 44718 38050
rect 44770 37998 44884 38050
rect 44716 37996 44884 37998
rect 45052 38164 45108 38782
rect 45164 38724 45220 39788
rect 45388 39620 45444 39630
rect 45388 39526 45444 39564
rect 45612 39508 45668 39518
rect 45276 39396 45332 39406
rect 45276 39302 45332 39340
rect 45500 39396 45556 39434
rect 45500 39330 45556 39340
rect 45500 38948 45556 38958
rect 45612 38948 45668 39452
rect 45836 39508 45892 39518
rect 45836 39414 45892 39452
rect 45948 39172 46004 40348
rect 46060 39394 46116 41020
rect 46956 41010 47012 41020
rect 46844 40740 46900 40750
rect 46844 40628 46900 40684
rect 47180 40628 47236 40638
rect 46844 40626 47236 40628
rect 46844 40574 46846 40626
rect 46898 40574 47182 40626
rect 47234 40574 47236 40626
rect 46844 40572 47236 40574
rect 46844 40562 46900 40572
rect 47180 40562 47236 40572
rect 46284 40514 46340 40526
rect 46284 40462 46286 40514
rect 46338 40462 46340 40514
rect 46284 39956 46340 40462
rect 46284 39890 46340 39900
rect 46956 40292 47012 40302
rect 46284 39620 46340 39630
rect 46284 39526 46340 39564
rect 46172 39508 46228 39518
rect 46172 39414 46228 39452
rect 46844 39506 46900 39518
rect 46844 39454 46846 39506
rect 46898 39454 46900 39506
rect 46060 39342 46062 39394
rect 46114 39342 46116 39394
rect 46060 39330 46116 39342
rect 45948 39116 46564 39172
rect 45500 38946 45668 38948
rect 45500 38894 45502 38946
rect 45554 38894 45668 38946
rect 45500 38892 45668 38894
rect 45948 38948 46004 38958
rect 45500 38882 45556 38892
rect 45948 38854 46004 38892
rect 45724 38724 45780 38734
rect 45164 38668 45444 38724
rect 45388 38612 45556 38668
rect 44716 37986 44772 37996
rect 44940 37938 44996 37950
rect 44940 37886 44942 37938
rect 44994 37886 44996 37938
rect 44492 37762 44548 37772
rect 44828 37828 44884 37838
rect 44380 37314 44436 37324
rect 44828 37266 44884 37772
rect 44828 37214 44830 37266
rect 44882 37214 44884 37266
rect 44828 37202 44884 37214
rect 43820 35138 44100 35140
rect 43820 35086 43822 35138
rect 43874 35086 44100 35138
rect 43820 35084 44100 35086
rect 44156 36428 44324 36484
rect 44828 36484 44884 36494
rect 44940 36484 44996 37886
rect 45052 37268 45108 38108
rect 45164 37940 45220 37950
rect 45164 37846 45220 37884
rect 45388 37940 45444 37950
rect 45388 37846 45444 37884
rect 45500 37604 45556 38612
rect 45724 38050 45780 38668
rect 46396 38724 46452 38762
rect 46396 38658 46452 38668
rect 45836 38274 45892 38286
rect 45836 38222 45838 38274
rect 45890 38222 45892 38274
rect 45836 38164 45892 38222
rect 45836 38098 45892 38108
rect 45724 37998 45726 38050
rect 45778 37998 45780 38050
rect 45724 37986 45780 37998
rect 45388 37548 45556 37604
rect 45612 37940 45668 37950
rect 45052 37212 45220 37268
rect 44828 36482 44996 36484
rect 44828 36430 44830 36482
rect 44882 36430 44996 36482
rect 44828 36428 44996 36430
rect 45164 36482 45220 37212
rect 45276 37156 45332 37166
rect 45276 37062 45332 37100
rect 45164 36430 45166 36482
rect 45218 36430 45220 36482
rect 43820 35074 43876 35084
rect 44156 34914 44212 36428
rect 44828 36418 44884 36428
rect 45164 36418 45220 36430
rect 45276 36484 45332 36494
rect 45388 36484 45444 37548
rect 45500 37044 45556 37054
rect 45612 37044 45668 37884
rect 45836 37940 45892 37950
rect 45836 37846 45892 37884
rect 46396 37940 46452 37950
rect 46396 37846 46452 37884
rect 45556 36988 45668 37044
rect 45724 37492 45780 37502
rect 45724 37378 45780 37436
rect 45724 37326 45726 37378
rect 45778 37326 45780 37378
rect 45500 36978 45556 36988
rect 45332 36428 45444 36484
rect 45500 36484 45556 36494
rect 45500 36482 45668 36484
rect 45500 36430 45502 36482
rect 45554 36430 45668 36482
rect 45500 36428 45668 36430
rect 45276 36390 45332 36428
rect 45500 36418 45556 36428
rect 44268 36258 44324 36270
rect 44268 36206 44270 36258
rect 44322 36206 44324 36258
rect 44268 35700 44324 36206
rect 44940 36260 44996 36270
rect 44268 35634 44324 35644
rect 44716 35700 44772 35710
rect 44716 35606 44772 35644
rect 44940 35698 44996 36204
rect 45164 36258 45220 36270
rect 45164 36206 45166 36258
rect 45218 36206 45220 36258
rect 45164 36148 45220 36206
rect 45164 36082 45220 36092
rect 45500 36260 45556 36270
rect 45612 36260 45668 36428
rect 45724 36482 45780 37326
rect 45836 37268 45892 37278
rect 45836 37174 45892 37212
rect 45724 36430 45726 36482
rect 45778 36430 45780 36482
rect 45724 36418 45780 36430
rect 46060 37044 46116 37054
rect 46060 36482 46116 36988
rect 46060 36430 46062 36482
rect 46114 36430 46116 36482
rect 46060 36418 46116 36430
rect 46172 36932 46228 36942
rect 45612 36204 45892 36260
rect 44940 35646 44942 35698
rect 44994 35646 44996 35698
rect 44940 35634 44996 35646
rect 45164 35924 45220 35934
rect 45164 35698 45220 35868
rect 45500 35922 45556 36204
rect 45500 35870 45502 35922
rect 45554 35870 45556 35922
rect 45500 35858 45556 35870
rect 45164 35646 45166 35698
rect 45218 35646 45220 35698
rect 45164 35634 45220 35646
rect 45724 35700 45780 35710
rect 45724 35606 45780 35644
rect 44380 35586 44436 35598
rect 44380 35534 44382 35586
rect 44434 35534 44436 35586
rect 44380 35252 44436 35534
rect 45612 35586 45668 35598
rect 45612 35534 45614 35586
rect 45666 35534 45668 35586
rect 44604 35476 44660 35486
rect 45612 35476 45668 35534
rect 44380 35186 44436 35196
rect 44492 35474 44660 35476
rect 44492 35422 44606 35474
rect 44658 35422 44660 35474
rect 44492 35420 44660 35422
rect 44156 34862 44158 34914
rect 44210 34862 44212 34914
rect 43932 34692 43988 34702
rect 43932 34598 43988 34636
rect 44156 34468 44212 34862
rect 43932 34412 44212 34468
rect 43820 34244 43876 34254
rect 43820 34150 43876 34188
rect 43932 33572 43988 34412
rect 44492 34356 44548 35420
rect 44604 35410 44660 35420
rect 45164 35420 45668 35476
rect 44716 34916 44772 34926
rect 43932 33506 43988 33516
rect 44044 34300 44548 34356
rect 44604 34914 44772 34916
rect 44604 34862 44718 34914
rect 44770 34862 44772 34914
rect 44604 34860 44772 34862
rect 44044 33570 44100 34300
rect 44604 33684 44660 34860
rect 44716 34850 44772 34860
rect 45164 34914 45220 35420
rect 45836 35364 45892 36204
rect 45948 35924 46004 35934
rect 45948 35830 46004 35868
rect 45612 35308 45892 35364
rect 45276 35252 45332 35262
rect 45276 35138 45332 35196
rect 45276 35086 45278 35138
rect 45330 35086 45332 35138
rect 45276 35074 45332 35086
rect 45164 34862 45166 34914
rect 45218 34862 45220 34914
rect 45164 34850 45220 34862
rect 45500 34916 45556 34926
rect 45612 34916 45668 35308
rect 46172 35028 46228 36876
rect 46396 36820 46452 36830
rect 46508 36820 46564 39116
rect 46844 39060 46900 39454
rect 46956 39506 47012 40236
rect 47292 39844 47348 43036
rect 47404 42756 47460 42766
rect 47404 41188 47460 42700
rect 48188 42756 48244 44044
rect 49084 44100 49140 44940
rect 51660 44930 51716 44940
rect 52332 44996 52388 45006
rect 52332 44902 52388 44940
rect 49084 44034 49140 44044
rect 50876 44098 50932 44110
rect 50876 44046 50878 44098
rect 50930 44046 50932 44098
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50092 43652 50148 43662
rect 50428 43652 50484 43662
rect 49644 43650 50148 43652
rect 49644 43598 50094 43650
rect 50146 43598 50148 43650
rect 49644 43596 50148 43598
rect 49084 43538 49140 43550
rect 49084 43486 49086 43538
rect 49138 43486 49140 43538
rect 48188 42690 48244 42700
rect 48748 43428 48804 43438
rect 48076 42642 48132 42654
rect 48076 42590 48078 42642
rect 48130 42590 48132 42642
rect 47740 41188 47796 41198
rect 47404 41186 47796 41188
rect 47404 41134 47742 41186
rect 47794 41134 47796 41186
rect 47404 41132 47796 41134
rect 48076 41188 48132 42590
rect 48748 41860 48804 43372
rect 49084 42644 49140 43486
rect 49644 43538 49700 43596
rect 49644 43486 49646 43538
rect 49698 43486 49700 43538
rect 49644 43474 49700 43486
rect 49084 42578 49140 42588
rect 49756 43426 49812 43438
rect 49756 43374 49758 43426
rect 49810 43374 49812 43426
rect 49756 42644 49812 43374
rect 50092 42868 50148 43596
rect 50316 43650 50484 43652
rect 50316 43598 50430 43650
rect 50482 43598 50484 43650
rect 50316 43596 50484 43598
rect 50204 42868 50260 42878
rect 50092 42866 50260 42868
rect 50092 42814 50206 42866
rect 50258 42814 50260 42866
rect 50092 42812 50260 42814
rect 50204 42802 50260 42812
rect 49420 41970 49476 41982
rect 49420 41918 49422 41970
rect 49474 41918 49476 41970
rect 48748 41300 48804 41804
rect 48860 41860 48916 41870
rect 48860 41858 49028 41860
rect 48860 41806 48862 41858
rect 48914 41806 49028 41858
rect 48860 41804 49028 41806
rect 48860 41794 48916 41804
rect 48860 41300 48916 41310
rect 48748 41298 48916 41300
rect 48748 41246 48862 41298
rect 48914 41246 48916 41298
rect 48748 41244 48916 41246
rect 48076 41132 48804 41188
rect 47740 40964 47796 41132
rect 48188 40964 48244 40974
rect 47740 40962 48356 40964
rect 47740 40910 48190 40962
rect 48242 40910 48356 40962
rect 47740 40908 48356 40910
rect 48188 40898 48244 40908
rect 48188 40628 48244 40638
rect 48188 40402 48244 40572
rect 48188 40350 48190 40402
rect 48242 40350 48244 40402
rect 47740 40292 47796 40302
rect 47796 40236 48132 40292
rect 47740 40198 47796 40236
rect 47292 39778 47348 39788
rect 47852 39844 47908 39854
rect 47180 39620 47236 39630
rect 47516 39620 47572 39630
rect 47180 39618 47572 39620
rect 47180 39566 47182 39618
rect 47234 39566 47518 39618
rect 47570 39566 47572 39618
rect 47180 39564 47572 39566
rect 47180 39554 47236 39564
rect 47516 39554 47572 39564
rect 46956 39454 46958 39506
rect 47010 39454 47012 39506
rect 46956 39442 47012 39454
rect 47852 39284 47908 39788
rect 47852 39218 47908 39228
rect 47964 39620 48020 39630
rect 46956 39060 47012 39070
rect 46844 39058 47012 39060
rect 46844 39006 46958 39058
rect 47010 39006 47012 39058
rect 46844 39004 47012 39006
rect 46956 38948 47012 39004
rect 46956 38882 47012 38892
rect 47740 39060 47796 39070
rect 47740 38946 47796 39004
rect 47740 38894 47742 38946
rect 47794 38894 47796 38946
rect 47740 38882 47796 38894
rect 47852 38948 47908 38958
rect 47852 38854 47908 38892
rect 47964 38946 48020 39564
rect 47964 38894 47966 38946
rect 48018 38894 48020 38946
rect 47964 38882 48020 38894
rect 46620 38836 46676 38846
rect 46620 38668 46676 38780
rect 48076 38668 48132 40236
rect 46620 38612 47124 38668
rect 47068 38050 47124 38612
rect 47292 38612 47348 38622
rect 47964 38612 48132 38668
rect 47292 38610 47796 38612
rect 47292 38558 47294 38610
rect 47346 38558 47796 38610
rect 47292 38556 47796 38558
rect 47292 38546 47348 38556
rect 47068 37998 47070 38050
rect 47122 37998 47124 38050
rect 47068 37986 47124 37998
rect 46452 36764 46564 36820
rect 46620 37268 46676 37278
rect 45500 34914 45668 34916
rect 45500 34862 45502 34914
rect 45554 34862 45668 34914
rect 45500 34860 45668 34862
rect 45836 34972 46228 35028
rect 46284 36708 46340 36718
rect 45164 34690 45220 34702
rect 45164 34638 45166 34690
rect 45218 34638 45220 34690
rect 45164 34244 45220 34638
rect 45164 34178 45220 34188
rect 44044 33518 44046 33570
rect 44098 33518 44100 33570
rect 44044 33506 44100 33518
rect 44156 33628 44660 33684
rect 44716 33796 44772 33806
rect 43932 33348 43988 33358
rect 44156 33348 44212 33628
rect 44716 33572 44772 33740
rect 45500 33796 45556 34860
rect 45724 34804 45780 34814
rect 45724 34710 45780 34748
rect 45836 33796 45892 34972
rect 46284 34916 46340 36652
rect 46396 36370 46452 36764
rect 46396 36318 46398 36370
rect 46450 36318 46452 36370
rect 46396 36306 46452 36318
rect 46620 35812 46676 37212
rect 47404 37156 47460 37166
rect 46844 37044 46900 37054
rect 46844 36594 46900 36988
rect 46844 36542 46846 36594
rect 46898 36542 46900 36594
rect 46844 36530 46900 36542
rect 47180 36484 47236 36494
rect 45500 33730 45556 33740
rect 45724 33740 45892 33796
rect 45948 34914 46340 34916
rect 45948 34862 46286 34914
rect 46338 34862 46340 34914
rect 45948 34860 46340 34862
rect 45948 34018 46004 34860
rect 46284 34850 46340 34860
rect 46508 35756 46676 35812
rect 47068 36372 47124 36382
rect 47068 35924 47124 36316
rect 47068 35810 47124 35868
rect 47068 35758 47070 35810
rect 47122 35758 47124 35810
rect 46396 34804 46452 34814
rect 46396 34710 46452 34748
rect 46396 34356 46452 34366
rect 46508 34356 46564 35756
rect 47068 35746 47124 35758
rect 46620 35586 46676 35598
rect 46620 35534 46622 35586
rect 46674 35534 46676 35586
rect 46620 34692 46676 35534
rect 47068 35364 47124 35374
rect 47068 34914 47124 35308
rect 47180 35026 47236 36428
rect 47180 34974 47182 35026
rect 47234 34974 47236 35026
rect 47180 34962 47236 34974
rect 47292 35476 47348 35486
rect 47068 34862 47070 34914
rect 47122 34862 47124 34914
rect 47068 34850 47124 34862
rect 47292 34914 47348 35420
rect 47292 34862 47294 34914
rect 47346 34862 47348 34914
rect 47292 34850 47348 34862
rect 46844 34692 46900 34702
rect 46620 34690 46900 34692
rect 46620 34638 46846 34690
rect 46898 34638 46900 34690
rect 46620 34636 46900 34638
rect 46396 34354 46564 34356
rect 46396 34302 46398 34354
rect 46450 34302 46564 34354
rect 46396 34300 46564 34302
rect 46396 34290 46452 34300
rect 45948 33966 45950 34018
rect 46002 33966 46004 34018
rect 43932 33346 44212 33348
rect 43932 33294 43934 33346
rect 43986 33294 44212 33346
rect 43932 33292 44212 33294
rect 44604 33516 44772 33572
rect 43932 33282 43988 33292
rect 43260 31266 43316 31276
rect 43372 32508 43540 32564
rect 43596 32844 43764 32900
rect 43820 33122 43876 33134
rect 43820 33070 43822 33122
rect 43874 33070 43876 33122
rect 43148 31166 43150 31218
rect 43202 31166 43204 31218
rect 42364 30212 42420 30222
rect 42476 30212 42532 30380
rect 42420 30156 42532 30212
rect 42588 30212 42644 30222
rect 43036 30212 43092 30222
rect 43148 30212 43204 31166
rect 43372 30884 43428 32508
rect 43484 31332 43540 31342
rect 43484 31218 43540 31276
rect 43484 31166 43486 31218
rect 43538 31166 43540 31218
rect 43484 31154 43540 31166
rect 43372 30828 43540 30884
rect 42588 30210 43204 30212
rect 42588 30158 42590 30210
rect 42642 30158 43038 30210
rect 43090 30158 43204 30210
rect 42588 30156 43204 30158
rect 42364 30146 42420 30156
rect 42588 30146 42644 30156
rect 43036 30146 43092 30156
rect 43372 30100 43428 30110
rect 42252 29362 42308 29372
rect 43260 29988 43316 29998
rect 42476 28812 42756 28868
rect 42364 28756 42420 28766
rect 42476 28756 42532 28812
rect 42364 28754 42532 28756
rect 42364 28702 42366 28754
rect 42418 28702 42532 28754
rect 42364 28700 42532 28702
rect 42364 28690 42420 28700
rect 42588 28644 42644 28654
rect 41804 27134 41806 27186
rect 41858 27134 41860 27186
rect 41132 26962 41188 26974
rect 41132 26910 41134 26962
rect 41186 26910 41188 26962
rect 41132 26628 41188 26910
rect 41244 26852 41300 26862
rect 41244 26758 41300 26796
rect 41132 26562 41188 26572
rect 41020 26348 41188 26404
rect 40908 26290 40964 26302
rect 40908 26238 40910 26290
rect 40962 26238 40964 26290
rect 40796 25508 40852 25518
rect 40796 25414 40852 25452
rect 40908 25172 40964 26238
rect 40908 25106 40964 25116
rect 41020 26178 41076 26190
rect 41020 26126 41022 26178
rect 41074 26126 41076 26178
rect 41020 24948 41076 26126
rect 41132 25060 41188 26348
rect 41244 26290 41300 26302
rect 41244 26238 41246 26290
rect 41298 26238 41300 26290
rect 41244 25844 41300 26238
rect 41356 26292 41412 27132
rect 41804 27122 41860 27134
rect 42028 27244 42140 27300
rect 41916 27076 41972 27086
rect 41916 26982 41972 27020
rect 41692 26962 41748 26974
rect 41692 26910 41694 26962
rect 41746 26910 41748 26962
rect 41692 26908 41748 26910
rect 42028 26908 42084 27244
rect 42140 27234 42196 27244
rect 42252 28418 42308 28430
rect 42252 28366 42254 28418
rect 42306 28366 42308 28418
rect 41692 26852 42084 26908
rect 42140 27074 42196 27086
rect 42140 27022 42142 27074
rect 42194 27022 42196 27074
rect 41356 26226 41412 26236
rect 41468 26290 41524 26302
rect 41468 26238 41470 26290
rect 41522 26238 41524 26290
rect 41244 25788 41412 25844
rect 41244 25618 41300 25630
rect 41244 25566 41246 25618
rect 41298 25566 41300 25618
rect 41244 25396 41300 25566
rect 41244 25330 41300 25340
rect 41356 25284 41412 25788
rect 41356 25218 41412 25228
rect 41132 24994 41188 25004
rect 40684 24892 41076 24948
rect 40684 23716 40740 24892
rect 41244 24836 41300 24846
rect 40684 23650 40740 23660
rect 40796 24724 40852 24734
rect 40796 23380 40852 24668
rect 41020 24724 41076 24734
rect 41020 24630 41076 24668
rect 41132 24722 41188 24734
rect 41132 24670 41134 24722
rect 41186 24670 41188 24722
rect 41132 24164 41188 24670
rect 41244 24722 41300 24780
rect 41244 24670 41246 24722
rect 41298 24670 41300 24722
rect 41244 24658 41300 24670
rect 41132 24108 41300 24164
rect 40796 23314 40852 23324
rect 40908 23828 40964 23838
rect 40572 22652 40852 22708
rect 40572 22484 40628 22494
rect 40460 22482 40628 22484
rect 40460 22430 40574 22482
rect 40626 22430 40628 22482
rect 40460 22428 40628 22430
rect 40572 22418 40628 22428
rect 40684 22372 40740 22382
rect 40796 22372 40852 22652
rect 40908 22594 40964 23772
rect 41132 23826 41188 23838
rect 41132 23774 41134 23826
rect 41186 23774 41188 23826
rect 41132 22708 41188 23774
rect 41132 22642 41188 22652
rect 41244 23268 41300 24108
rect 41356 23828 41412 23838
rect 41468 23828 41524 26238
rect 41916 26292 41972 26302
rect 41916 26198 41972 26236
rect 41692 25508 41748 25518
rect 41692 24946 41748 25452
rect 42140 25396 42196 27022
rect 42252 27076 42308 28366
rect 42476 28420 42532 28430
rect 42476 28326 42532 28364
rect 42588 28196 42644 28588
rect 42364 28140 42644 28196
rect 42364 27970 42420 28140
rect 42364 27918 42366 27970
rect 42418 27918 42420 27970
rect 42364 27906 42420 27918
rect 42700 27524 42756 28812
rect 42924 28644 42980 28654
rect 43260 28644 43316 29932
rect 43372 28756 43428 30044
rect 43484 29428 43540 30828
rect 43596 30212 43652 32844
rect 43820 32788 43876 33070
rect 43820 32722 43876 32732
rect 43708 32564 43764 32574
rect 43708 32470 43764 32508
rect 43932 32562 43988 32574
rect 43932 32510 43934 32562
rect 43986 32510 43988 32562
rect 43820 32452 43876 32462
rect 43820 32358 43876 32396
rect 43932 31668 43988 32510
rect 44380 32562 44436 32574
rect 44380 32510 44382 32562
rect 44434 32510 44436 32562
rect 44268 31890 44324 31902
rect 44268 31838 44270 31890
rect 44322 31838 44324 31890
rect 43932 31602 43988 31612
rect 44044 31780 44100 31790
rect 44044 30884 44100 31724
rect 44268 31780 44324 31838
rect 44268 31714 44324 31724
rect 44268 31220 44324 31230
rect 44380 31220 44436 32510
rect 44268 31218 44436 31220
rect 44268 31166 44270 31218
rect 44322 31166 44436 31218
rect 44268 31164 44436 31166
rect 44268 31154 44324 31164
rect 44156 31108 44212 31118
rect 44156 31014 44212 31052
rect 44380 30994 44436 31006
rect 44380 30942 44382 30994
rect 44434 30942 44436 30994
rect 44380 30884 44436 30942
rect 44044 30828 44436 30884
rect 43596 30156 43876 30212
rect 43484 29362 43540 29372
rect 43596 28980 43652 28990
rect 43372 28662 43428 28700
rect 43484 28924 43596 28980
rect 42924 28642 43316 28644
rect 42924 28590 42926 28642
rect 42978 28590 43316 28642
rect 42924 28588 43316 28590
rect 42924 28578 42980 28588
rect 43484 28532 43540 28924
rect 43596 28914 43652 28924
rect 43820 28868 43876 30156
rect 44492 29316 44548 29326
rect 44492 29222 44548 29260
rect 43820 28754 43876 28812
rect 44268 29092 44324 29102
rect 44604 29092 44660 33516
rect 45388 33012 45444 33022
rect 44828 32340 44884 32350
rect 44716 31106 44772 31118
rect 44716 31054 44718 31106
rect 44770 31054 44772 31106
rect 44716 30996 44772 31054
rect 44716 30930 44772 30940
rect 44828 29540 44884 32284
rect 44940 31892 44996 31902
rect 44940 31798 44996 31836
rect 45388 31332 45444 32956
rect 44940 31220 44996 31230
rect 44940 30994 44996 31164
rect 44940 30942 44942 30994
rect 44994 30942 44996 30994
rect 44940 30930 44996 30942
rect 45276 30996 45332 31006
rect 45388 30996 45444 31276
rect 45500 31220 45556 31230
rect 45724 31220 45780 33740
rect 45836 33572 45892 33582
rect 45836 32562 45892 33516
rect 45836 32510 45838 32562
rect 45890 32510 45892 32562
rect 45836 32498 45892 32510
rect 45948 32564 46004 33966
rect 46508 33348 46564 33358
rect 46508 33234 46564 33292
rect 46508 33182 46510 33234
rect 46562 33182 46564 33234
rect 46508 33170 46564 33182
rect 46732 33234 46788 33246
rect 46732 33182 46734 33234
rect 46786 33182 46788 33234
rect 46620 33122 46676 33134
rect 46620 33070 46622 33122
rect 46674 33070 46676 33122
rect 46396 32788 46452 32798
rect 46396 32694 46452 32732
rect 46620 32676 46676 33070
rect 46732 32788 46788 33182
rect 46844 33012 46900 34636
rect 47068 33684 47124 33694
rect 47068 33346 47124 33628
rect 47068 33294 47070 33346
rect 47122 33294 47124 33346
rect 47068 33282 47124 33294
rect 47180 33570 47236 33582
rect 47180 33518 47182 33570
rect 47234 33518 47236 33570
rect 47180 33348 47236 33518
rect 47180 33282 47236 33292
rect 47180 33124 47236 33134
rect 47180 33030 47236 33068
rect 46844 32946 46900 32956
rect 47404 32900 47460 37100
rect 47628 36596 47684 36606
rect 47516 36372 47572 36382
rect 47516 36278 47572 36316
rect 47628 35924 47684 36540
rect 47740 36482 47796 38556
rect 47740 36430 47742 36482
rect 47794 36430 47796 36482
rect 47740 36260 47796 36430
rect 47740 36194 47796 36204
rect 47964 35924 48020 38612
rect 48188 37940 48244 40350
rect 48300 38836 48356 40908
rect 48748 40740 48804 41132
rect 48860 41076 48916 41244
rect 48860 41010 48916 41020
rect 48748 40684 48916 40740
rect 48748 40402 48804 40414
rect 48748 40350 48750 40402
rect 48802 40350 48804 40402
rect 48412 39620 48468 39630
rect 48636 39620 48692 39630
rect 48412 39618 48692 39620
rect 48412 39566 48414 39618
rect 48466 39566 48638 39618
rect 48690 39566 48692 39618
rect 48412 39564 48692 39566
rect 48412 39554 48468 39564
rect 48636 39554 48692 39564
rect 48748 38948 48804 40350
rect 48860 39730 48916 40684
rect 48860 39678 48862 39730
rect 48914 39678 48916 39730
rect 48860 39666 48916 39678
rect 48972 40626 49028 41804
rect 49420 41748 49476 41918
rect 49756 41970 49812 42588
rect 49756 41918 49758 41970
rect 49810 41918 49812 41970
rect 49756 41906 49812 41918
rect 50316 42532 50372 43596
rect 50428 43586 50484 43596
rect 50876 43428 50932 44046
rect 51100 43428 51156 43438
rect 50876 43372 51100 43428
rect 51100 43334 51156 43372
rect 51324 43314 51380 43326
rect 51660 43316 51716 43326
rect 51324 43262 51326 43314
rect 51378 43262 51380 43314
rect 51324 43204 51380 43262
rect 51324 43138 51380 43148
rect 51548 43260 51660 43316
rect 49420 41682 49476 41692
rect 49980 41412 50036 41422
rect 49980 41318 50036 41356
rect 49980 41076 50036 41086
rect 49980 40982 50036 41020
rect 50092 41076 50148 41086
rect 50316 41076 50372 42476
rect 50428 42756 50484 42766
rect 50540 42756 50596 42766
rect 50484 42754 50596 42756
rect 50484 42702 50542 42754
rect 50594 42702 50596 42754
rect 50484 42700 50596 42702
rect 50428 42196 50484 42700
rect 50540 42690 50596 42700
rect 50764 42754 50820 42766
rect 50764 42702 50766 42754
rect 50818 42702 50820 42754
rect 50764 42532 50820 42702
rect 51100 42644 51156 42654
rect 51436 42644 51492 42654
rect 51100 42642 51492 42644
rect 51100 42590 51102 42642
rect 51154 42590 51438 42642
rect 51490 42590 51492 42642
rect 51100 42588 51492 42590
rect 51100 42578 51156 42588
rect 51436 42578 51492 42588
rect 50764 42466 50820 42476
rect 50988 42532 51044 42542
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50428 42140 50596 42196
rect 50428 41076 50484 41086
rect 50092 41074 50260 41076
rect 50092 41022 50094 41074
rect 50146 41022 50260 41074
rect 50092 41020 50260 41022
rect 50316 41074 50484 41076
rect 50316 41022 50430 41074
rect 50482 41022 50484 41074
rect 50316 41020 50484 41022
rect 50092 41010 50148 41020
rect 49420 40962 49476 40974
rect 49420 40910 49422 40962
rect 49474 40910 49476 40962
rect 48972 40574 48974 40626
rect 49026 40574 49028 40626
rect 48748 38882 48804 38892
rect 48972 39620 49028 40574
rect 49196 40628 49252 40638
rect 49196 40534 49252 40572
rect 49420 40516 49476 40910
rect 48300 38770 48356 38780
rect 48300 38612 48356 38622
rect 48300 38050 48356 38556
rect 48300 37998 48302 38050
rect 48354 37998 48356 38050
rect 48300 37986 48356 37998
rect 48972 38050 49028 39564
rect 48972 37998 48974 38050
rect 49026 37998 49028 38050
rect 48972 37986 49028 37998
rect 49084 40292 49140 40302
rect 49084 39508 49140 40236
rect 48188 37154 48244 37884
rect 48860 37938 48916 37950
rect 48860 37886 48862 37938
rect 48914 37886 48916 37938
rect 48860 37492 48916 37886
rect 48188 37102 48190 37154
rect 48242 37102 48244 37154
rect 48188 36484 48244 37102
rect 48524 37436 48916 37492
rect 48188 36482 48356 36484
rect 48188 36430 48190 36482
rect 48242 36430 48356 36482
rect 48188 36428 48356 36430
rect 48188 36418 48244 36428
rect 47516 35868 47684 35924
rect 47740 35868 48020 35924
rect 48076 36148 48132 36158
rect 47516 35364 47572 35868
rect 47516 35298 47572 35308
rect 47628 35698 47684 35710
rect 47628 35646 47630 35698
rect 47682 35646 47684 35698
rect 47628 34804 47684 35646
rect 47628 34130 47684 34748
rect 47628 34078 47630 34130
rect 47682 34078 47684 34130
rect 47628 34066 47684 34078
rect 47180 32844 47460 32900
rect 46844 32788 46900 32798
rect 46732 32786 46900 32788
rect 46732 32734 46846 32786
rect 46898 32734 46900 32786
rect 46732 32732 46900 32734
rect 46844 32722 46900 32732
rect 47180 32786 47236 32844
rect 47180 32734 47182 32786
rect 47234 32734 47236 32786
rect 47180 32722 47236 32734
rect 47516 32788 47572 32798
rect 46956 32676 47012 32686
rect 46620 32620 46788 32676
rect 46060 32564 46116 32574
rect 45948 32562 46116 32564
rect 45948 32510 46062 32562
rect 46114 32510 46116 32562
rect 45948 32508 46116 32510
rect 46060 32498 46116 32508
rect 46284 32340 46340 32350
rect 46284 32246 46340 32284
rect 46508 32340 46564 32350
rect 46508 32338 46676 32340
rect 46508 32286 46510 32338
rect 46562 32286 46676 32338
rect 46508 32284 46676 32286
rect 46508 32274 46564 32284
rect 46284 31892 46340 31902
rect 45724 31164 46116 31220
rect 45500 31126 45556 31164
rect 45388 30940 45556 30996
rect 45052 30772 45108 30782
rect 45052 30678 45108 30716
rect 44828 29484 44996 29540
rect 44716 29428 44772 29438
rect 44772 29372 44884 29428
rect 44716 29362 44772 29372
rect 44828 29314 44884 29372
rect 44828 29262 44830 29314
rect 44882 29262 44884 29314
rect 44828 29250 44884 29262
rect 44324 29036 44660 29092
rect 43820 28702 43822 28754
rect 43874 28702 43876 28754
rect 43820 28690 43876 28702
rect 44044 28756 44100 28766
rect 43148 28476 43540 28532
rect 42364 27468 42756 27524
rect 43036 27524 43092 27534
rect 42364 27298 42420 27468
rect 42364 27246 42366 27298
rect 42418 27246 42420 27298
rect 42364 27234 42420 27246
rect 42924 27300 42980 27310
rect 42252 27010 42308 27020
rect 42812 27076 42868 27086
rect 42812 26982 42868 27020
rect 42700 26962 42756 26974
rect 42700 26910 42702 26962
rect 42754 26910 42756 26962
rect 42700 26908 42756 26910
rect 42476 26852 42756 26908
rect 42476 25844 42532 26852
rect 42476 25778 42532 25788
rect 42588 26628 42644 26638
rect 42252 25508 42308 25518
rect 42252 25414 42308 25452
rect 42028 25340 42196 25396
rect 42588 25394 42644 26572
rect 42700 26516 42756 26526
rect 42924 26516 42980 27244
rect 42700 26514 42980 26516
rect 42700 26462 42702 26514
rect 42754 26462 42980 26514
rect 42700 26460 42980 26462
rect 43036 26962 43092 27468
rect 43036 26910 43038 26962
rect 43090 26910 43092 26962
rect 42700 26450 42756 26460
rect 43036 25844 43092 26910
rect 42588 25342 42590 25394
rect 42642 25342 42644 25394
rect 42028 25284 42084 25340
rect 42028 25218 42084 25228
rect 42476 25284 42532 25294
rect 41692 24894 41694 24946
rect 41746 24894 41748 24946
rect 41692 24882 41748 24894
rect 42140 25172 42196 25182
rect 41804 24164 41860 24174
rect 41412 23772 41524 23828
rect 41692 23938 41748 23950
rect 41692 23886 41694 23938
rect 41746 23886 41748 23938
rect 41356 23762 41412 23772
rect 41692 23604 41748 23886
rect 41692 23538 41748 23548
rect 41804 23716 41860 24108
rect 42028 23938 42084 23950
rect 42028 23886 42030 23938
rect 42082 23886 42084 23938
rect 42028 23828 42084 23886
rect 42028 23762 42084 23772
rect 42140 23828 42196 25116
rect 42476 24610 42532 25228
rect 42476 24558 42478 24610
rect 42530 24558 42532 24610
rect 42140 23826 42308 23828
rect 42140 23774 42142 23826
rect 42194 23774 42308 23826
rect 42140 23772 42308 23774
rect 42140 23762 42196 23772
rect 41804 23378 41860 23660
rect 41804 23326 41806 23378
rect 41858 23326 41860 23378
rect 41804 23314 41860 23326
rect 40908 22542 40910 22594
rect 40962 22542 40964 22594
rect 40908 22530 40964 22542
rect 41244 22596 41300 23212
rect 42252 23268 42308 23772
rect 42140 23044 42196 23054
rect 42140 22950 42196 22988
rect 42028 22708 42084 22718
rect 42084 22652 42196 22708
rect 42028 22642 42084 22652
rect 41244 22530 41300 22540
rect 42028 22484 42084 22494
rect 42028 22390 42084 22428
rect 40796 22316 41636 22372
rect 40684 22278 40740 22316
rect 40236 22194 40292 22204
rect 41020 22148 41076 22158
rect 38892 21758 38894 21810
rect 38946 21758 38948 21810
rect 38892 21746 38948 21758
rect 40124 22036 40180 22046
rect 39900 21700 39956 21710
rect 39900 21586 39956 21644
rect 39900 21534 39902 21586
rect 39954 21534 39956 21586
rect 39900 21522 39956 21534
rect 40124 21586 40180 21980
rect 41020 21700 41076 22092
rect 40124 21534 40126 21586
rect 40178 21534 40180 21586
rect 40124 21522 40180 21534
rect 40460 21698 41076 21700
rect 40460 21646 41022 21698
rect 41074 21646 41076 21698
rect 40460 21644 41076 21646
rect 40460 21586 40516 21644
rect 41020 21634 41076 21644
rect 40460 21534 40462 21586
rect 40514 21534 40516 21586
rect 40460 21522 40516 21534
rect 40236 21476 40292 21486
rect 40236 21382 40292 21420
rect 37212 20914 37492 20916
rect 37212 20862 37214 20914
rect 37266 20862 37492 20914
rect 37212 20860 37492 20862
rect 37212 20850 37268 20860
rect 38444 20802 38500 20814
rect 38444 20750 38446 20802
rect 38498 20750 38500 20802
rect 36988 20076 37492 20132
rect 36988 19348 37044 20076
rect 37436 20018 37492 20076
rect 37436 19966 37438 20018
rect 37490 19966 37492 20018
rect 37436 19954 37492 19966
rect 37100 19908 37156 19918
rect 38444 19908 38500 20750
rect 39116 20690 39172 20702
rect 39116 20638 39118 20690
rect 39170 20638 39172 20690
rect 39116 20580 39172 20638
rect 39116 20514 39172 20524
rect 41132 20242 41188 22316
rect 41244 21588 41300 21598
rect 41244 20916 41300 21532
rect 41244 20914 41524 20916
rect 41244 20862 41246 20914
rect 41298 20862 41524 20914
rect 41244 20860 41524 20862
rect 41244 20850 41300 20860
rect 41132 20190 41134 20242
rect 41186 20190 41188 20242
rect 41132 20178 41188 20190
rect 41468 20132 41524 20860
rect 41580 20802 41636 22316
rect 42028 21586 42084 21598
rect 42028 21534 42030 21586
rect 42082 21534 42084 21586
rect 41804 21476 41860 21486
rect 41804 21026 41860 21420
rect 41804 20974 41806 21026
rect 41858 20974 41860 21026
rect 41804 20962 41860 20974
rect 42028 20804 42084 21534
rect 42140 21474 42196 22652
rect 42252 22148 42308 23212
rect 42252 22082 42308 22092
rect 42476 22932 42532 24558
rect 42588 23826 42644 25342
rect 42588 23774 42590 23826
rect 42642 23774 42644 23826
rect 42588 23762 42644 23774
rect 42700 25788 43092 25844
rect 42700 24834 42756 25788
rect 43148 25732 43204 28476
rect 43260 28308 43316 28318
rect 43260 27074 43316 28252
rect 43596 27524 43652 27534
rect 43596 27186 43652 27468
rect 43596 27134 43598 27186
rect 43650 27134 43652 27186
rect 43596 27122 43652 27134
rect 43260 27022 43262 27074
rect 43314 27022 43316 27074
rect 43260 26964 43316 27022
rect 44044 27076 44100 28700
rect 44268 28754 44324 29036
rect 44268 28702 44270 28754
rect 44322 28702 44324 28754
rect 44268 28532 44324 28702
rect 44268 28466 44324 28476
rect 44828 28756 44884 28766
rect 44828 27858 44884 28700
rect 44940 28084 44996 29484
rect 45164 29428 45220 29466
rect 45164 29362 45220 29372
rect 45276 29428 45332 30940
rect 45388 29428 45444 29438
rect 45276 29426 45444 29428
rect 45276 29374 45390 29426
rect 45442 29374 45444 29426
rect 45276 29372 45444 29374
rect 45164 29204 45220 29214
rect 45164 28866 45220 29148
rect 45164 28814 45166 28866
rect 45218 28814 45220 28866
rect 45164 28802 45220 28814
rect 44940 28018 44996 28028
rect 45052 28530 45108 28542
rect 45052 28478 45054 28530
rect 45106 28478 45108 28530
rect 44828 27806 44830 27858
rect 44882 27806 44884 27858
rect 44828 27794 44884 27806
rect 44492 27746 44548 27758
rect 44492 27694 44494 27746
rect 44546 27694 44548 27746
rect 44492 27636 44548 27694
rect 45052 27636 45108 28478
rect 43260 26898 43316 26908
rect 43484 26964 43540 26974
rect 43484 26516 43540 26908
rect 43932 26852 43988 26862
rect 43596 26516 43652 26526
rect 43484 26514 43652 26516
rect 43484 26462 43598 26514
rect 43650 26462 43652 26514
rect 43484 26460 43652 26462
rect 43596 26450 43652 26460
rect 42924 25676 43204 25732
rect 43484 25844 43540 25854
rect 42812 25508 42868 25518
rect 42812 25414 42868 25452
rect 42700 24782 42702 24834
rect 42754 24782 42756 24834
rect 42700 24724 42756 24782
rect 42588 23268 42644 23278
rect 42700 23268 42756 24668
rect 42588 23266 42756 23268
rect 42588 23214 42590 23266
rect 42642 23214 42756 23266
rect 42588 23212 42756 23214
rect 42812 23380 42868 23390
rect 42588 23202 42644 23212
rect 42476 22036 42532 22876
rect 42588 22484 42644 22494
rect 42588 22370 42644 22428
rect 42588 22318 42590 22370
rect 42642 22318 42644 22370
rect 42588 22306 42644 22318
rect 42812 22370 42868 23324
rect 42812 22318 42814 22370
rect 42866 22318 42868 22370
rect 42812 22148 42868 22318
rect 42812 22082 42868 22092
rect 42476 21970 42532 21980
rect 42140 21422 42142 21474
rect 42194 21422 42196 21474
rect 42140 21410 42196 21422
rect 42812 20916 42868 20926
rect 42924 20916 42980 25676
rect 43148 25506 43204 25518
rect 43148 25454 43150 25506
rect 43202 25454 43204 25506
rect 43036 23714 43092 23726
rect 43036 23662 43038 23714
rect 43090 23662 43092 23714
rect 43036 23156 43092 23662
rect 43036 23090 43092 23100
rect 43148 22372 43204 25454
rect 43484 24722 43540 25788
rect 43484 24670 43486 24722
rect 43538 24670 43540 24722
rect 43484 24658 43540 24670
rect 43596 25620 43652 25630
rect 43148 22306 43204 22316
rect 43484 23604 43540 23614
rect 43372 22260 43428 22270
rect 43372 22166 43428 22204
rect 43036 21588 43092 21598
rect 43036 21494 43092 21532
rect 43484 21474 43540 23548
rect 43596 23154 43652 25564
rect 43708 25508 43764 25518
rect 43708 24050 43764 25452
rect 43932 24722 43988 26796
rect 44044 26514 44100 27020
rect 44044 26462 44046 26514
rect 44098 26462 44100 26514
rect 44044 26450 44100 26462
rect 44156 27580 45108 27636
rect 44156 27074 44212 27580
rect 45276 27524 45332 29372
rect 45388 29362 45444 29372
rect 45500 29204 45556 30940
rect 45612 30994 45668 31006
rect 45612 30942 45614 30994
rect 45666 30942 45668 30994
rect 45612 30772 45668 30942
rect 45612 30100 45668 30716
rect 46060 30100 46116 31164
rect 45612 30034 45668 30044
rect 45836 30098 46116 30100
rect 45836 30046 46062 30098
rect 46114 30046 46116 30098
rect 45836 30044 46116 30046
rect 45724 29986 45780 29998
rect 45724 29934 45726 29986
rect 45778 29934 45780 29986
rect 45724 29876 45780 29934
rect 45724 29810 45780 29820
rect 45836 29764 45892 30044
rect 46060 30034 46116 30044
rect 45836 29698 45892 29708
rect 46060 29652 46116 29662
rect 45836 29540 45892 29550
rect 45724 29428 45780 29438
rect 45388 29148 45556 29204
rect 45612 29314 45668 29326
rect 45612 29262 45614 29314
rect 45666 29262 45668 29314
rect 45388 28756 45444 29148
rect 45388 28690 45444 28700
rect 45500 28868 45556 28878
rect 44828 27468 45332 27524
rect 44828 27186 44884 27468
rect 45052 27300 45108 27310
rect 45052 27206 45108 27244
rect 44828 27134 44830 27186
rect 44882 27134 44884 27186
rect 44828 27122 44884 27134
rect 45276 27188 45332 27198
rect 44156 27022 44158 27074
rect 44210 27022 44212 27074
rect 44156 25620 44212 27022
rect 45276 26516 45332 27132
rect 45276 26450 45332 26460
rect 45388 27186 45444 27198
rect 45388 27134 45390 27186
rect 45442 27134 45444 27186
rect 44492 26402 44548 26414
rect 44492 26350 44494 26402
rect 44546 26350 44548 26402
rect 44380 26292 44436 26302
rect 43932 24670 43934 24722
rect 43986 24670 43988 24722
rect 43932 24658 43988 24670
rect 44044 25564 44212 25620
rect 44268 26290 44436 26292
rect 44268 26238 44382 26290
rect 44434 26238 44436 26290
rect 44268 26236 44436 26238
rect 44044 25396 44100 25564
rect 44268 25508 44324 26236
rect 44380 26226 44436 26236
rect 43932 24164 43988 24174
rect 44044 24164 44100 25340
rect 44156 25452 44324 25508
rect 44156 25394 44212 25452
rect 44156 25342 44158 25394
rect 44210 25342 44212 25394
rect 44156 25284 44212 25342
rect 44156 25218 44212 25228
rect 44268 25282 44324 25294
rect 44268 25230 44270 25282
rect 44322 25230 44324 25282
rect 44268 24612 44324 25230
rect 44268 24546 44324 24556
rect 43932 24162 44100 24164
rect 43932 24110 43934 24162
rect 43986 24110 44100 24162
rect 43932 24108 44100 24110
rect 43932 24098 43988 24108
rect 43708 23998 43710 24050
rect 43762 23998 43764 24050
rect 43708 23986 43764 23998
rect 44492 23940 44548 26350
rect 45388 26292 45444 27134
rect 45388 26226 45444 26236
rect 45388 25844 45444 25854
rect 45276 25788 45388 25844
rect 45276 25618 45332 25788
rect 45388 25778 45444 25788
rect 45276 25566 45278 25618
rect 45330 25566 45332 25618
rect 45276 25554 45332 25566
rect 44940 25508 44996 25518
rect 44940 25414 44996 25452
rect 45388 24722 45444 24734
rect 45388 24670 45390 24722
rect 45442 24670 45444 24722
rect 43932 23884 44548 23940
rect 44940 24612 44996 24622
rect 44940 23938 44996 24556
rect 45388 24164 45444 24670
rect 45276 24108 45444 24164
rect 44940 23886 44942 23938
rect 44994 23886 44996 23938
rect 43596 23102 43598 23154
rect 43650 23102 43652 23154
rect 43596 23090 43652 23102
rect 43820 23156 43876 23166
rect 43820 23062 43876 23100
rect 43484 21422 43486 21474
rect 43538 21422 43540 21474
rect 43484 21410 43540 21422
rect 43932 21476 43988 23884
rect 44940 23874 44996 23886
rect 45164 23940 45220 23950
rect 45164 23846 45220 23884
rect 44268 23714 44324 23726
rect 44268 23662 44270 23714
rect 44322 23662 44324 23714
rect 44268 22260 44324 23662
rect 45276 23156 45332 24108
rect 45388 23940 45444 23950
rect 45500 23940 45556 28812
rect 45612 28642 45668 29262
rect 45612 28590 45614 28642
rect 45666 28590 45668 28642
rect 45612 28578 45668 28590
rect 45724 28420 45780 29372
rect 45612 28364 45780 28420
rect 45836 29426 45892 29484
rect 46060 29538 46116 29596
rect 46060 29486 46062 29538
rect 46114 29486 46116 29538
rect 46060 29474 46116 29486
rect 45836 29374 45838 29426
rect 45890 29374 45892 29426
rect 45612 26908 45668 28364
rect 45836 27300 45892 29374
rect 46172 29314 46228 29326
rect 46172 29262 46174 29314
rect 46226 29262 46228 29314
rect 46172 28644 46228 29262
rect 46172 28578 46228 28588
rect 46284 27746 46340 31836
rect 46508 30996 46564 31006
rect 46508 30436 46564 30940
rect 46508 30370 46564 30380
rect 46396 30212 46452 30250
rect 46396 30146 46452 30156
rect 46620 29652 46676 32284
rect 46732 32116 46788 32620
rect 46956 32582 47012 32620
rect 47516 32562 47572 32732
rect 47516 32510 47518 32562
rect 47570 32510 47572 32562
rect 47516 32498 47572 32510
rect 47740 32564 47796 35868
rect 47740 32498 47796 32508
rect 47852 35700 47908 35710
rect 46788 32060 47012 32116
rect 46732 32022 46788 32060
rect 46956 32002 47012 32060
rect 46956 31950 46958 32002
rect 47010 31950 47012 32002
rect 46956 31938 47012 31950
rect 46732 31778 46788 31790
rect 46732 31726 46734 31778
rect 46786 31726 46788 31778
rect 46732 31444 46788 31726
rect 47180 31778 47236 31790
rect 47180 31726 47182 31778
rect 47234 31726 47236 31778
rect 46844 31444 46900 31454
rect 46732 31388 46844 31444
rect 46844 31378 46900 31388
rect 47180 30996 47236 31726
rect 47628 31556 47684 31566
rect 47628 31462 47684 31500
rect 47180 30930 47236 30940
rect 47404 30994 47460 31006
rect 47404 30942 47406 30994
rect 47458 30942 47460 30994
rect 46732 30884 46788 30894
rect 46732 30790 46788 30828
rect 46956 30772 47012 30782
rect 46844 30770 47012 30772
rect 46844 30718 46958 30770
rect 47010 30718 47012 30770
rect 46844 30716 47012 30718
rect 46844 30324 46900 30716
rect 46956 30706 47012 30716
rect 47068 30772 47124 30782
rect 47404 30772 47460 30942
rect 47068 30770 47460 30772
rect 47068 30718 47070 30770
rect 47122 30718 47460 30770
rect 47068 30716 47460 30718
rect 47068 30436 47124 30716
rect 46844 30258 46900 30268
rect 46956 30380 47124 30436
rect 46956 30212 47012 30380
rect 47740 30324 47796 30334
rect 47740 30230 47796 30268
rect 46956 30146 47012 30156
rect 47068 30212 47124 30222
rect 47068 30210 47236 30212
rect 47068 30158 47070 30210
rect 47122 30158 47236 30210
rect 47068 30156 47236 30158
rect 47068 30146 47124 30156
rect 46732 29988 46788 29998
rect 46732 29986 47012 29988
rect 46732 29934 46734 29986
rect 46786 29934 47012 29986
rect 46732 29932 47012 29934
rect 46732 29922 46788 29932
rect 46956 29876 47012 29932
rect 46956 29820 47068 29876
rect 47012 29662 47068 29820
rect 46396 29596 46676 29652
rect 46956 29652 47068 29662
rect 47012 29596 47068 29652
rect 47180 29652 47236 30156
rect 47852 30210 47908 35644
rect 47964 35700 48020 35710
rect 48076 35700 48132 36092
rect 47964 35698 48132 35700
rect 47964 35646 47966 35698
rect 48018 35646 48132 35698
rect 47964 35644 48132 35646
rect 47964 35634 48020 35644
rect 48076 34130 48132 35644
rect 48188 34244 48244 34254
rect 48188 34150 48244 34188
rect 48076 34078 48078 34130
rect 48130 34078 48132 34130
rect 48076 34066 48132 34078
rect 47964 32900 48020 32910
rect 47964 31666 48020 32844
rect 48300 31892 48356 36428
rect 48524 34914 48580 37436
rect 48748 37266 48804 37278
rect 48748 37214 48750 37266
rect 48802 37214 48804 37266
rect 48748 36484 48804 37214
rect 48972 37266 49028 37278
rect 48972 37214 48974 37266
rect 49026 37214 49028 37266
rect 48860 36932 48916 36942
rect 48860 36706 48916 36876
rect 48860 36654 48862 36706
rect 48914 36654 48916 36706
rect 48860 36642 48916 36654
rect 48972 36596 49028 37214
rect 48972 36530 49028 36540
rect 48748 36418 48804 36428
rect 48636 36258 48692 36270
rect 48636 36206 48638 36258
rect 48690 36206 48692 36258
rect 48636 35252 48692 36206
rect 48748 36258 48804 36270
rect 48748 36206 48750 36258
rect 48802 36206 48804 36258
rect 48748 35698 48804 36206
rect 49084 35812 49140 39452
rect 49196 40290 49252 40302
rect 49196 40238 49198 40290
rect 49250 40238 49252 40290
rect 49196 38834 49252 40238
rect 49420 39844 49476 40460
rect 49420 39778 49476 39788
rect 49532 40402 49588 40414
rect 49532 40350 49534 40402
rect 49586 40350 49588 40402
rect 49532 39732 49588 40350
rect 49756 40404 49812 40414
rect 49756 40310 49812 40348
rect 50092 40402 50148 40414
rect 50092 40350 50094 40402
rect 50146 40350 50148 40402
rect 49644 40292 49700 40302
rect 49644 40198 49700 40236
rect 50092 40292 50148 40350
rect 50204 40404 50260 41020
rect 50428 40628 50484 41020
rect 50540 41074 50596 42140
rect 50764 41860 50820 41870
rect 50764 41858 50932 41860
rect 50764 41806 50766 41858
rect 50818 41806 50932 41858
rect 50764 41804 50932 41806
rect 50764 41794 50820 41804
rect 50540 41022 50542 41074
rect 50594 41022 50596 41074
rect 50540 41010 50596 41022
rect 50764 40964 50820 41002
rect 50764 40898 50820 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50876 40628 50932 41804
rect 50988 41186 51044 42476
rect 51548 41636 51604 43260
rect 51660 43222 51716 43260
rect 53788 43316 53844 43326
rect 51660 42644 51716 42654
rect 51660 42550 51716 42588
rect 51996 42642 52052 42654
rect 51996 42590 51998 42642
rect 52050 42590 52052 42642
rect 51772 42530 51828 42542
rect 51772 42478 51774 42530
rect 51826 42478 51828 42530
rect 51772 41970 51828 42478
rect 51772 41918 51774 41970
rect 51826 41918 51828 41970
rect 51772 41906 51828 41918
rect 51884 42084 51940 42094
rect 50988 41134 50990 41186
rect 51042 41134 51044 41186
rect 50988 41122 51044 41134
rect 51212 41580 51604 41636
rect 51660 41858 51716 41870
rect 51660 41806 51662 41858
rect 51714 41806 51716 41858
rect 51212 41186 51268 41580
rect 51212 41134 51214 41186
rect 51266 41134 51268 41186
rect 51212 41122 51268 41134
rect 51324 41412 51380 41422
rect 51324 41186 51380 41356
rect 51324 41134 51326 41186
rect 51378 41134 51380 41186
rect 50428 40572 50596 40628
rect 50204 40338 50260 40348
rect 50316 40402 50372 40414
rect 50316 40350 50318 40402
rect 50370 40350 50372 40402
rect 50092 40226 50148 40236
rect 50316 39956 50372 40350
rect 50204 39844 50260 39854
rect 50092 39788 50204 39844
rect 50092 39732 50148 39788
rect 50204 39778 50260 39788
rect 49532 39666 49588 39676
rect 49868 39676 50148 39732
rect 49308 39620 49364 39630
rect 49308 39526 49364 39564
rect 49756 39620 49812 39630
rect 49756 39526 49812 39564
rect 49868 39618 49924 39676
rect 50316 39620 50372 39900
rect 49868 39566 49870 39618
rect 49922 39566 49924 39618
rect 49868 39554 49924 39566
rect 50092 39618 50372 39620
rect 50092 39566 50318 39618
rect 50370 39566 50372 39618
rect 50092 39564 50372 39566
rect 49644 39508 49700 39518
rect 49644 39414 49700 39452
rect 49196 38782 49198 38834
rect 49250 38782 49252 38834
rect 49196 38770 49252 38782
rect 49644 39060 49700 39070
rect 49644 38834 49700 39004
rect 49756 38948 49812 38958
rect 49756 38854 49812 38892
rect 49644 38782 49646 38834
rect 49698 38782 49700 38834
rect 49644 38050 49700 38782
rect 49644 37998 49646 38050
rect 49698 37998 49700 38050
rect 49644 37986 49700 37998
rect 49420 37266 49476 37278
rect 49420 37214 49422 37266
rect 49474 37214 49476 37266
rect 48748 35646 48750 35698
rect 48802 35646 48804 35698
rect 48748 35634 48804 35646
rect 48860 35756 49140 35812
rect 49196 37154 49252 37166
rect 49196 37102 49198 37154
rect 49250 37102 49252 37154
rect 48748 35476 48804 35486
rect 48748 35382 48804 35420
rect 48636 35196 48804 35252
rect 48524 34862 48526 34914
rect 48578 34862 48580 34914
rect 48524 34356 48580 34862
rect 48748 34804 48804 35196
rect 48748 34738 48804 34748
rect 48524 34290 48580 34300
rect 48748 34132 48804 34142
rect 48860 34132 48916 35756
rect 49196 35700 49252 37102
rect 48972 35644 49252 35700
rect 49420 35700 49476 37214
rect 50092 36820 50148 39564
rect 50316 39554 50372 39564
rect 50428 40180 50484 40190
rect 50428 39060 50484 40124
rect 50540 39844 50596 40572
rect 50652 40572 50932 40628
rect 50652 40180 50708 40572
rect 50988 40516 51044 40526
rect 50988 40422 51044 40460
rect 51324 40516 51380 41134
rect 51436 40626 51492 41580
rect 51436 40574 51438 40626
rect 51490 40574 51492 40626
rect 51436 40562 51492 40574
rect 51660 40626 51716 41806
rect 51772 41412 51828 41422
rect 51884 41412 51940 42028
rect 51996 41748 52052 42590
rect 53004 42084 53060 42094
rect 53004 41990 53060 42028
rect 53788 42082 53844 43260
rect 53788 42030 53790 42082
rect 53842 42030 53844 42082
rect 53788 42018 53844 42030
rect 51996 41682 52052 41692
rect 52220 41972 52276 41982
rect 51772 41410 51940 41412
rect 51772 41358 51774 41410
rect 51826 41358 51940 41410
rect 51772 41356 51940 41358
rect 51772 41346 51828 41356
rect 51884 40964 51940 40974
rect 51940 40908 52052 40964
rect 51884 40898 51940 40908
rect 51660 40574 51662 40626
rect 51714 40574 51716 40626
rect 51660 40562 51716 40574
rect 51996 40626 52052 40908
rect 51996 40574 51998 40626
rect 52050 40574 52052 40626
rect 51996 40562 52052 40574
rect 52220 40626 52276 41916
rect 52780 41970 52836 41982
rect 52780 41918 52782 41970
rect 52834 41918 52836 41970
rect 52780 41748 52836 41918
rect 53676 41972 53732 41982
rect 53676 41878 53732 41916
rect 52780 41682 52836 41692
rect 53564 41858 53620 41870
rect 53564 41806 53566 41858
rect 53618 41806 53620 41858
rect 52220 40574 52222 40626
rect 52274 40574 52276 40626
rect 52220 40562 52276 40574
rect 52556 40628 52612 40638
rect 52556 40534 52612 40572
rect 51324 40422 51380 40460
rect 51884 40516 51940 40526
rect 51884 40422 51940 40460
rect 50764 40404 50820 40414
rect 50764 40310 50820 40348
rect 51660 40404 51716 40414
rect 50876 40292 50932 40302
rect 50876 40198 50932 40236
rect 50652 40114 50708 40124
rect 50988 40068 51044 40078
rect 51044 40012 51156 40068
rect 50988 40002 51044 40012
rect 50652 39844 50708 39854
rect 50540 39788 50652 39844
rect 50652 39618 50708 39788
rect 50652 39566 50654 39618
rect 50706 39566 50708 39618
rect 50652 39554 50708 39566
rect 50988 39394 51044 39406
rect 50988 39342 50990 39394
rect 51042 39342 51044 39394
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50428 38994 50484 39004
rect 50316 38836 50372 38846
rect 50428 38836 50484 38846
rect 50372 38834 50484 38836
rect 50372 38782 50430 38834
rect 50482 38782 50484 38834
rect 50372 38780 50484 38782
rect 50204 37492 50260 37502
rect 50316 37492 50372 38780
rect 50428 38770 50484 38780
rect 50988 38164 51044 39342
rect 51100 38948 51156 40012
rect 51212 39508 51268 39518
rect 51212 39506 51380 39508
rect 51212 39454 51214 39506
rect 51266 39454 51380 39506
rect 51212 39452 51380 39454
rect 51212 39442 51268 39452
rect 51212 38948 51268 38958
rect 51100 38946 51268 38948
rect 51100 38894 51214 38946
rect 51266 38894 51268 38946
rect 51100 38892 51268 38894
rect 51212 38882 51268 38892
rect 51324 38276 51380 39452
rect 51660 39506 51716 40348
rect 51660 39454 51662 39506
rect 51714 39454 51716 39506
rect 51660 38724 51716 39454
rect 51660 38658 51716 38668
rect 53340 38724 53396 38734
rect 53340 38630 53396 38668
rect 51324 38220 51828 38276
rect 50876 38108 51044 38164
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50204 37490 50372 37492
rect 50204 37438 50206 37490
rect 50258 37438 50372 37490
rect 50204 37436 50372 37438
rect 50204 37426 50260 37436
rect 50428 37154 50484 37166
rect 50428 37102 50430 37154
rect 50482 37102 50484 37154
rect 50428 36932 50484 37102
rect 50428 36866 50484 36876
rect 50092 36764 50372 36820
rect 49868 36708 49924 36718
rect 49868 36482 49924 36652
rect 49868 36430 49870 36482
rect 49922 36430 49924 36482
rect 49868 36418 49924 36430
rect 50204 36596 50260 36606
rect 50204 36482 50260 36540
rect 50204 36430 50206 36482
rect 50258 36430 50260 36482
rect 50204 36148 50260 36430
rect 50204 36082 50260 36092
rect 48972 35252 49028 35644
rect 49420 35634 49476 35644
rect 49644 35698 49700 35710
rect 49644 35646 49646 35698
rect 49698 35646 49700 35698
rect 48972 35186 49028 35196
rect 49084 35474 49140 35486
rect 49084 35422 49086 35474
rect 49138 35422 49140 35474
rect 48972 34692 49028 34702
rect 48972 34354 49028 34636
rect 49084 34580 49140 35422
rect 49308 34916 49364 34926
rect 49308 34822 49364 34860
rect 49532 34914 49588 34926
rect 49532 34862 49534 34914
rect 49586 34862 49588 34914
rect 49084 34514 49140 34524
rect 49420 34804 49476 34814
rect 48972 34302 48974 34354
rect 49026 34302 49028 34354
rect 48972 34290 49028 34302
rect 48860 34076 49028 34132
rect 48748 34038 48804 34076
rect 48860 32450 48916 32462
rect 48860 32398 48862 32450
rect 48914 32398 48916 32450
rect 48300 31836 48580 31892
rect 47964 31614 47966 31666
rect 48018 31614 48020 31666
rect 47964 31602 48020 31614
rect 48188 31668 48244 31678
rect 48188 31108 48244 31612
rect 48412 31668 48468 31678
rect 48412 31574 48468 31612
rect 48188 31042 48244 31052
rect 48300 31554 48356 31566
rect 48300 31502 48302 31554
rect 48354 31502 48356 31554
rect 47964 30882 48020 30894
rect 47964 30830 47966 30882
rect 48018 30830 48020 30882
rect 47964 30324 48020 30830
rect 47964 30258 48020 30268
rect 47852 30158 47854 30210
rect 47906 30158 47908 30210
rect 47852 30146 47908 30158
rect 47292 30098 47348 30110
rect 47292 30046 47294 30098
rect 47346 30046 47348 30098
rect 47292 29876 47348 30046
rect 47292 29810 47348 29820
rect 47628 29986 47684 29998
rect 47628 29934 47630 29986
rect 47682 29934 47684 29986
rect 47404 29652 47460 29662
rect 47180 29596 47348 29652
rect 46396 29426 46452 29596
rect 46956 29558 47012 29596
rect 46396 29374 46398 29426
rect 46450 29374 46452 29426
rect 46396 29204 46452 29374
rect 46620 29428 46676 29438
rect 46620 29334 46676 29372
rect 47068 29428 47124 29438
rect 47068 29334 47124 29372
rect 47180 29426 47236 29438
rect 47180 29374 47182 29426
rect 47234 29374 47236 29426
rect 46396 29138 46452 29148
rect 47180 29204 47236 29374
rect 47180 29138 47236 29148
rect 46620 28868 46676 28878
rect 46284 27694 46286 27746
rect 46338 27694 46340 27746
rect 46284 27682 46340 27694
rect 46396 28756 46452 28766
rect 45836 27234 45892 27244
rect 45724 27076 45780 27086
rect 45724 26982 45780 27020
rect 45612 26852 45892 26908
rect 45836 25620 45892 26852
rect 46060 26404 46116 26414
rect 45836 25554 45892 25564
rect 45948 26180 46004 26190
rect 45724 25506 45780 25518
rect 45724 25454 45726 25506
rect 45778 25454 45780 25506
rect 45724 25396 45780 25454
rect 45948 25506 46004 26124
rect 45948 25454 45950 25506
rect 46002 25454 46004 25506
rect 45948 25442 46004 25454
rect 46060 25506 46116 26348
rect 46060 25454 46062 25506
rect 46114 25454 46116 25506
rect 46060 25442 46116 25454
rect 46172 25844 46228 25854
rect 45724 25330 45780 25340
rect 45948 24612 46004 24622
rect 45388 23938 45556 23940
rect 45388 23886 45390 23938
rect 45442 23886 45556 23938
rect 45388 23884 45556 23886
rect 45612 24164 45668 24174
rect 45612 23938 45668 24108
rect 45612 23886 45614 23938
rect 45666 23886 45668 23938
rect 45388 23716 45444 23884
rect 45612 23874 45668 23886
rect 45948 23938 46004 24556
rect 45948 23886 45950 23938
rect 46002 23886 46004 23938
rect 45948 23874 46004 23886
rect 46172 23938 46228 25788
rect 46396 24276 46452 28700
rect 46620 28530 46676 28812
rect 47292 28756 47348 29596
rect 47404 29558 47460 29596
rect 47180 28700 47348 28756
rect 47404 29316 47460 29326
rect 46620 28478 46622 28530
rect 46674 28478 46676 28530
rect 46620 28466 46676 28478
rect 46844 28642 46900 28654
rect 46844 28590 46846 28642
rect 46898 28590 46900 28642
rect 46732 27972 46788 27982
rect 46620 27076 46676 27086
rect 46508 25732 46564 25742
rect 46620 25732 46676 27020
rect 46732 26514 46788 27916
rect 46732 26462 46734 26514
rect 46786 26462 46788 26514
rect 46732 26404 46788 26462
rect 46732 26338 46788 26348
rect 46844 26292 46900 28590
rect 46956 28420 47012 28430
rect 46956 28326 47012 28364
rect 46844 26226 46900 26236
rect 46508 25730 46676 25732
rect 46508 25678 46510 25730
rect 46562 25678 46676 25730
rect 46508 25676 46676 25678
rect 46508 25666 46564 25676
rect 46956 25620 47012 25630
rect 46956 25526 47012 25564
rect 47180 25284 47236 28700
rect 47292 28532 47348 28542
rect 47292 28438 47348 28476
rect 47404 27188 47460 29260
rect 47628 28868 47684 29934
rect 48076 29988 48132 29998
rect 48076 29894 48132 29932
rect 48300 29316 48356 31502
rect 48524 31556 48580 31836
rect 48748 31556 48804 31566
rect 48524 31554 48804 31556
rect 48524 31502 48750 31554
rect 48802 31502 48804 31554
rect 48524 31500 48804 31502
rect 48748 30212 48804 31500
rect 48860 31332 48916 32398
rect 48860 31266 48916 31276
rect 48748 30146 48804 30156
rect 48860 30100 48916 30110
rect 48972 30100 49028 34076
rect 49196 34130 49252 34142
rect 49196 34078 49198 34130
rect 49250 34078 49252 34130
rect 49084 34018 49140 34030
rect 49084 33966 49086 34018
rect 49138 33966 49140 34018
rect 49084 32900 49140 33966
rect 49084 32834 49140 32844
rect 49196 33124 49252 34078
rect 49420 34130 49476 34748
rect 49420 34078 49422 34130
rect 49474 34078 49476 34130
rect 49420 34020 49476 34078
rect 49420 33954 49476 33964
rect 49196 32788 49252 33068
rect 49532 32900 49588 34862
rect 49644 34244 49700 35646
rect 49980 35700 50036 35710
rect 49644 34178 49700 34188
rect 49756 34580 49812 34590
rect 49756 34020 49812 34524
rect 49980 34354 50036 35644
rect 49980 34302 49982 34354
rect 50034 34302 50036 34354
rect 49868 34020 49924 34030
rect 49756 34018 49924 34020
rect 49756 33966 49870 34018
rect 49922 33966 49924 34018
rect 49756 33964 49924 33966
rect 49868 33954 49924 33964
rect 49980 33346 50036 34302
rect 50092 34804 50148 34814
rect 50092 33570 50148 34748
rect 50204 34244 50260 34254
rect 50204 34150 50260 34188
rect 50092 33518 50094 33570
rect 50146 33518 50148 33570
rect 50092 33506 50148 33518
rect 50204 33908 50260 33918
rect 49980 33294 49982 33346
rect 50034 33294 50036 33346
rect 49980 33282 50036 33294
rect 50204 32900 50260 33852
rect 49196 32722 49252 32732
rect 49308 32844 49588 32900
rect 50092 32844 50260 32900
rect 49308 32564 49364 32844
rect 50092 32676 50148 32844
rect 49868 32674 50148 32676
rect 49868 32622 50094 32674
rect 50146 32622 50148 32674
rect 49868 32620 50148 32622
rect 49084 32562 49364 32564
rect 49084 32510 49310 32562
rect 49362 32510 49364 32562
rect 49084 32508 49364 32510
rect 49084 31778 49140 32508
rect 49308 32498 49364 32508
rect 49532 32564 49588 32574
rect 49084 31726 49086 31778
rect 49138 31726 49140 31778
rect 49084 31556 49140 31726
rect 49084 31490 49140 31500
rect 49420 31220 49476 31230
rect 49420 31126 49476 31164
rect 49196 30994 49252 31006
rect 49196 30942 49198 30994
rect 49250 30942 49252 30994
rect 49196 30436 49252 30942
rect 49420 30994 49476 31006
rect 49420 30942 49422 30994
rect 49474 30942 49476 30994
rect 49420 30884 49476 30942
rect 49420 30818 49476 30828
rect 49532 30436 49588 32508
rect 49756 32564 49812 32574
rect 49756 32470 49812 32508
rect 49756 32340 49812 32350
rect 49644 32284 49756 32340
rect 49644 30660 49700 32284
rect 49756 32274 49812 32284
rect 49756 31554 49812 31566
rect 49756 31502 49758 31554
rect 49810 31502 49812 31554
rect 49756 31332 49812 31502
rect 49756 31266 49812 31276
rect 49756 30996 49812 31006
rect 49868 30996 49924 32620
rect 50092 32610 50148 32620
rect 50204 32674 50260 32686
rect 50204 32622 50206 32674
rect 50258 32622 50260 32674
rect 50204 32564 50260 32622
rect 50204 32498 50260 32508
rect 50204 32338 50260 32350
rect 50204 32286 50206 32338
rect 50258 32286 50260 32338
rect 49756 30994 49924 30996
rect 49756 30942 49758 30994
rect 49810 30942 49924 30994
rect 49756 30940 49924 30942
rect 49756 30930 49812 30940
rect 49868 30660 49924 30940
rect 49980 31554 50036 31566
rect 49980 31502 49982 31554
rect 50034 31502 50036 31554
rect 49980 30772 50036 31502
rect 50092 31554 50148 31566
rect 50092 31502 50094 31554
rect 50146 31502 50148 31554
rect 50092 30994 50148 31502
rect 50204 31556 50260 32286
rect 50316 32340 50372 36764
rect 50876 36596 50932 38108
rect 51324 38052 51380 38062
rect 51212 38050 51380 38052
rect 51212 37998 51326 38050
rect 51378 37998 51380 38050
rect 51212 37996 51380 37998
rect 50988 37940 51044 37950
rect 50988 37490 51044 37884
rect 50988 37438 50990 37490
rect 51042 37438 51044 37490
rect 50988 37426 51044 37438
rect 51100 37828 51156 37838
rect 51100 37268 51156 37772
rect 51100 37202 51156 37212
rect 50428 36540 50932 36596
rect 50428 35924 50484 36540
rect 50876 36370 50932 36382
rect 50876 36318 50878 36370
rect 50930 36318 50932 36370
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50764 35924 50820 35934
rect 50428 35868 50596 35924
rect 50428 35586 50484 35598
rect 50428 35534 50430 35586
rect 50482 35534 50484 35586
rect 50428 34916 50484 35534
rect 50428 34850 50484 34860
rect 50540 34692 50596 35868
rect 50764 35700 50820 35868
rect 50876 35700 50932 36318
rect 51212 35924 51268 37996
rect 51324 37986 51380 37996
rect 51324 37156 51380 37166
rect 51436 37156 51492 38220
rect 51772 38052 51828 38220
rect 51772 37958 51828 37996
rect 52780 38052 52836 38062
rect 52556 37940 52612 37950
rect 52556 37268 52612 37884
rect 52780 37938 52836 37996
rect 52780 37886 52782 37938
rect 52834 37886 52836 37938
rect 52780 37874 52836 37886
rect 52892 38050 52948 38062
rect 52892 37998 52894 38050
rect 52946 37998 52948 38050
rect 52556 37212 52836 37268
rect 51324 37154 51492 37156
rect 51324 37102 51326 37154
rect 51378 37102 51492 37154
rect 51324 37100 51492 37102
rect 51324 37090 51380 37100
rect 52556 36932 52612 36942
rect 51660 36820 51716 36830
rect 51660 36594 51716 36764
rect 51660 36542 51662 36594
rect 51714 36542 51716 36594
rect 51660 36530 51716 36542
rect 52332 36820 52388 36830
rect 52108 36260 52164 36270
rect 52108 36166 52164 36204
rect 51212 35858 51268 35868
rect 51436 35700 51492 35710
rect 50876 35698 51492 35700
rect 50876 35646 51438 35698
rect 51490 35646 51492 35698
rect 50876 35644 51492 35646
rect 50764 35606 50820 35644
rect 50988 34914 51044 35644
rect 51436 35634 51492 35644
rect 51548 35364 51604 35374
rect 51548 35138 51604 35308
rect 51548 35086 51550 35138
rect 51602 35086 51604 35138
rect 51548 35074 51604 35086
rect 50988 34862 50990 34914
rect 51042 34862 51044 34914
rect 50988 34850 51044 34862
rect 51100 35026 51156 35038
rect 51100 34974 51102 35026
rect 51154 34974 51156 35026
rect 51100 34804 51156 34974
rect 51100 34738 51156 34748
rect 51772 34916 51828 34926
rect 50428 34636 50596 34692
rect 50428 34132 50484 34636
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 51660 34356 51716 34366
rect 50652 34244 50708 34254
rect 50652 34150 50708 34188
rect 50428 34066 50484 34076
rect 51100 34132 51156 34142
rect 50988 33796 51044 33806
rect 50876 33348 50932 33358
rect 50876 33254 50932 33292
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50764 32564 50820 32574
rect 50764 32470 50820 32508
rect 50316 32274 50372 32284
rect 50988 32228 51044 33740
rect 51100 33346 51156 34076
rect 51660 34020 51716 34300
rect 51772 34130 51828 34860
rect 52332 34916 52388 36764
rect 52556 35698 52612 36876
rect 52668 36482 52724 36494
rect 52668 36430 52670 36482
rect 52722 36430 52724 36482
rect 52668 36372 52724 36430
rect 52668 36306 52724 36316
rect 52556 35646 52558 35698
rect 52610 35646 52612 35698
rect 52556 35634 52612 35646
rect 52332 34850 52388 34860
rect 52668 35140 52724 35150
rect 52668 34914 52724 35084
rect 52668 34862 52670 34914
rect 52722 34862 52724 34914
rect 52668 34850 52724 34862
rect 52780 34916 52836 37212
rect 52892 36708 52948 37998
rect 53564 38052 53620 41806
rect 55020 38162 55076 38174
rect 55020 38110 55022 38162
rect 55074 38110 55076 38162
rect 53564 37986 53620 37996
rect 54572 38052 54628 38062
rect 54572 37958 54628 37996
rect 53340 37938 53396 37950
rect 53340 37886 53342 37938
rect 53394 37886 53396 37938
rect 53340 37380 53396 37886
rect 53340 37324 53620 37380
rect 52892 36642 52948 36652
rect 53452 37154 53508 37166
rect 53452 37102 53454 37154
rect 53506 37102 53508 37154
rect 52892 36370 52948 36382
rect 52892 36318 52894 36370
rect 52946 36318 52948 36370
rect 52892 35924 52948 36318
rect 52892 35858 52948 35868
rect 53116 36258 53172 36270
rect 53116 36206 53118 36258
rect 53170 36206 53172 36258
rect 52892 35252 52948 35262
rect 52892 35138 52948 35196
rect 52892 35086 52894 35138
rect 52946 35086 52948 35138
rect 52892 35074 52948 35086
rect 52780 34860 53060 34916
rect 51772 34078 51774 34130
rect 51826 34078 51828 34130
rect 51772 34066 51828 34078
rect 51212 33908 51268 33946
rect 51212 33842 51268 33852
rect 51212 33684 51268 33694
rect 51212 33458 51268 33628
rect 51212 33406 51214 33458
rect 51266 33406 51268 33458
rect 51212 33394 51268 33406
rect 51660 33458 51716 33964
rect 51660 33406 51662 33458
rect 51714 33406 51716 33458
rect 51660 33394 51716 33406
rect 51100 33294 51102 33346
rect 51154 33294 51156 33346
rect 51100 33282 51156 33294
rect 52108 33236 52164 33246
rect 52108 33142 52164 33180
rect 53004 33234 53060 34860
rect 53116 34130 53172 36206
rect 53340 35586 53396 35598
rect 53340 35534 53342 35586
rect 53394 35534 53396 35586
rect 53340 35252 53396 35534
rect 53340 35186 53396 35196
rect 53340 35028 53396 35038
rect 53452 35028 53508 37102
rect 53340 35026 53508 35028
rect 53340 34974 53342 35026
rect 53394 34974 53508 35026
rect 53340 34972 53508 34974
rect 53564 37044 53620 37324
rect 54124 37268 54180 37278
rect 54124 37174 54180 37212
rect 55020 37266 55076 38110
rect 56140 37380 56196 37390
rect 56140 37378 56868 37380
rect 56140 37326 56142 37378
rect 56194 37326 56868 37378
rect 56140 37324 56868 37326
rect 56140 37314 56196 37324
rect 55020 37214 55022 37266
rect 55074 37214 55076 37266
rect 53340 34962 53396 34972
rect 53228 34804 53284 34814
rect 53228 34710 53284 34748
rect 53452 34804 53508 34814
rect 53452 34710 53508 34748
rect 53564 34580 53620 36988
rect 54572 37154 54628 37166
rect 54572 37102 54574 37154
rect 54626 37102 54628 37154
rect 54572 36708 54628 37102
rect 54796 37044 54852 37054
rect 54572 36642 54628 36652
rect 54684 36932 54740 36942
rect 54684 36594 54740 36876
rect 54684 36542 54686 36594
rect 54738 36542 54740 36594
rect 54012 36484 54068 36494
rect 54012 36258 54068 36428
rect 54124 36482 54180 36494
rect 54124 36430 54126 36482
rect 54178 36430 54180 36482
rect 54124 36372 54180 36430
rect 54572 36484 54628 36494
rect 54124 36306 54180 36316
rect 54460 36372 54516 36382
rect 54012 36206 54014 36258
rect 54066 36206 54068 36258
rect 54012 36194 54068 36206
rect 54236 36260 54292 36270
rect 53116 34078 53118 34130
rect 53170 34078 53172 34130
rect 53116 34066 53172 34078
rect 53452 34524 53620 34580
rect 53676 35252 53732 35262
rect 53452 33348 53508 34524
rect 53676 34356 53732 35196
rect 53676 34290 53732 34300
rect 54124 35026 54180 35038
rect 54124 34974 54126 35026
rect 54178 34974 54180 35026
rect 53564 34132 53620 34142
rect 53564 34130 53844 34132
rect 53564 34078 53566 34130
rect 53618 34078 53844 34130
rect 53564 34076 53844 34078
rect 53564 34066 53620 34076
rect 53564 33348 53620 33358
rect 53452 33346 53620 33348
rect 53452 33294 53566 33346
rect 53618 33294 53620 33346
rect 53452 33292 53620 33294
rect 53004 33182 53006 33234
rect 53058 33182 53060 33234
rect 53004 33170 53060 33182
rect 53564 33236 53620 33292
rect 53564 33170 53620 33180
rect 52220 32788 52276 32798
rect 52220 32694 52276 32732
rect 51660 32676 51716 32686
rect 51660 32582 51716 32620
rect 52780 32674 52836 32686
rect 52780 32622 52782 32674
rect 52834 32622 52836 32674
rect 51772 32564 51828 32574
rect 51772 32470 51828 32508
rect 52108 32562 52164 32574
rect 52108 32510 52110 32562
rect 52162 32510 52164 32562
rect 51324 32452 51380 32462
rect 51324 32450 51604 32452
rect 51324 32398 51326 32450
rect 51378 32398 51604 32450
rect 51324 32396 51604 32398
rect 51324 32386 51380 32396
rect 50988 32162 51044 32172
rect 50988 32002 51044 32014
rect 50988 31950 50990 32002
rect 51042 31950 51044 32002
rect 50988 31948 51044 31950
rect 50876 31892 51044 31948
rect 51324 32004 51380 32014
rect 50204 31554 50372 31556
rect 50204 31502 50206 31554
rect 50258 31502 50372 31554
rect 50204 31500 50372 31502
rect 50204 31490 50260 31500
rect 50316 31108 50372 31500
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50540 31108 50596 31118
rect 50316 31106 50596 31108
rect 50316 31054 50542 31106
rect 50594 31054 50596 31106
rect 50316 31052 50596 31054
rect 50540 31042 50596 31052
rect 50092 30942 50094 30994
rect 50146 30942 50148 30994
rect 50092 30930 50148 30942
rect 50204 30994 50260 31006
rect 50204 30942 50206 30994
rect 50258 30942 50260 30994
rect 50204 30884 50260 30942
rect 50204 30772 50260 30828
rect 50428 30884 50484 30894
rect 50876 30884 50932 31892
rect 50428 30882 50932 30884
rect 50428 30830 50430 30882
rect 50482 30830 50932 30882
rect 50428 30828 50932 30830
rect 50988 31778 51044 31790
rect 50988 31726 50990 31778
rect 51042 31726 51044 31778
rect 50988 30882 51044 31726
rect 51324 31778 51380 31948
rect 51324 31726 51326 31778
rect 51378 31726 51380 31778
rect 51324 31714 51380 31726
rect 51548 31666 51604 32396
rect 51996 32004 52052 32014
rect 52108 31948 52164 32510
rect 51548 31614 51550 31666
rect 51602 31614 51604 31666
rect 51436 31556 51492 31566
rect 51436 31462 51492 31500
rect 50988 30830 50990 30882
rect 51042 30830 51044 30882
rect 50428 30818 50484 30828
rect 49980 30716 50260 30772
rect 50204 30660 50260 30716
rect 50988 30660 51044 30830
rect 49644 30604 49812 30660
rect 49868 30604 50148 30660
rect 50204 30604 50484 30660
rect 49756 30548 49812 30604
rect 49756 30492 49924 30548
rect 49532 30380 49812 30436
rect 49196 30370 49252 30380
rect 49532 30212 49588 30222
rect 48860 30098 49028 30100
rect 48860 30046 48862 30098
rect 48914 30046 49028 30098
rect 48860 30044 49028 30046
rect 48860 30034 48916 30044
rect 48524 29988 48580 29998
rect 48524 29894 48580 29932
rect 48300 29250 48356 29260
rect 48972 29204 49028 30044
rect 49084 30210 49588 30212
rect 49084 30158 49534 30210
rect 49586 30158 49588 30210
rect 49084 30156 49588 30158
rect 49084 29426 49140 30156
rect 49532 30146 49588 30156
rect 49420 29988 49476 29998
rect 49420 29894 49476 29932
rect 49644 29988 49700 29998
rect 49644 29894 49700 29932
rect 49308 29650 49364 29662
rect 49308 29598 49310 29650
rect 49362 29598 49364 29650
rect 49084 29374 49086 29426
rect 49138 29374 49140 29426
rect 49084 29362 49140 29374
rect 49196 29426 49252 29438
rect 49196 29374 49198 29426
rect 49250 29374 49252 29426
rect 49196 29204 49252 29374
rect 48972 29148 49252 29204
rect 47404 27094 47460 27132
rect 47516 28812 47684 28868
rect 47516 25844 47572 28812
rect 49308 28754 49364 29598
rect 49532 29428 49588 29438
rect 49308 28702 49310 28754
rect 49362 28702 49364 28754
rect 49308 28690 49364 28702
rect 49420 29426 49588 29428
rect 49420 29374 49534 29426
rect 49586 29374 49588 29426
rect 49420 29372 49588 29374
rect 49756 29428 49812 30380
rect 49868 30098 49924 30492
rect 49868 30046 49870 30098
rect 49922 30046 49924 30098
rect 49868 29652 49924 30046
rect 49868 29586 49924 29596
rect 49756 29372 49924 29428
rect 47628 28644 47684 28654
rect 47628 28642 47796 28644
rect 47628 28590 47630 28642
rect 47682 28590 47796 28642
rect 47628 28588 47796 28590
rect 47628 28578 47684 28588
rect 47740 28082 47796 28588
rect 48524 28642 48580 28654
rect 48524 28590 48526 28642
rect 48578 28590 48580 28642
rect 47740 28030 47742 28082
rect 47794 28030 47796 28082
rect 47740 28018 47796 28030
rect 48188 28420 48244 28430
rect 48524 28420 48580 28590
rect 48188 28418 48580 28420
rect 48188 28366 48190 28418
rect 48242 28366 48580 28418
rect 48188 28364 48580 28366
rect 47852 27860 47908 27870
rect 47852 26628 47908 27804
rect 48188 27188 48244 28364
rect 48860 28308 48916 28318
rect 48860 28082 48916 28252
rect 48860 28030 48862 28082
rect 48914 28030 48916 28082
rect 48860 28018 48916 28030
rect 48972 27860 49028 27870
rect 48972 27858 49364 27860
rect 48972 27806 48974 27858
rect 49026 27806 49364 27858
rect 48972 27804 49364 27806
rect 48972 27794 49028 27804
rect 49084 27636 49140 27646
rect 48188 26740 48244 27132
rect 48972 27634 49140 27636
rect 48972 27582 49086 27634
rect 49138 27582 49140 27634
rect 48972 27580 49140 27582
rect 48748 27076 48804 27114
rect 48748 27010 48804 27020
rect 48972 26908 49028 27580
rect 49084 27570 49140 27580
rect 49196 27636 49252 27646
rect 48524 26852 48580 26862
rect 48972 26852 49140 26908
rect 48524 26758 48580 26796
rect 48188 26684 48468 26740
rect 47852 26572 48244 26628
rect 47628 26404 47684 26414
rect 47628 26310 47684 26348
rect 48188 26290 48244 26572
rect 48188 26238 48190 26290
rect 48242 26238 48244 26290
rect 48188 26226 48244 26238
rect 47516 25778 47572 25788
rect 47292 25618 47348 25630
rect 47292 25566 47294 25618
rect 47346 25566 47348 25618
rect 47292 25508 47348 25566
rect 47516 25620 47572 25630
rect 47292 25442 47348 25452
rect 47404 25506 47460 25518
rect 47404 25454 47406 25506
rect 47458 25454 47460 25506
rect 47068 25228 47236 25284
rect 46508 24724 46564 24734
rect 46508 24630 46564 24668
rect 46732 24612 46788 24622
rect 46172 23886 46174 23938
rect 46226 23886 46228 23938
rect 46172 23874 46228 23886
rect 46284 24220 46452 24276
rect 46620 24610 46788 24612
rect 46620 24558 46734 24610
rect 46786 24558 46788 24610
rect 46620 24556 46788 24558
rect 45388 23650 45444 23660
rect 45500 23714 45556 23726
rect 45500 23662 45502 23714
rect 45554 23662 45556 23714
rect 45388 23156 45444 23166
rect 45276 23100 45388 23156
rect 45388 23062 45444 23100
rect 44828 22708 44884 22718
rect 44828 22594 44884 22652
rect 44828 22542 44830 22594
rect 44882 22542 44884 22594
rect 44828 22530 44884 22542
rect 45500 22484 45556 23662
rect 46284 23492 46340 24220
rect 46396 24052 46452 24062
rect 46396 23714 46452 23996
rect 46508 23828 46564 23838
rect 46508 23734 46564 23772
rect 46396 23662 46398 23714
rect 46450 23662 46452 23714
rect 46396 23650 46452 23662
rect 46284 23436 46452 23492
rect 46060 23268 46116 23278
rect 46060 23174 46116 23212
rect 46396 23268 46452 23436
rect 46508 23268 46564 23278
rect 46396 23266 46564 23268
rect 46396 23214 46510 23266
rect 46562 23214 46564 23266
rect 46396 23212 46564 23214
rect 46284 23154 46340 23166
rect 46284 23102 46286 23154
rect 46338 23102 46340 23154
rect 46172 23042 46228 23054
rect 46172 22990 46174 23042
rect 46226 22990 46228 23042
rect 46060 22596 46116 22606
rect 45500 22428 45668 22484
rect 44268 22194 44324 22204
rect 45276 22260 45332 22270
rect 45276 22166 45332 22204
rect 45388 22258 45444 22270
rect 45388 22206 45390 22258
rect 45442 22206 45444 22258
rect 43932 21382 43988 21420
rect 44044 22148 44100 22158
rect 41580 20750 41582 20802
rect 41634 20750 41636 20802
rect 41580 20738 41636 20750
rect 41692 20802 42084 20804
rect 41692 20750 42030 20802
rect 42082 20750 42084 20802
rect 41692 20748 42084 20750
rect 41580 20580 41636 20590
rect 41580 20486 41636 20524
rect 41580 20132 41636 20142
rect 41468 20130 41636 20132
rect 41468 20078 41582 20130
rect 41634 20078 41636 20130
rect 41468 20076 41636 20078
rect 41580 20066 41636 20076
rect 41692 20130 41748 20748
rect 42028 20738 42084 20748
rect 42364 20914 42980 20916
rect 42364 20862 42814 20914
rect 42866 20862 42980 20914
rect 42364 20860 42980 20862
rect 44044 20914 44100 22092
rect 45388 22148 45444 22206
rect 45500 22260 45556 22270
rect 45500 22166 45556 22204
rect 45388 22082 45444 22092
rect 44044 20862 44046 20914
rect 44098 20862 44100 20914
rect 42364 20802 42420 20860
rect 42812 20850 42868 20860
rect 44044 20850 44100 20862
rect 44268 21364 44324 21374
rect 44268 20914 44324 21308
rect 44268 20862 44270 20914
rect 44322 20862 44324 20914
rect 44268 20850 44324 20862
rect 44940 20916 44996 20926
rect 42364 20750 42366 20802
rect 42418 20750 42420 20802
rect 42364 20738 42420 20750
rect 44940 20802 44996 20860
rect 45612 20914 45668 22428
rect 46060 22372 46116 22540
rect 46060 22306 46116 22316
rect 46060 22148 46116 22158
rect 46060 21698 46116 22092
rect 46060 21646 46062 21698
rect 46114 21646 46116 21698
rect 46060 21634 46116 21646
rect 46172 21700 46228 22990
rect 46284 22932 46340 23102
rect 46284 22866 46340 22876
rect 46172 21634 46228 21644
rect 45612 20862 45614 20914
rect 45666 20862 45668 20914
rect 45612 20850 45668 20862
rect 44940 20750 44942 20802
rect 44994 20750 44996 20802
rect 44940 20738 44996 20750
rect 45836 20244 45892 20254
rect 46396 20244 46452 23212
rect 46508 23202 46564 23212
rect 46508 22484 46564 22494
rect 46620 22484 46676 24556
rect 46732 24546 46788 24556
rect 46732 24276 46788 24286
rect 46732 23938 46788 24220
rect 47068 24052 47124 25228
rect 47180 25060 47236 25070
rect 47180 24834 47236 25004
rect 47180 24782 47182 24834
rect 47234 24782 47236 24834
rect 47180 24770 47236 24782
rect 47180 24276 47236 24286
rect 47180 24162 47236 24220
rect 47180 24110 47182 24162
rect 47234 24110 47236 24162
rect 47180 24098 47236 24110
rect 47068 23986 47124 23996
rect 47292 24052 47348 24062
rect 46732 23886 46734 23938
rect 46786 23886 46788 23938
rect 46732 23874 46788 23886
rect 46564 22428 46676 22484
rect 47068 23492 47124 23502
rect 47068 23154 47124 23436
rect 47068 23102 47070 23154
rect 47122 23102 47124 23154
rect 47068 22484 47124 23102
rect 47292 22820 47348 23996
rect 47404 23940 47460 25454
rect 47516 24834 47572 25564
rect 47516 24782 47518 24834
rect 47570 24782 47572 24834
rect 47516 24770 47572 24782
rect 47628 25506 47684 25518
rect 47628 25454 47630 25506
rect 47682 25454 47684 25506
rect 47628 24276 47684 25454
rect 47628 24210 47684 24220
rect 47740 25284 47796 25294
rect 47740 24052 47796 25228
rect 47852 24722 47908 24734
rect 47852 24670 47854 24722
rect 47906 24670 47908 24722
rect 47852 24388 47908 24670
rect 48188 24722 48244 24734
rect 48188 24670 48190 24722
rect 48242 24670 48244 24722
rect 47964 24612 48020 24622
rect 47964 24518 48020 24556
rect 48188 24500 48244 24670
rect 48412 24612 48468 26684
rect 48636 26516 48692 26526
rect 48524 26460 48636 26516
rect 48524 25172 48580 26460
rect 48636 26450 48692 26460
rect 48860 26516 48916 26526
rect 48860 26422 48916 26460
rect 48972 26292 49028 26302
rect 48524 25116 48804 25172
rect 48636 24612 48692 24622
rect 48412 24556 48636 24612
rect 48636 24546 48692 24556
rect 48188 24434 48244 24444
rect 47908 24332 48132 24388
rect 47852 24322 47908 24332
rect 47740 23996 47908 24052
rect 47404 23042 47460 23884
rect 47628 23826 47684 23838
rect 47628 23774 47630 23826
rect 47682 23774 47684 23826
rect 47628 23492 47684 23774
rect 47628 23426 47684 23436
rect 47740 23826 47796 23838
rect 47740 23774 47742 23826
rect 47794 23774 47796 23826
rect 47404 22990 47406 23042
rect 47458 22990 47460 23042
rect 47404 22978 47460 22990
rect 47516 23268 47572 23278
rect 47740 23268 47796 23774
rect 47516 23266 47796 23268
rect 47516 23214 47518 23266
rect 47570 23214 47796 23266
rect 47516 23212 47796 23214
rect 47292 22764 47460 22820
rect 46508 22390 46564 22428
rect 47068 22418 47124 22428
rect 47292 21700 47348 21710
rect 46844 21586 46900 21598
rect 46844 21534 46846 21586
rect 46898 21534 46900 21586
rect 46844 20916 46900 21534
rect 47292 21586 47348 21644
rect 47404 21698 47460 22764
rect 47516 22370 47572 23212
rect 47852 23044 47908 23996
rect 47740 22988 47908 23044
rect 47964 23938 48020 23950
rect 47964 23886 47966 23938
rect 48018 23886 48020 23938
rect 47964 23492 48020 23886
rect 47964 23154 48020 23436
rect 47964 23102 47966 23154
rect 48018 23102 48020 23154
rect 47516 22318 47518 22370
rect 47570 22318 47572 22370
rect 47516 22036 47572 22318
rect 47516 21970 47572 21980
rect 47628 22372 47684 22382
rect 47628 21810 47684 22316
rect 47628 21758 47630 21810
rect 47682 21758 47684 21810
rect 47628 21746 47684 21758
rect 47404 21646 47406 21698
rect 47458 21646 47460 21698
rect 47404 21634 47460 21646
rect 47292 21534 47294 21586
rect 47346 21534 47348 21586
rect 47292 21522 47348 21534
rect 47740 21588 47796 22988
rect 47852 22484 47908 22494
rect 47852 22370 47908 22428
rect 47852 22318 47854 22370
rect 47906 22318 47908 22370
rect 47852 22306 47908 22318
rect 47964 22260 48020 23102
rect 48076 22482 48132 24332
rect 48748 23826 48804 25116
rect 48972 24834 49028 26236
rect 48972 24782 48974 24834
rect 49026 24782 49028 24834
rect 48972 24770 49028 24782
rect 49084 24724 49140 26852
rect 49196 25732 49252 27580
rect 49308 26180 49364 27804
rect 49420 26402 49476 29372
rect 49532 29362 49588 29372
rect 49644 29316 49700 29326
rect 49532 28308 49588 28318
rect 49532 28082 49588 28252
rect 49532 28030 49534 28082
rect 49586 28030 49588 28082
rect 49532 28018 49588 28030
rect 49644 27074 49700 29260
rect 49644 27022 49646 27074
rect 49698 27022 49700 27074
rect 49644 27010 49700 27022
rect 49756 29204 49812 29214
rect 49756 26962 49812 29148
rect 49756 26910 49758 26962
rect 49810 26910 49812 26962
rect 49756 26898 49812 26910
rect 49868 26908 49924 29372
rect 50092 29426 50148 30604
rect 50092 29374 50094 29426
rect 50146 29374 50148 29426
rect 50092 29362 50148 29374
rect 50204 29876 50260 29886
rect 49980 28532 50036 28542
rect 49980 27970 50036 28476
rect 49980 27918 49982 27970
rect 50034 27918 50036 27970
rect 49980 27636 50036 27918
rect 49980 27570 50036 27580
rect 49868 26852 50036 26908
rect 49420 26350 49422 26402
rect 49474 26350 49476 26402
rect 49420 26338 49476 26350
rect 49868 26740 49924 26750
rect 49532 26290 49588 26302
rect 49868 26292 49924 26684
rect 49532 26238 49534 26290
rect 49586 26238 49588 26290
rect 49532 26180 49588 26238
rect 49308 26124 49588 26180
rect 49756 26290 49924 26292
rect 49756 26238 49870 26290
rect 49922 26238 49924 26290
rect 49756 26236 49924 26238
rect 49196 25676 49364 25732
rect 49196 25506 49252 25518
rect 49196 25454 49198 25506
rect 49250 25454 49252 25506
rect 49196 25060 49252 25454
rect 49196 24994 49252 25004
rect 49084 24658 49140 24668
rect 49196 24724 49252 24734
rect 49308 24724 49364 25676
rect 49196 24722 49364 24724
rect 49196 24670 49198 24722
rect 49250 24670 49364 24722
rect 49196 24668 49364 24670
rect 49420 25060 49476 25070
rect 49196 24658 49252 24668
rect 49084 24500 49140 24510
rect 48748 23774 48750 23826
rect 48802 23774 48804 23826
rect 48748 23762 48804 23774
rect 48972 23828 49028 23838
rect 48300 23714 48356 23726
rect 48300 23662 48302 23714
rect 48354 23662 48356 23714
rect 48076 22430 48078 22482
rect 48130 22430 48132 22482
rect 48076 22418 48132 22430
rect 48188 23604 48244 23614
rect 48300 23604 48356 23662
rect 48244 23548 48356 23604
rect 48412 23714 48468 23726
rect 48412 23662 48414 23714
rect 48466 23662 48468 23714
rect 47964 22194 48020 22204
rect 46844 20850 46900 20860
rect 47180 20916 47236 20926
rect 45836 20242 46452 20244
rect 45836 20190 45838 20242
rect 45890 20190 46452 20242
rect 45836 20188 46452 20190
rect 47180 20242 47236 20860
rect 47740 20914 47796 21532
rect 47852 21812 47908 21822
rect 47852 21586 47908 21756
rect 47852 21534 47854 21586
rect 47906 21534 47908 21586
rect 47852 21522 47908 21534
rect 47740 20862 47742 20914
rect 47794 20862 47796 20914
rect 47740 20850 47796 20862
rect 48188 20916 48244 23548
rect 48412 23156 48468 23662
rect 48524 23714 48580 23726
rect 48524 23662 48526 23714
rect 48578 23662 48580 23714
rect 48524 23492 48580 23662
rect 48524 23426 48580 23436
rect 48972 23492 49028 23772
rect 49084 23492 49140 24444
rect 49420 24500 49476 25004
rect 49532 24948 49588 24958
rect 49532 24854 49588 24892
rect 49532 24724 49588 24734
rect 49532 24630 49588 24668
rect 49420 24498 49588 24500
rect 49420 24446 49422 24498
rect 49474 24446 49588 24498
rect 49420 24444 49588 24446
rect 49420 24434 49476 24444
rect 49196 24276 49252 24286
rect 49196 24162 49252 24220
rect 49196 24110 49198 24162
rect 49250 24110 49252 24162
rect 49196 24098 49252 24110
rect 49420 23940 49476 23950
rect 49308 23828 49364 23838
rect 49308 23714 49364 23772
rect 49420 23826 49476 23884
rect 49420 23774 49422 23826
rect 49474 23774 49476 23826
rect 49420 23762 49476 23774
rect 49532 23828 49588 24444
rect 49644 23828 49700 23838
rect 49532 23772 49644 23828
rect 49644 23762 49700 23772
rect 49308 23662 49310 23714
rect 49362 23662 49364 23714
rect 49308 23650 49364 23662
rect 49532 23604 49588 23614
rect 49084 23436 49252 23492
rect 48972 23426 49028 23436
rect 49196 23378 49252 23436
rect 49196 23326 49198 23378
rect 49250 23326 49252 23378
rect 49196 23314 49252 23326
rect 48636 23268 48692 23278
rect 48636 23156 48692 23212
rect 48412 23100 48580 23156
rect 48524 22932 48580 23100
rect 48636 23154 48916 23156
rect 48636 23102 48638 23154
rect 48690 23102 48916 23154
rect 48636 23100 48916 23102
rect 48636 23090 48692 23100
rect 48524 22876 48804 22932
rect 48748 22594 48804 22876
rect 48748 22542 48750 22594
rect 48802 22542 48804 22594
rect 48748 22530 48804 22542
rect 48860 22484 48916 23100
rect 49084 23154 49140 23166
rect 49084 23102 49086 23154
rect 49138 23102 49140 23154
rect 49084 22932 49140 23102
rect 49308 23156 49364 23166
rect 49308 23062 49364 23100
rect 49084 22866 49140 22876
rect 48860 22418 48916 22428
rect 48412 22372 48468 22382
rect 48412 22278 48468 22316
rect 49420 22260 49476 22270
rect 49420 22166 49476 22204
rect 48636 22148 48692 22158
rect 48636 22054 48692 22092
rect 49084 22146 49140 22158
rect 49084 22094 49086 22146
rect 49138 22094 49140 22146
rect 48748 22036 48804 22046
rect 48748 21810 48804 21980
rect 48748 21758 48750 21810
rect 48802 21758 48804 21810
rect 48748 21746 48804 21758
rect 49084 21812 49140 22094
rect 49532 22036 49588 23548
rect 49644 23380 49700 23390
rect 49644 23266 49700 23324
rect 49644 23214 49646 23266
rect 49698 23214 49700 23266
rect 49644 23202 49700 23214
rect 49756 23268 49812 26236
rect 49868 26226 49924 26236
rect 49980 26068 50036 26852
rect 49868 26012 50036 26068
rect 49868 24722 49924 26012
rect 50204 25060 50260 29820
rect 50428 29538 50484 30604
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50428 29486 50430 29538
rect 50482 29486 50484 29538
rect 50428 29474 50484 29486
rect 50876 29314 50932 29326
rect 50876 29262 50878 29314
rect 50930 29262 50932 29314
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50428 28084 50484 28094
rect 50652 28084 50708 28094
rect 50428 27858 50484 28028
rect 50428 27806 50430 27858
rect 50482 27806 50484 27858
rect 50428 27636 50484 27806
rect 50428 27570 50484 27580
rect 50540 28028 50652 28084
rect 50540 27188 50596 28028
rect 50652 28018 50708 28028
rect 50764 27746 50820 27758
rect 50764 27694 50766 27746
rect 50818 27694 50820 27746
rect 50764 27412 50820 27694
rect 50764 27346 50820 27356
rect 50316 27132 50596 27188
rect 50316 26404 50372 27132
rect 50540 27074 50596 27132
rect 50540 27022 50542 27074
rect 50594 27022 50596 27074
rect 50540 27010 50596 27022
rect 50316 26338 50372 26348
rect 50428 26962 50484 26974
rect 50428 26910 50430 26962
rect 50482 26910 50484 26962
rect 50428 25844 50484 26910
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50876 25844 50932 29262
rect 50988 27188 51044 30604
rect 51548 30324 51604 31614
rect 51324 30268 51604 30324
rect 51660 31892 51716 31902
rect 51212 28868 51268 28878
rect 51324 28868 51380 30268
rect 51548 30100 51604 30110
rect 51268 28812 51380 28868
rect 51436 29988 51492 29998
rect 51212 28802 51268 28812
rect 51436 28756 51492 29932
rect 51548 29986 51604 30044
rect 51548 29934 51550 29986
rect 51602 29934 51604 29986
rect 51548 29922 51604 29934
rect 51660 29652 51716 31836
rect 51996 31892 52164 31948
rect 52780 31892 52836 32622
rect 53116 31892 53172 31902
rect 51996 31890 52052 31892
rect 51996 31838 51998 31890
rect 52050 31838 52052 31890
rect 51996 31826 52052 31838
rect 52780 31890 53172 31892
rect 52780 31838 53118 31890
rect 53170 31838 53172 31890
rect 52780 31836 53172 31838
rect 52668 31780 52724 31790
rect 52668 31686 52724 31724
rect 51884 31668 51940 31678
rect 51940 31612 52164 31668
rect 51884 31574 51940 31612
rect 51884 31108 51940 31118
rect 51884 31014 51940 31052
rect 52108 31108 52164 31612
rect 52108 31014 52164 31052
rect 52556 31332 52612 31342
rect 52556 30994 52612 31276
rect 52780 31220 52836 31836
rect 53116 31826 53172 31836
rect 52780 31154 52836 31164
rect 53452 31780 53508 31790
rect 52556 30942 52558 30994
rect 52610 30942 52612 30994
rect 52556 30930 52612 30942
rect 52332 30882 52388 30894
rect 52332 30830 52334 30882
rect 52386 30830 52388 30882
rect 51884 30212 51940 30222
rect 51884 30118 51940 30156
rect 51324 28754 51492 28756
rect 51324 28702 51438 28754
rect 51490 28702 51492 28754
rect 51324 28700 51492 28702
rect 51324 27636 51380 28700
rect 51436 28690 51492 28700
rect 51548 29596 51716 29652
rect 52108 30100 52164 30110
rect 52332 30100 52388 30830
rect 52780 30884 52836 30894
rect 52780 30790 52836 30828
rect 53452 30322 53508 31724
rect 53788 31332 53844 34076
rect 53900 34130 53956 34142
rect 53900 34078 53902 34130
rect 53954 34078 53956 34130
rect 53900 33684 53956 34078
rect 54124 34132 54180 34974
rect 54124 34066 54180 34076
rect 54236 33796 54292 36204
rect 54460 35810 54516 36316
rect 54572 35922 54628 36428
rect 54684 36036 54740 36542
rect 54796 36482 54852 36988
rect 55020 36596 55076 37214
rect 56700 37156 56756 37166
rect 56588 37154 56756 37156
rect 56588 37102 56702 37154
rect 56754 37102 56756 37154
rect 56588 37100 56756 37102
rect 55468 37042 55524 37054
rect 55468 36990 55470 37042
rect 55522 36990 55524 37042
rect 55468 36820 55524 36990
rect 55468 36754 55524 36764
rect 56364 36820 56420 36830
rect 55020 36530 55076 36540
rect 55412 36596 55468 36606
rect 55468 36540 55524 36596
rect 55412 36530 55524 36540
rect 54796 36430 54798 36482
rect 54850 36430 54852 36482
rect 54796 36418 54852 36430
rect 55468 36482 55524 36530
rect 55468 36430 55470 36482
rect 55522 36430 55524 36482
rect 54684 35970 54740 35980
rect 54572 35870 54574 35922
rect 54626 35870 54628 35922
rect 54572 35858 54628 35870
rect 55132 35924 55188 35934
rect 54460 35758 54462 35810
rect 54514 35758 54516 35810
rect 54460 35746 54516 35758
rect 54796 35700 54852 35710
rect 54796 35606 54852 35644
rect 55132 35586 55188 35868
rect 55356 35700 55412 35710
rect 55356 35606 55412 35644
rect 55132 35534 55134 35586
rect 55186 35534 55188 35586
rect 55132 35364 55188 35534
rect 55468 35308 55524 36430
rect 55580 36594 55636 36606
rect 55580 36542 55582 36594
rect 55634 36542 55636 36594
rect 55580 36372 55636 36542
rect 55580 36306 55636 36316
rect 56028 36482 56084 36494
rect 56028 36430 56030 36482
rect 56082 36430 56084 36482
rect 56028 36372 56084 36430
rect 56364 36482 56420 36764
rect 56364 36430 56366 36482
rect 56418 36430 56420 36482
rect 56364 36418 56420 36430
rect 56028 36306 56084 36316
rect 56252 36258 56308 36270
rect 56252 36206 56254 36258
rect 56306 36206 56308 36258
rect 55132 35298 55188 35308
rect 55356 35252 55524 35308
rect 55580 36148 55636 36158
rect 56140 36148 56196 36158
rect 54460 34916 54516 34926
rect 54236 33730 54292 33740
rect 54348 34802 54404 34814
rect 54348 34750 54350 34802
rect 54402 34750 54404 34802
rect 53900 33618 53956 33628
rect 54012 33346 54068 33358
rect 54012 33294 54014 33346
rect 54066 33294 54068 33346
rect 54012 32564 54068 33294
rect 54236 33348 54292 33358
rect 54348 33348 54404 34750
rect 54292 33292 54404 33348
rect 54012 31778 54068 32508
rect 54012 31726 54014 31778
rect 54066 31726 54068 31778
rect 54012 31714 54068 31726
rect 54124 33122 54180 33134
rect 54124 33070 54126 33122
rect 54178 33070 54180 33122
rect 53788 31266 53844 31276
rect 53788 31108 53844 31118
rect 53788 30994 53844 31052
rect 53788 30942 53790 30994
rect 53842 30942 53844 30994
rect 53788 30930 53844 30942
rect 53900 30882 53956 30894
rect 53900 30830 53902 30882
rect 53954 30830 53956 30882
rect 53452 30270 53454 30322
rect 53506 30270 53508 30322
rect 53452 30258 53508 30270
rect 53676 30324 53732 30334
rect 53676 30230 53732 30268
rect 53116 30212 53172 30222
rect 52108 30098 52388 30100
rect 52108 30046 52110 30098
rect 52162 30046 52388 30098
rect 52108 30044 52388 30046
rect 53004 30100 53060 30110
rect 50988 26292 51044 27132
rect 51212 27580 51380 27636
rect 51436 27636 51492 27646
rect 51212 27076 51268 27580
rect 51212 26962 51268 27020
rect 51436 27074 51492 27580
rect 51436 27022 51438 27074
rect 51490 27022 51492 27074
rect 51436 27010 51492 27022
rect 51212 26910 51214 26962
rect 51266 26910 51268 26962
rect 51212 26898 51268 26910
rect 51548 26908 51604 29596
rect 51660 29426 51716 29438
rect 51660 29374 51662 29426
rect 51714 29374 51716 29426
rect 51660 28532 51716 29374
rect 52108 29316 52164 30044
rect 53004 30006 53060 30044
rect 52780 29988 52836 29998
rect 52780 29894 52836 29932
rect 52892 29986 52948 29998
rect 52892 29934 52894 29986
rect 52946 29934 52948 29986
rect 52892 29540 52948 29934
rect 52892 29474 52948 29484
rect 53116 29428 53172 30156
rect 53788 30100 53844 30110
rect 53564 29988 53620 29998
rect 52108 29260 53060 29316
rect 51772 28868 51828 28878
rect 51828 28812 51940 28868
rect 51772 28802 51828 28812
rect 51660 28466 51716 28476
rect 51772 28530 51828 28542
rect 51772 28478 51774 28530
rect 51826 28478 51828 28530
rect 51772 28196 51828 28478
rect 51660 28140 51828 28196
rect 51660 28084 51716 28140
rect 51660 28018 51716 28028
rect 51772 27972 51828 27982
rect 51772 27878 51828 27916
rect 51660 27858 51716 27870
rect 51660 27806 51662 27858
rect 51714 27806 51716 27858
rect 51660 27636 51716 27806
rect 51660 27570 51716 27580
rect 51660 27412 51716 27422
rect 51716 27356 51828 27412
rect 51660 27346 51716 27356
rect 51772 27074 51828 27356
rect 51772 27022 51774 27074
rect 51826 27022 51828 27074
rect 51772 27010 51828 27022
rect 50988 26198 51044 26236
rect 51100 26850 51156 26862
rect 51548 26852 51828 26908
rect 51100 26798 51102 26850
rect 51154 26798 51156 26850
rect 50428 25788 50596 25844
rect 50540 25284 50596 25788
rect 50876 25778 50932 25788
rect 50988 26066 51044 26078
rect 50988 26014 50990 26066
rect 51042 26014 51044 26066
rect 50876 25620 50932 25630
rect 50876 25526 50932 25564
rect 50652 25508 50708 25518
rect 50652 25414 50708 25452
rect 50204 24994 50260 25004
rect 50428 25228 50596 25284
rect 49868 24670 49870 24722
rect 49922 24670 49924 24722
rect 49868 24276 49924 24670
rect 49868 23716 49924 24220
rect 49868 23650 49924 23660
rect 49980 24836 50036 24846
rect 49980 23548 50036 24780
rect 50316 24724 50372 24734
rect 50428 24724 50484 25228
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50988 24948 51044 26014
rect 51100 25396 51156 26798
rect 51548 26516 51604 26526
rect 51324 26292 51380 26302
rect 51324 26198 51380 26236
rect 51548 26290 51604 26460
rect 51548 26238 51550 26290
rect 51602 26238 51604 26290
rect 51436 26178 51492 26190
rect 51436 26126 51438 26178
rect 51490 26126 51492 26178
rect 51324 25620 51380 25630
rect 51100 25340 51268 25396
rect 50988 24882 51044 24892
rect 51100 24836 51156 24846
rect 51100 24742 51156 24780
rect 50372 24668 50484 24724
rect 50988 24724 51044 24734
rect 50316 24658 50372 24668
rect 50092 24612 50148 24622
rect 50092 23604 50148 24556
rect 50204 24610 50260 24622
rect 50204 24558 50206 24610
rect 50258 24558 50260 24610
rect 50204 24388 50260 24558
rect 50988 24612 51044 24668
rect 50988 24556 51156 24612
rect 50428 24500 50484 24510
rect 50428 24406 50484 24444
rect 50764 24498 50820 24510
rect 50764 24446 50766 24498
rect 50818 24446 50820 24498
rect 50204 24322 50260 24332
rect 50764 24052 50820 24446
rect 50764 23986 50820 23996
rect 50428 23938 50484 23950
rect 50428 23886 50430 23938
rect 50482 23886 50484 23938
rect 50428 23604 50484 23886
rect 50876 23940 50932 23950
rect 50876 23846 50932 23884
rect 50092 23548 50260 23604
rect 49980 23482 50036 23492
rect 49756 23212 50148 23268
rect 50092 23154 50148 23212
rect 50092 23102 50094 23154
rect 50146 23102 50148 23154
rect 50092 23090 50148 23102
rect 49756 23042 49812 23054
rect 49756 22990 49758 23042
rect 49810 22990 49812 23042
rect 49756 22820 49812 22990
rect 49756 22754 49812 22764
rect 49868 23044 49924 23054
rect 49868 22482 49924 22988
rect 49980 23042 50036 23054
rect 49980 22990 49982 23042
rect 50034 22990 50036 23042
rect 49980 22932 50036 22990
rect 50092 22932 50148 22942
rect 49980 22876 50092 22932
rect 50092 22866 50148 22876
rect 49868 22430 49870 22482
rect 49922 22430 49924 22482
rect 49868 22418 49924 22430
rect 49756 22258 49812 22270
rect 49756 22206 49758 22258
rect 49810 22206 49812 22258
rect 49756 22036 49812 22206
rect 49980 22260 50036 22270
rect 49980 22166 50036 22204
rect 49532 21980 49700 22036
rect 49532 21812 49588 21822
rect 49084 21810 49588 21812
rect 49084 21758 49534 21810
rect 49586 21758 49588 21810
rect 49084 21756 49588 21758
rect 48972 21588 49028 21598
rect 48972 21494 49028 21532
rect 48300 21474 48356 21486
rect 48300 21422 48302 21474
rect 48354 21422 48356 21474
rect 48300 21252 48356 21422
rect 49084 21476 49140 21756
rect 49532 21746 49588 21756
rect 49644 21812 49700 21980
rect 49756 21970 49812 21980
rect 49644 21746 49700 21756
rect 49644 21588 49700 21598
rect 50204 21588 50260 23548
rect 50316 23548 50484 23604
rect 50988 23826 51044 23838
rect 50988 23774 50990 23826
rect 51042 23774 51044 23826
rect 50556 23548 50820 23558
rect 50316 23380 50372 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50316 23314 50372 23324
rect 50764 23380 50820 23390
rect 50764 23266 50820 23324
rect 50764 23214 50766 23266
rect 50818 23214 50820 23266
rect 50764 23202 50820 23214
rect 50876 23378 50932 23390
rect 50876 23326 50878 23378
rect 50930 23326 50932 23378
rect 50540 23156 50596 23166
rect 50540 23062 50596 23100
rect 50764 23044 50820 23054
rect 50764 22596 50820 22988
rect 50428 22372 50484 22382
rect 50428 22258 50484 22316
rect 50764 22370 50820 22540
rect 50764 22318 50766 22370
rect 50818 22318 50820 22370
rect 50764 22306 50820 22318
rect 50428 22206 50430 22258
rect 50482 22206 50484 22258
rect 50428 22194 50484 22206
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50876 21700 50932 23326
rect 50988 22594 51044 23774
rect 51100 23156 51156 24556
rect 51212 23938 51268 25340
rect 51324 24722 51380 25564
rect 51436 25284 51492 26126
rect 51548 25732 51604 26238
rect 51548 25676 51716 25732
rect 51436 25218 51492 25228
rect 51548 25508 51604 25518
rect 51324 24670 51326 24722
rect 51378 24670 51380 24722
rect 51324 24658 51380 24670
rect 51212 23886 51214 23938
rect 51266 23886 51268 23938
rect 51212 23874 51268 23886
rect 51436 23940 51492 23950
rect 51436 23846 51492 23884
rect 51436 23268 51492 23278
rect 51548 23268 51604 25452
rect 51660 25396 51716 25676
rect 51660 25330 51716 25340
rect 51660 23826 51716 23838
rect 51660 23774 51662 23826
rect 51714 23774 51716 23826
rect 51660 23380 51716 23774
rect 51772 23380 51828 26852
rect 51884 26516 51940 28812
rect 52108 28756 52164 28766
rect 52108 28754 52948 28756
rect 52108 28702 52110 28754
rect 52162 28702 52948 28754
rect 52108 28700 52948 28702
rect 52108 28690 52164 28700
rect 52780 28532 52836 28542
rect 51996 28420 52052 28430
rect 51996 28418 52164 28420
rect 51996 28366 51998 28418
rect 52050 28366 52164 28418
rect 51996 28364 52164 28366
rect 51996 28354 52052 28364
rect 52108 28084 52164 28364
rect 52108 28028 52612 28084
rect 52332 27860 52388 27870
rect 52332 27766 52388 27804
rect 52220 27634 52276 27646
rect 52220 27582 52222 27634
rect 52274 27582 52276 27634
rect 52108 26962 52164 26974
rect 52108 26910 52110 26962
rect 52162 26910 52164 26962
rect 51996 26852 52052 26862
rect 51996 26758 52052 26796
rect 51884 26450 51940 26460
rect 52108 25956 52164 26910
rect 52220 26178 52276 27582
rect 52332 27076 52388 27086
rect 52332 26290 52388 27020
rect 52332 26238 52334 26290
rect 52386 26238 52388 26290
rect 52332 26226 52388 26238
rect 52556 26292 52612 28028
rect 52780 27858 52836 28476
rect 52892 28084 52948 28700
rect 53004 28642 53060 29260
rect 53116 28754 53172 29372
rect 53228 29426 53284 29438
rect 53228 29374 53230 29426
rect 53282 29374 53284 29426
rect 53228 28866 53284 29374
rect 53228 28814 53230 28866
rect 53282 28814 53284 28866
rect 53228 28802 53284 28814
rect 53564 28980 53620 29932
rect 53116 28702 53118 28754
rect 53170 28702 53172 28754
rect 53116 28690 53172 28702
rect 53004 28590 53006 28642
rect 53058 28590 53060 28642
rect 53004 28578 53060 28590
rect 52892 28028 53508 28084
rect 52780 27806 52782 27858
rect 52834 27806 52836 27858
rect 52780 27794 52836 27806
rect 53452 27858 53508 28028
rect 53452 27806 53454 27858
rect 53506 27806 53508 27858
rect 53452 27794 53508 27806
rect 53228 27636 53284 27646
rect 53116 27634 53284 27636
rect 53116 27582 53230 27634
rect 53282 27582 53284 27634
rect 53116 27580 53284 27582
rect 52780 27188 52836 27198
rect 52780 27094 52836 27132
rect 53116 26908 53172 27580
rect 53228 27570 53284 27580
rect 53228 27412 53284 27422
rect 53564 27412 53620 28924
rect 53284 27356 53620 27412
rect 53676 28868 53732 28878
rect 53228 27298 53284 27356
rect 53228 27246 53230 27298
rect 53282 27246 53284 27298
rect 53228 27234 53284 27246
rect 53340 27076 53396 27086
rect 53116 26852 53284 26908
rect 52220 26126 52222 26178
rect 52274 26126 52276 26178
rect 52220 26114 52276 26126
rect 52444 26066 52500 26078
rect 52444 26014 52446 26066
rect 52498 26014 52500 26066
rect 52444 25956 52500 26014
rect 52108 25900 52500 25956
rect 52444 25508 52500 25900
rect 52556 25732 52612 26236
rect 52556 25666 52612 25676
rect 52892 25620 52948 25630
rect 52892 25526 52948 25564
rect 52780 25508 52836 25518
rect 52444 25506 52836 25508
rect 52444 25454 52782 25506
rect 52834 25454 52836 25506
rect 52444 25452 52836 25454
rect 52780 25442 52836 25452
rect 51996 25396 52052 25406
rect 51884 25340 51996 25396
rect 51884 24052 51940 25340
rect 51996 25330 52052 25340
rect 52668 25284 52724 25294
rect 52556 24836 52612 24846
rect 52444 24780 52556 24836
rect 51996 24724 52052 24734
rect 51996 24630 52052 24668
rect 51884 23996 52052 24052
rect 51996 23940 52052 23996
rect 51996 23884 52164 23940
rect 51884 23828 51940 23838
rect 51884 23826 52052 23828
rect 51884 23774 51886 23826
rect 51938 23774 52052 23826
rect 51884 23772 52052 23774
rect 51884 23762 51940 23772
rect 51884 23380 51940 23390
rect 51772 23378 51940 23380
rect 51772 23326 51886 23378
rect 51938 23326 51940 23378
rect 51772 23324 51940 23326
rect 51660 23314 51716 23324
rect 51492 23212 51604 23268
rect 51884 23268 51940 23324
rect 51436 23202 51492 23212
rect 51884 23202 51940 23212
rect 51324 23156 51380 23166
rect 51100 23154 51380 23156
rect 51100 23102 51326 23154
rect 51378 23102 51380 23154
rect 51100 23100 51380 23102
rect 51324 23044 51380 23100
rect 51324 22988 51492 23044
rect 51100 22932 51156 22942
rect 51100 22838 51156 22876
rect 50988 22542 50990 22594
rect 51042 22542 51044 22594
rect 50988 22530 51044 22542
rect 51212 22484 51268 22494
rect 51212 22390 51268 22428
rect 51436 22372 51492 22988
rect 51772 23042 51828 23054
rect 51772 22990 51774 23042
rect 51826 22990 51828 23042
rect 51660 22930 51716 22942
rect 51660 22878 51662 22930
rect 51714 22878 51716 22930
rect 51660 22594 51716 22878
rect 51772 22932 51828 22990
rect 51772 22866 51828 22876
rect 51660 22542 51662 22594
rect 51714 22542 51716 22594
rect 51660 22530 51716 22542
rect 51660 22372 51716 22382
rect 51436 22370 51716 22372
rect 51436 22318 51662 22370
rect 51714 22318 51716 22370
rect 51436 22316 51716 22318
rect 51660 22306 51716 22316
rect 51996 22372 52052 23772
rect 52108 23156 52164 23884
rect 52332 23380 52388 23390
rect 52332 23286 52388 23324
rect 52444 23268 52500 24780
rect 52556 24770 52612 24780
rect 52668 24834 52724 25228
rect 52668 24782 52670 24834
rect 52722 24782 52724 24834
rect 52668 24770 52724 24782
rect 53228 24500 53284 26852
rect 53340 26290 53396 27020
rect 53676 27074 53732 28812
rect 53788 28756 53844 30044
rect 53900 29426 53956 30830
rect 53900 29374 53902 29426
rect 53954 29374 53956 29426
rect 53900 29316 53956 29374
rect 53900 29250 53956 29260
rect 54012 29986 54068 29998
rect 54012 29934 54014 29986
rect 54066 29934 54068 29986
rect 53788 28642 53844 28700
rect 53788 28590 53790 28642
rect 53842 28590 53844 28642
rect 53788 28578 53844 28590
rect 54012 28644 54068 29934
rect 53676 27022 53678 27074
rect 53730 27022 53732 27074
rect 53676 27010 53732 27022
rect 53788 27972 53844 27982
rect 53788 27074 53844 27916
rect 53900 27972 53956 27982
rect 54012 27972 54068 28588
rect 53900 27970 54068 27972
rect 53900 27918 53902 27970
rect 53954 27918 54068 27970
rect 53900 27916 54068 27918
rect 54124 28084 54180 33070
rect 54236 32562 54292 33292
rect 54236 32510 54238 32562
rect 54290 32510 54292 32562
rect 54236 32498 54292 32510
rect 54460 31948 54516 34860
rect 55356 34916 55412 35252
rect 55580 35140 55636 36092
rect 56028 36092 56140 36148
rect 56028 35810 56084 36092
rect 56140 36082 56196 36092
rect 56028 35758 56030 35810
rect 56082 35758 56084 35810
rect 56028 35746 56084 35758
rect 55580 35074 55636 35084
rect 55804 35588 55860 35598
rect 55356 34850 55412 34860
rect 54684 34692 54740 34702
rect 54684 33234 54740 34636
rect 55580 34020 55636 34030
rect 55020 34018 55636 34020
rect 55020 33966 55582 34018
rect 55634 33966 55636 34018
rect 55020 33964 55636 33966
rect 55020 33348 55076 33964
rect 55580 33954 55636 33964
rect 55804 33458 55860 35532
rect 55916 35476 55972 35486
rect 55916 34690 55972 35420
rect 56028 34804 56084 34814
rect 56252 34804 56308 36206
rect 56028 34802 56308 34804
rect 56028 34750 56030 34802
rect 56082 34750 56308 34802
rect 56028 34748 56308 34750
rect 56588 35698 56644 37100
rect 56700 37090 56756 37100
rect 56700 36370 56756 36382
rect 56700 36318 56702 36370
rect 56754 36318 56756 36370
rect 56700 35924 56756 36318
rect 56812 35924 56868 37324
rect 57260 37154 57316 37166
rect 57260 37102 57262 37154
rect 57314 37102 57316 37154
rect 57036 36370 57092 36382
rect 57036 36318 57038 36370
rect 57090 36318 57092 36370
rect 57036 36148 57092 36318
rect 57036 36082 57092 36092
rect 57148 36258 57204 36270
rect 57148 36206 57150 36258
rect 57202 36206 57204 36258
rect 57148 35924 57204 36206
rect 57260 36260 57316 37102
rect 57260 36166 57316 36204
rect 57820 36260 57876 36270
rect 57372 36036 57428 36046
rect 56812 35868 57092 35924
rect 57148 35868 57316 35924
rect 56700 35858 56756 35868
rect 56588 35646 56590 35698
rect 56642 35646 56644 35698
rect 56588 34804 56644 35646
rect 56924 35698 56980 35710
rect 56924 35646 56926 35698
rect 56978 35646 56980 35698
rect 56700 35588 56756 35598
rect 56700 35494 56756 35532
rect 56812 34916 56868 34926
rect 56812 34822 56868 34860
rect 56028 34738 56084 34748
rect 55916 34638 55918 34690
rect 55970 34638 55972 34690
rect 55916 34626 55972 34638
rect 56588 34356 56644 34748
rect 56812 34692 56868 34702
rect 56924 34692 56980 35646
rect 57036 35700 57092 35868
rect 57148 35700 57204 35710
rect 57036 35698 57204 35700
rect 57036 35646 57150 35698
rect 57202 35646 57204 35698
rect 57036 35644 57204 35646
rect 57036 35140 57092 35644
rect 57148 35634 57204 35644
rect 57148 35474 57204 35486
rect 57148 35422 57150 35474
rect 57202 35422 57204 35474
rect 57148 35364 57204 35422
rect 57148 35298 57204 35308
rect 57036 34916 57092 35084
rect 57148 35140 57204 35150
rect 57260 35140 57316 35868
rect 57148 35138 57316 35140
rect 57148 35086 57150 35138
rect 57202 35086 57316 35138
rect 57148 35084 57316 35086
rect 57148 35074 57204 35084
rect 57148 34916 57204 34926
rect 57036 34914 57204 34916
rect 57036 34862 57150 34914
rect 57202 34862 57204 34914
rect 57036 34860 57204 34862
rect 56868 34636 56980 34692
rect 57036 34690 57092 34702
rect 57036 34638 57038 34690
rect 57090 34638 57092 34690
rect 56812 34626 56868 34636
rect 56588 34300 56756 34356
rect 56028 34244 56084 34254
rect 56028 34150 56084 34188
rect 56476 34130 56532 34142
rect 56476 34078 56478 34130
rect 56530 34078 56532 34130
rect 56476 34020 56532 34078
rect 56476 33954 56532 33964
rect 55804 33406 55806 33458
rect 55858 33406 55860 33458
rect 55804 33394 55860 33406
rect 54684 33182 54686 33234
rect 54738 33182 54740 33234
rect 54684 33170 54740 33182
rect 54908 33346 55076 33348
rect 54908 33294 55022 33346
rect 55074 33294 55076 33346
rect 54908 33292 55076 33294
rect 54796 32676 54852 32686
rect 54796 32582 54852 32620
rect 54348 31892 54516 31948
rect 54236 31668 54292 31678
rect 54348 31668 54404 31892
rect 54796 31780 54852 31790
rect 54236 31666 54404 31668
rect 54236 31614 54238 31666
rect 54290 31614 54404 31666
rect 54236 31612 54404 31614
rect 54684 31778 54852 31780
rect 54684 31726 54798 31778
rect 54850 31726 54852 31778
rect 54684 31724 54852 31726
rect 54236 31602 54292 31612
rect 54572 31554 54628 31566
rect 54572 31502 54574 31554
rect 54626 31502 54628 31554
rect 54348 31332 54404 31342
rect 54348 29652 54404 31276
rect 54572 31108 54628 31502
rect 54572 31042 54628 31052
rect 54572 30324 54628 30334
rect 54684 30324 54740 31724
rect 54796 31714 54852 31724
rect 54908 30996 54964 33292
rect 55020 33282 55076 33292
rect 56700 32786 56756 34300
rect 56812 34132 56868 34142
rect 56812 34038 56868 34076
rect 56700 32734 56702 32786
rect 56754 32734 56756 32786
rect 56700 32722 56756 32734
rect 55244 32676 55300 32686
rect 55244 31890 55300 32620
rect 57036 31948 57092 34638
rect 57148 34244 57204 34860
rect 57148 34178 57204 34188
rect 57260 34916 57316 34926
rect 57260 34130 57316 34860
rect 57260 34078 57262 34130
rect 57314 34078 57316 34130
rect 57260 34066 57316 34078
rect 57372 34018 57428 35980
rect 57820 35924 57876 36204
rect 57932 35924 57988 35934
rect 57820 35922 57988 35924
rect 57820 35870 57934 35922
rect 57986 35870 57988 35922
rect 57820 35868 57988 35870
rect 57932 35858 57988 35868
rect 57820 35586 57876 35598
rect 57820 35534 57822 35586
rect 57874 35534 57876 35586
rect 57708 35476 57764 35486
rect 57708 35382 57764 35420
rect 57820 35364 57876 35534
rect 57820 35298 57876 35308
rect 57820 34804 57876 34814
rect 57820 34802 57988 34804
rect 57820 34750 57822 34802
rect 57874 34750 57988 34802
rect 57820 34748 57988 34750
rect 57820 34738 57876 34748
rect 57708 34692 57764 34702
rect 57708 34598 57764 34636
rect 57372 33966 57374 34018
rect 57426 33966 57428 34018
rect 57372 33954 57428 33966
rect 57932 33458 57988 34748
rect 57932 33406 57934 33458
rect 57986 33406 57988 33458
rect 57932 33348 57988 33406
rect 57932 33282 57988 33292
rect 57036 31892 57428 31948
rect 55244 31838 55246 31890
rect 55298 31838 55300 31890
rect 55244 31826 55300 31838
rect 57372 31890 57428 31892
rect 57372 31838 57374 31890
rect 57426 31838 57428 31890
rect 57372 31826 57428 31838
rect 58044 31778 58100 31790
rect 58044 31726 58046 31778
rect 58098 31726 58100 31778
rect 56700 31556 56756 31566
rect 54908 30902 54964 30940
rect 55356 30996 55412 31006
rect 55356 30902 55412 30940
rect 54628 30268 54740 30324
rect 54572 30230 54628 30268
rect 56700 30210 56756 31500
rect 56700 30158 56702 30210
rect 56754 30158 56756 30210
rect 56700 30146 56756 30158
rect 57372 30996 57428 31006
rect 57372 30210 57428 30940
rect 58044 30996 58100 31726
rect 58044 30930 58100 30940
rect 57372 30158 57374 30210
rect 57426 30158 57428 30210
rect 57372 30146 57428 30158
rect 54348 29596 55412 29652
rect 54348 29314 54404 29596
rect 54796 29428 54852 29438
rect 54796 29334 54852 29372
rect 54348 29262 54350 29314
rect 54402 29262 54404 29314
rect 54348 29250 54404 29262
rect 54460 29316 54516 29326
rect 54236 28980 54292 28990
rect 54236 28642 54292 28924
rect 54236 28590 54238 28642
rect 54290 28590 54292 28642
rect 54236 28578 54292 28590
rect 54124 27970 54180 28028
rect 54124 27918 54126 27970
rect 54178 27918 54180 27970
rect 53900 27906 53956 27916
rect 54124 27906 54180 27918
rect 54460 27972 54516 29260
rect 54908 28756 54964 28766
rect 54908 28662 54964 28700
rect 55020 28530 55076 29596
rect 55356 29426 55412 29596
rect 55356 29374 55358 29426
rect 55410 29374 55412 29426
rect 55356 29362 55412 29374
rect 55132 29202 55188 29214
rect 55132 29150 55134 29202
rect 55186 29150 55188 29202
rect 55132 28868 55188 29150
rect 55356 28868 55412 28878
rect 55132 28812 55356 28868
rect 55356 28642 55412 28812
rect 56252 28868 56308 28878
rect 55356 28590 55358 28642
rect 55410 28590 55412 28642
rect 55356 28578 55412 28590
rect 55692 28642 55748 28654
rect 55692 28590 55694 28642
rect 55746 28590 55748 28642
rect 55020 28478 55022 28530
rect 55074 28478 55076 28530
rect 55020 28466 55076 28478
rect 55468 28420 55524 28430
rect 54460 27906 54516 27916
rect 55020 28196 55076 28206
rect 55020 27860 55076 28140
rect 55020 27766 55076 27804
rect 54236 27748 54292 27758
rect 54124 27692 54236 27748
rect 53788 27022 53790 27074
rect 53842 27022 53844 27074
rect 53788 27010 53844 27022
rect 54012 27076 54068 27086
rect 54124 27076 54180 27692
rect 54236 27654 54292 27692
rect 54012 27074 54180 27076
rect 54012 27022 54014 27074
rect 54066 27022 54180 27074
rect 54012 27020 54180 27022
rect 54348 27636 54404 27646
rect 54012 27010 54068 27020
rect 53676 26852 53732 26862
rect 53340 26238 53342 26290
rect 53394 26238 53396 26290
rect 53340 26226 53396 26238
rect 53452 26402 53508 26414
rect 53452 26350 53454 26402
rect 53506 26350 53508 26402
rect 53452 25508 53508 26350
rect 53340 25452 53508 25508
rect 53340 25394 53396 25452
rect 53340 25342 53342 25394
rect 53394 25342 53396 25394
rect 53340 24836 53396 25342
rect 53340 24770 53396 24780
rect 53676 24724 53732 26796
rect 53900 26404 53956 26414
rect 53900 26310 53956 26348
rect 54348 26290 54404 27580
rect 55468 27188 55524 28364
rect 55692 28196 55748 28590
rect 56252 28530 56308 28812
rect 56476 28644 56532 28654
rect 56476 28550 56532 28588
rect 56252 28478 56254 28530
rect 56306 28478 56308 28530
rect 56252 28466 56308 28478
rect 55692 28130 55748 28140
rect 56812 28084 56868 28094
rect 56588 27972 56644 27982
rect 56588 27878 56644 27916
rect 55580 27858 55636 27870
rect 55580 27806 55582 27858
rect 55634 27806 55636 27858
rect 55580 27748 55636 27806
rect 56812 27858 56868 28028
rect 56812 27806 56814 27858
rect 56866 27806 56868 27858
rect 56812 27794 56868 27806
rect 55580 27682 55636 27692
rect 57708 27748 57764 27758
rect 55580 27188 55636 27198
rect 55468 27186 55636 27188
rect 55468 27134 55582 27186
rect 55634 27134 55636 27186
rect 55468 27132 55636 27134
rect 55580 27122 55636 27132
rect 57708 27186 57764 27692
rect 57708 27134 57710 27186
rect 57762 27134 57764 27186
rect 57708 27122 57764 27134
rect 54908 27074 54964 27086
rect 54908 27022 54910 27074
rect 54962 27022 54964 27074
rect 54460 26964 54516 26974
rect 54460 26870 54516 26908
rect 54908 26964 54964 27022
rect 54908 26898 54964 26908
rect 54796 26292 54852 26302
rect 54348 26238 54350 26290
rect 54402 26238 54404 26290
rect 54348 26226 54404 26238
rect 54460 26290 54852 26292
rect 54460 26238 54798 26290
rect 54850 26238 54852 26290
rect 54460 26236 54852 26238
rect 53900 25732 53956 25742
rect 54460 25732 54516 26236
rect 53900 25638 53956 25676
rect 54012 25676 54516 25732
rect 54012 25618 54068 25676
rect 54012 25566 54014 25618
rect 54066 25566 54068 25618
rect 54012 25554 54068 25566
rect 54460 25396 54516 25406
rect 54460 25302 54516 25340
rect 53228 24444 53396 24500
rect 53228 24276 53284 24286
rect 53228 24050 53284 24220
rect 53228 23998 53230 24050
rect 53282 23998 53284 24050
rect 53228 23986 53284 23998
rect 52780 23828 52836 23838
rect 52780 23734 52836 23772
rect 53004 23268 53060 23278
rect 52444 23266 52948 23268
rect 52444 23214 52446 23266
rect 52498 23214 52948 23266
rect 52444 23212 52948 23214
rect 52444 23202 52500 23212
rect 52108 22482 52164 23100
rect 52892 23044 52948 23212
rect 53004 23174 53060 23212
rect 53340 23044 53396 24444
rect 53676 24050 53732 24668
rect 54796 24610 54852 26236
rect 54796 24558 54798 24610
rect 54850 24558 54852 24610
rect 54796 24546 54852 24558
rect 53676 23998 53678 24050
rect 53730 23998 53732 24050
rect 53676 23986 53732 23998
rect 52892 22988 53172 23044
rect 52108 22430 52110 22482
rect 52162 22430 52164 22482
rect 52108 22418 52164 22430
rect 51996 22306 52052 22316
rect 50988 21700 51044 21710
rect 50876 21698 51044 21700
rect 50876 21646 50990 21698
rect 51042 21646 51044 21698
rect 50876 21644 51044 21646
rect 50988 21634 51044 21644
rect 49644 21494 49700 21532
rect 49868 21586 50260 21588
rect 49868 21534 50206 21586
rect 50258 21534 50260 21586
rect 49868 21532 50260 21534
rect 49084 21410 49140 21420
rect 49532 21364 49588 21374
rect 49532 21270 49588 21308
rect 48300 21186 48356 21196
rect 48300 20916 48356 20926
rect 48188 20914 48356 20916
rect 48188 20862 48302 20914
rect 48354 20862 48356 20914
rect 48188 20860 48356 20862
rect 48300 20850 48356 20860
rect 48636 20916 48692 20926
rect 48636 20822 48692 20860
rect 49868 20916 49924 21532
rect 50204 21522 50260 21532
rect 53116 21474 53172 22988
rect 53340 22978 53396 22988
rect 53116 21422 53118 21474
rect 53170 21422 53172 21474
rect 53116 21410 53172 21422
rect 49868 20822 49924 20860
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 47180 20190 47182 20242
rect 47234 20190 47236 20242
rect 45836 20178 45892 20188
rect 47180 20178 47236 20190
rect 41692 20078 41694 20130
rect 41746 20078 41748 20130
rect 41692 20066 41748 20078
rect 38556 19908 38612 19918
rect 39788 19908 39844 19918
rect 38444 19852 38556 19908
rect 38612 19852 38724 19908
rect 37100 19814 37156 19852
rect 38556 19814 38612 19852
rect 37100 19348 37156 19358
rect 36988 19346 37156 19348
rect 36988 19294 37102 19346
rect 37154 19294 37156 19346
rect 36988 19292 37156 19294
rect 37100 19282 37156 19292
rect 35980 19236 36036 19246
rect 35420 19122 35588 19124
rect 35420 19070 35422 19122
rect 35474 19070 35588 19122
rect 35420 19068 35588 19070
rect 35756 19234 36036 19236
rect 35756 19182 35982 19234
rect 36034 19182 36036 19234
rect 35756 19180 36036 19182
rect 35420 19058 35476 19068
rect 35308 18946 35364 18956
rect 35308 18338 35364 18350
rect 35308 18286 35310 18338
rect 35362 18286 35364 18338
rect 35308 18228 35364 18286
rect 35756 18228 35812 19180
rect 35980 19170 36036 19180
rect 36316 19012 36372 19022
rect 35308 18172 35812 18228
rect 35868 19010 36372 19012
rect 35868 18958 36318 19010
rect 36370 18958 36372 19010
rect 35868 18956 36372 18958
rect 34860 18060 35140 18116
rect 35196 18060 35460 18070
rect 33852 17668 33908 17678
rect 33852 17666 34020 17668
rect 33852 17614 33854 17666
rect 33906 17614 34020 17666
rect 33852 17612 34020 17614
rect 33852 17602 33908 17612
rect 33628 16830 33630 16882
rect 33682 16830 33684 16882
rect 33628 16098 33684 16830
rect 33964 16324 34020 17612
rect 34076 17444 34132 17454
rect 34076 17442 34356 17444
rect 34076 17390 34078 17442
rect 34130 17390 34356 17442
rect 34076 17388 34356 17390
rect 34076 17378 34132 17388
rect 34300 16994 34356 17388
rect 34300 16942 34302 16994
rect 34354 16942 34356 16994
rect 34300 16930 34356 16942
rect 34188 16324 34244 16334
rect 33964 16322 34244 16324
rect 33964 16270 34190 16322
rect 34242 16270 34244 16322
rect 33964 16268 34244 16270
rect 34188 16258 34244 16268
rect 33628 16046 33630 16098
rect 33682 16046 33684 16098
rect 33628 15540 33684 16046
rect 34524 16098 34580 16110
rect 34524 16046 34526 16098
rect 34578 16046 34580 16098
rect 33628 15474 33684 15484
rect 33852 15652 33908 15662
rect 33852 15538 33908 15596
rect 33852 15486 33854 15538
rect 33906 15486 33908 15538
rect 33852 15474 33908 15486
rect 34524 15316 34580 16046
rect 34748 16100 34804 16110
rect 34748 15986 34804 16044
rect 34748 15934 34750 15986
rect 34802 15934 34804 15986
rect 34748 15922 34804 15934
rect 34860 15426 34916 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35084 16660 35140 16670
rect 35084 15986 35140 16604
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35084 15934 35086 15986
rect 35138 15934 35140 15986
rect 35084 15922 35140 15934
rect 35532 16100 35588 16110
rect 34860 15374 34862 15426
rect 34914 15374 34916 15426
rect 34860 15362 34916 15374
rect 34188 15204 34244 15242
rect 34188 15138 34244 15148
rect 34300 13858 34356 13870
rect 34300 13806 34302 13858
rect 34354 13806 34356 13858
rect 33516 13694 33518 13746
rect 33570 13694 33572 13746
rect 33516 13682 33572 13694
rect 33964 13746 34020 13758
rect 33964 13694 33966 13746
rect 34018 13694 34020 13746
rect 32732 13074 33012 13076
rect 32732 13022 32734 13074
rect 32786 13022 33012 13074
rect 32732 13020 33012 13022
rect 32732 13010 32788 13020
rect 31500 12910 31502 12962
rect 31554 12910 31556 12962
rect 31500 12898 31556 12910
rect 31276 12798 31278 12850
rect 31330 12798 31332 12850
rect 31276 12786 31332 12798
rect 30380 11620 30436 11630
rect 30380 11526 30436 11564
rect 30716 11620 30772 12348
rect 32956 12180 33012 13020
rect 33180 12964 33236 12974
rect 33180 12962 33348 12964
rect 33180 12910 33182 12962
rect 33234 12910 33348 12962
rect 33180 12908 33348 12910
rect 33180 12898 33236 12908
rect 33068 12180 33124 12190
rect 32956 12178 33236 12180
rect 32956 12126 33070 12178
rect 33122 12126 33236 12178
rect 32956 12124 33236 12126
rect 33068 12114 33124 12124
rect 30716 11554 30772 11564
rect 31500 11732 31556 11742
rect 30604 11508 30660 11518
rect 30604 11282 30660 11452
rect 30604 11230 30606 11282
rect 30658 11230 30660 11282
rect 30044 11170 30100 11182
rect 30044 11118 30046 11170
rect 30098 11118 30100 11170
rect 29932 10836 29988 10846
rect 29652 10834 29988 10836
rect 29652 10782 29934 10834
rect 29986 10782 29988 10834
rect 29652 10780 29988 10782
rect 29596 10742 29652 10780
rect 29932 10770 29988 10780
rect 29932 9828 29988 9838
rect 30044 9828 30100 11118
rect 30268 10836 30324 10846
rect 30268 10742 30324 10780
rect 30604 10612 30660 11230
rect 30940 11284 30996 11294
rect 30940 11190 30996 11228
rect 31500 10836 31556 11676
rect 30828 10724 30884 10734
rect 30716 10612 30772 10622
rect 30604 10610 30772 10612
rect 30604 10558 30718 10610
rect 30770 10558 30772 10610
rect 30604 10556 30772 10558
rect 30716 10546 30772 10556
rect 29932 9826 30100 9828
rect 29932 9774 29934 9826
rect 29986 9774 30100 9826
rect 29932 9772 30100 9774
rect 29932 9762 29988 9772
rect 30156 9604 30212 9614
rect 30156 9510 30212 9548
rect 29260 8878 29262 8930
rect 29314 8878 29316 8930
rect 29260 8866 29316 8878
rect 30716 8372 30772 8382
rect 30828 8372 30884 10668
rect 31500 10610 31556 10780
rect 31500 10558 31502 10610
rect 31554 10558 31556 10610
rect 31500 10546 31556 10558
rect 31836 10388 31892 10398
rect 31612 10386 31892 10388
rect 31612 10334 31838 10386
rect 31890 10334 31892 10386
rect 31612 10332 31892 10334
rect 31612 9940 31668 10332
rect 31836 10322 31892 10332
rect 31052 9884 31668 9940
rect 31052 9826 31108 9884
rect 31052 9774 31054 9826
rect 31106 9774 31108 9826
rect 31052 9762 31108 9774
rect 30716 8370 30884 8372
rect 30716 8318 30718 8370
rect 30770 8318 30884 8370
rect 30716 8316 30884 8318
rect 31276 9602 31332 9614
rect 31276 9550 31278 9602
rect 31330 9550 31332 9602
rect 31276 8372 31332 9550
rect 31388 9604 31444 9614
rect 31388 9154 31444 9548
rect 33180 9268 33236 12124
rect 33292 11618 33348 12908
rect 33404 12740 33460 12750
rect 33404 12738 33908 12740
rect 33404 12686 33406 12738
rect 33458 12686 33908 12738
rect 33404 12684 33908 12686
rect 33404 12674 33460 12684
rect 33852 12290 33908 12684
rect 33852 12238 33854 12290
rect 33906 12238 33908 12290
rect 33852 12226 33908 12238
rect 33964 11956 34020 13694
rect 33964 11890 34020 11900
rect 34300 12068 34356 13806
rect 33292 11566 33294 11618
rect 33346 11566 33348 11618
rect 33292 11554 33348 11566
rect 33628 11732 33684 11742
rect 33628 11618 33684 11676
rect 33628 11566 33630 11618
rect 33682 11566 33684 11618
rect 33628 11554 33684 11566
rect 33852 11396 33908 11406
rect 33852 11282 33908 11340
rect 33852 11230 33854 11282
rect 33906 11230 33908 11282
rect 33852 11218 33908 11230
rect 34300 11282 34356 12012
rect 34524 11732 34580 15260
rect 34972 15314 35028 15326
rect 34972 15262 34974 15314
rect 35026 15262 35028 15314
rect 34972 14084 35028 15262
rect 35084 15204 35140 15214
rect 35084 14418 35140 15148
rect 35420 15204 35476 15242
rect 35420 15138 35476 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35084 14366 35086 14418
rect 35138 14366 35140 14418
rect 35084 14354 35140 14366
rect 35532 14418 35588 16044
rect 35532 14366 35534 14418
rect 35586 14366 35588 14418
rect 35532 14354 35588 14366
rect 34972 14018 35028 14028
rect 35084 13636 35140 13646
rect 35084 13188 35140 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 13188 35252 13198
rect 35084 13186 35252 13188
rect 35084 13134 35198 13186
rect 35250 13134 35252 13186
rect 35084 13132 35252 13134
rect 35196 13122 35252 13132
rect 35532 13188 35588 13198
rect 35644 13188 35700 18172
rect 35868 17666 35924 18956
rect 36316 18946 36372 18956
rect 36988 19012 37044 19022
rect 35868 17614 35870 17666
rect 35922 17614 35924 17666
rect 35868 17602 35924 17614
rect 36988 18340 37044 18956
rect 37548 19012 37604 19022
rect 37548 18918 37604 18956
rect 38220 19012 38276 19022
rect 38220 18676 38276 18956
rect 38668 18676 38724 19852
rect 39788 19814 39844 19852
rect 42140 19908 42196 19918
rect 42140 19814 42196 19852
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 38220 18674 38724 18676
rect 38220 18622 38670 18674
rect 38722 18622 38724 18674
rect 38220 18620 38724 18622
rect 38220 18450 38276 18620
rect 38220 18398 38222 18450
rect 38274 18398 38276 18450
rect 38220 18386 38276 18398
rect 36092 17556 36148 17566
rect 36092 17462 36148 17500
rect 36876 17108 36932 17118
rect 36988 17108 37044 18284
rect 37436 18338 37492 18350
rect 37436 18286 37438 18338
rect 37490 18286 37492 18338
rect 37436 17556 37492 18286
rect 37436 17490 37492 17500
rect 36876 17106 37044 17108
rect 36876 17054 36878 17106
rect 36930 17054 37044 17106
rect 36876 17052 37044 17054
rect 36876 17042 36932 17052
rect 36428 16770 36484 16782
rect 36428 16718 36430 16770
rect 36482 16718 36484 16770
rect 36428 16660 36484 16718
rect 36428 16594 36484 16604
rect 35868 16100 35924 16110
rect 35868 16098 36260 16100
rect 35868 16046 35870 16098
rect 35922 16046 36260 16098
rect 35868 16044 36260 16046
rect 35868 16034 35924 16044
rect 36092 15876 36148 15886
rect 36092 15782 36148 15820
rect 36204 14754 36260 16044
rect 37548 15876 37604 15886
rect 37548 15426 37604 15820
rect 38668 15540 38724 18620
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 38780 15540 38836 15550
rect 37548 15374 37550 15426
rect 37602 15374 37604 15426
rect 37548 15362 37604 15374
rect 38556 15538 39172 15540
rect 38556 15486 38782 15538
rect 38834 15486 39172 15538
rect 38556 15484 39172 15486
rect 38332 15316 38388 15326
rect 38556 15316 38612 15484
rect 38780 15474 38836 15484
rect 38332 15314 38612 15316
rect 38332 15262 38334 15314
rect 38386 15262 38612 15314
rect 38332 15260 38612 15262
rect 38332 15250 38388 15260
rect 36204 14702 36206 14754
rect 36258 14702 36260 14754
rect 36204 14690 36260 14702
rect 35868 14530 35924 14542
rect 35868 14478 35870 14530
rect 35922 14478 35924 14530
rect 35532 13186 35700 13188
rect 35532 13134 35534 13186
rect 35586 13134 35700 13186
rect 35532 13132 35700 13134
rect 35756 14084 35812 14094
rect 35532 13122 35588 13132
rect 35756 12850 35812 14028
rect 35756 12798 35758 12850
rect 35810 12798 35812 12850
rect 35756 12786 35812 12798
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34524 11666 34580 11676
rect 35532 11620 35588 11630
rect 35868 11620 35924 14478
rect 36316 12850 36372 12862
rect 36316 12798 36318 12850
rect 36370 12798 36372 12850
rect 35980 12068 36036 12078
rect 35980 11974 36036 12012
rect 36316 12066 36372 12798
rect 39116 12404 39172 15484
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 39676 12404 39732 12414
rect 39116 12402 39732 12404
rect 39116 12350 39678 12402
rect 39730 12350 39732 12402
rect 39116 12348 39732 12350
rect 36316 12014 36318 12066
rect 36370 12014 36372 12066
rect 35588 11564 35924 11620
rect 35980 11844 36036 11854
rect 35532 11526 35588 11564
rect 34300 11230 34302 11282
rect 34354 11230 34356 11282
rect 34300 11218 34356 11230
rect 35756 11396 35812 11406
rect 35756 11282 35812 11340
rect 35756 11230 35758 11282
rect 35810 11230 35812 11282
rect 35756 11218 35812 11230
rect 35196 11172 35252 11182
rect 35196 11170 35700 11172
rect 35196 11118 35198 11170
rect 35250 11118 35700 11170
rect 35196 11116 35700 11118
rect 35196 11106 35252 11116
rect 35644 10722 35700 11116
rect 35980 10834 36036 11788
rect 36316 11282 36372 12014
rect 37100 12180 37156 12190
rect 37100 11506 37156 12124
rect 39116 12180 39172 12348
rect 39676 12338 39732 12348
rect 39116 12086 39172 12124
rect 38444 12066 38500 12078
rect 38444 12014 38446 12066
rect 38498 12014 38500 12066
rect 38444 11844 38500 12014
rect 38444 11778 38500 11788
rect 37100 11454 37102 11506
rect 37154 11454 37156 11506
rect 37100 11442 37156 11454
rect 36316 11230 36318 11282
rect 36370 11230 36372 11282
rect 36316 11218 36372 11230
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 35980 10782 35982 10834
rect 36034 10782 36036 10834
rect 35980 10770 36036 10782
rect 35644 10670 35646 10722
rect 35698 10670 35700 10722
rect 35644 10658 35700 10670
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 31388 9102 31390 9154
rect 31442 9102 31444 9154
rect 31388 9090 31444 9102
rect 32172 9266 33572 9268
rect 32172 9214 33182 9266
rect 33234 9214 33572 9266
rect 32172 9212 33572 9214
rect 32172 9042 32228 9212
rect 33180 9202 33236 9212
rect 32172 8990 32174 9042
rect 32226 8990 32228 9042
rect 32172 8978 32228 8990
rect 30716 8306 30772 8316
rect 31276 8306 31332 8316
rect 32844 8372 32900 8382
rect 32844 8278 32900 8316
rect 33516 8260 33572 9212
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 33628 8260 33684 8270
rect 34188 8260 34244 8270
rect 33516 8258 34244 8260
rect 33516 8206 33630 8258
rect 33682 8206 34190 8258
rect 34242 8206 34244 8258
rect 33516 8204 34244 8206
rect 33628 8194 33684 8204
rect 34188 8194 34244 8204
rect 27916 7534 27918 7586
rect 27970 7534 27972 7586
rect 27916 7522 27972 7534
rect 28588 7980 28868 8036
rect 27244 6636 27636 6692
rect 27244 6468 27300 6478
rect 27244 6466 27524 6468
rect 27244 6414 27246 6466
rect 27298 6414 27524 6466
rect 27244 6412 27524 6414
rect 27244 6402 27300 6412
rect 27132 5854 27134 5906
rect 27186 5854 27188 5906
rect 27132 5842 27188 5854
rect 27020 5796 27076 5806
rect 26684 4564 26740 4574
rect 26684 4338 26740 4508
rect 26684 4286 26686 4338
rect 26738 4286 26740 4338
rect 26684 4274 26740 4286
rect 26572 3726 26574 3778
rect 26626 3726 26628 3778
rect 26572 3714 26628 3726
rect 27020 3444 27076 5740
rect 27468 4450 27524 6412
rect 27468 4398 27470 4450
rect 27522 4398 27524 4450
rect 27468 4386 27524 4398
rect 27580 5906 27636 6636
rect 28588 6690 28644 7980
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 28588 6638 28590 6690
rect 28642 6638 28644 6690
rect 28588 6626 28644 6638
rect 28476 6578 28532 6590
rect 28476 6526 28478 6578
rect 28530 6526 28532 6578
rect 27580 5854 27582 5906
rect 27634 5854 27636 5906
rect 27580 4228 27636 5854
rect 27244 4172 27636 4228
rect 27916 6020 27972 6030
rect 28476 6020 28532 6526
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 27916 6018 28532 6020
rect 27916 5966 27918 6018
rect 27970 5966 28532 6018
rect 27916 5964 28532 5966
rect 27916 4228 27972 5964
rect 28252 5796 28308 5806
rect 28252 5234 28308 5740
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 28252 5182 28254 5234
rect 28306 5182 28308 5234
rect 28252 5170 28308 5182
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 27244 3554 27300 4172
rect 27916 4162 27972 4172
rect 29596 4228 29652 4238
rect 29596 4134 29652 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 27244 3502 27246 3554
rect 27298 3502 27300 3554
rect 27244 3490 27300 3502
rect 27132 3444 27188 3454
rect 27020 3442 27188 3444
rect 27020 3390 27134 3442
rect 27186 3390 27188 3442
rect 27020 3388 27188 3390
rect 27132 3378 27188 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
<< via2 >>
rect 4620 56306 4676 56308
rect 4620 56254 4622 56306
rect 4622 56254 4674 56306
rect 4674 56254 4676 56306
rect 4620 56252 4676 56254
rect 5516 56252 5572 56308
rect 5852 56194 5908 56196
rect 5852 56142 5854 56194
rect 5854 56142 5906 56194
rect 5906 56142 5908 56194
rect 5852 56140 5908 56142
rect 8428 56140 8484 56196
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 14812 56028 14868 56084
rect 4060 53788 4116 53844
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 3276 52780 3332 52836
rect 2492 51884 2548 51940
rect 2492 48748 2548 48804
rect 3612 51996 3668 52052
rect 3836 52946 3892 52948
rect 3836 52894 3838 52946
rect 3838 52894 3890 52946
rect 3890 52894 3892 52946
rect 3836 52892 3892 52894
rect 4508 52946 4564 52948
rect 4508 52894 4510 52946
rect 4510 52894 4562 52946
rect 4562 52894 4564 52946
rect 4508 52892 4564 52894
rect 4956 52892 5012 52948
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4396 52386 4452 52388
rect 4396 52334 4398 52386
rect 4398 52334 4450 52386
rect 4450 52334 4452 52386
rect 4396 52332 4452 52334
rect 4956 52220 5012 52276
rect 4396 51996 4452 52052
rect 4284 51938 4340 51940
rect 4284 51886 4286 51938
rect 4286 51886 4338 51938
rect 4338 51886 4340 51938
rect 4284 51884 4340 51886
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 3836 50764 3892 50820
rect 4620 50764 4676 50820
rect 4956 50652 5012 50708
rect 4060 50540 4116 50596
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4844 49420 4900 49476
rect 4684 49364 4740 49366
rect 3948 49084 4004 49140
rect 4732 49026 4788 49028
rect 4732 48974 4734 49026
rect 4734 48974 4786 49026
rect 4786 48974 4788 49026
rect 4732 48972 4788 48974
rect 4620 48802 4676 48804
rect 4620 48750 4622 48802
rect 4622 48750 4674 48802
rect 4674 48750 4676 48802
rect 4620 48748 4676 48750
rect 6188 52780 6244 52836
rect 6412 52332 6468 52388
rect 6300 52220 6356 52276
rect 6636 52162 6692 52164
rect 6636 52110 6638 52162
rect 6638 52110 6690 52162
rect 6690 52110 6692 52162
rect 6636 52108 6692 52110
rect 6748 52220 6804 52276
rect 8092 53058 8148 53060
rect 8092 53006 8094 53058
rect 8094 53006 8146 53058
rect 8146 53006 8148 53058
rect 8092 53004 8148 53006
rect 5964 50594 6020 50596
rect 5964 50542 5966 50594
rect 5966 50542 6018 50594
rect 6018 50542 6020 50594
rect 5964 50540 6020 50542
rect 4956 48860 5012 48916
rect 3052 48300 3108 48356
rect 4060 48242 4116 48244
rect 4060 48190 4062 48242
rect 4062 48190 4114 48242
rect 4114 48190 4116 48242
rect 4060 48188 4116 48190
rect 4956 48076 5012 48132
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 3388 46396 3444 46452
rect 1820 45948 1876 46004
rect 2268 45164 2324 45220
rect 2492 45218 2548 45220
rect 2492 45166 2494 45218
rect 2494 45166 2546 45218
rect 2546 45166 2548 45218
rect 2492 45164 2548 45166
rect 2716 45106 2772 45108
rect 2716 45054 2718 45106
rect 2718 45054 2770 45106
rect 2770 45054 2772 45106
rect 2716 45052 2772 45054
rect 3500 45164 3556 45220
rect 3388 44492 3444 44548
rect 3388 43484 3444 43540
rect 4284 46396 4340 46452
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4060 45164 4116 45220
rect 3948 45052 4004 45108
rect 4620 45052 4676 45108
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 3612 44044 3668 44100
rect 2828 41970 2884 41972
rect 2828 41918 2830 41970
rect 2830 41918 2882 41970
rect 2882 41918 2884 41970
rect 2828 41916 2884 41918
rect 5964 50316 6020 50372
rect 5628 48972 5684 49028
rect 5740 50092 5796 50148
rect 5740 49084 5796 49140
rect 5852 48860 5908 48916
rect 6748 50764 6804 50820
rect 6636 50706 6692 50708
rect 6636 50654 6638 50706
rect 6638 50654 6690 50706
rect 6690 50654 6692 50706
rect 6636 50652 6692 50654
rect 6188 50092 6244 50148
rect 6860 50594 6916 50596
rect 6860 50542 6862 50594
rect 6862 50542 6914 50594
rect 6914 50542 6916 50594
rect 6860 50540 6916 50542
rect 6076 49026 6132 49028
rect 6076 48974 6078 49026
rect 6078 48974 6130 49026
rect 6130 48974 6132 49026
rect 6076 48972 6132 48974
rect 5068 45948 5124 46004
rect 4956 45106 5012 45108
rect 4956 45054 4958 45106
rect 4958 45054 5010 45106
rect 5010 45054 5012 45106
rect 4956 45052 5012 45054
rect 5068 44098 5124 44100
rect 5068 44046 5070 44098
rect 5070 44046 5122 44098
rect 5122 44046 5124 44098
rect 5068 44044 5124 44046
rect 4620 43708 4676 43764
rect 4956 43708 5012 43764
rect 4732 43372 4788 43428
rect 4844 43596 4900 43652
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 6524 48748 6580 48804
rect 7532 52332 7588 52388
rect 7196 52162 7252 52164
rect 7196 52110 7198 52162
rect 7198 52110 7250 52162
rect 7250 52110 7252 52162
rect 7196 52108 7252 52110
rect 8540 53004 8596 53060
rect 7420 50370 7476 50372
rect 7420 50318 7422 50370
rect 7422 50318 7474 50370
rect 7474 50318 7476 50370
rect 7420 50316 7476 50318
rect 6972 48300 7028 48356
rect 7084 48860 7140 48916
rect 7644 48914 7700 48916
rect 7644 48862 7646 48914
rect 7646 48862 7698 48914
rect 7698 48862 7700 48914
rect 7644 48860 7700 48862
rect 7196 48748 7252 48804
rect 15148 55916 15204 55972
rect 15596 57036 15652 57092
rect 15708 56252 15764 56308
rect 9212 54460 9268 54516
rect 9996 54460 10052 54516
rect 9324 53788 9380 53844
rect 9212 52050 9268 52052
rect 9212 51998 9214 52050
rect 9214 51998 9266 52050
rect 9266 51998 9268 52050
rect 9212 51996 9268 51998
rect 8764 51100 8820 51156
rect 12124 54514 12180 54516
rect 12124 54462 12126 54514
rect 12126 54462 12178 54514
rect 12178 54462 12180 54514
rect 12124 54460 12180 54462
rect 17500 57036 17556 57092
rect 17052 55916 17108 55972
rect 16492 55356 16548 55412
rect 16604 55244 16660 55300
rect 16828 55186 16884 55188
rect 16828 55134 16830 55186
rect 16830 55134 16882 55186
rect 16882 55134 16884 55186
rect 16828 55132 16884 55134
rect 12908 53900 12964 53956
rect 10668 53788 10724 53844
rect 9548 53004 9604 53060
rect 11452 52946 11508 52948
rect 11452 52894 11454 52946
rect 11454 52894 11506 52946
rect 11506 52894 11508 52946
rect 11452 52892 11508 52894
rect 10892 52834 10948 52836
rect 10892 52782 10894 52834
rect 10894 52782 10946 52834
rect 10946 52782 10948 52834
rect 10892 52780 10948 52782
rect 12012 52834 12068 52836
rect 12012 52782 12014 52834
rect 12014 52782 12066 52834
rect 12066 52782 12068 52834
rect 12012 52780 12068 52782
rect 10332 51436 10388 51492
rect 11564 52220 11620 52276
rect 11340 51436 11396 51492
rect 10108 51154 10164 51156
rect 10108 51102 10110 51154
rect 10110 51102 10162 51154
rect 10162 51102 10164 51154
rect 10108 51100 10164 51102
rect 10220 50988 10276 51044
rect 9996 50428 10052 50484
rect 8652 48972 8708 49028
rect 7868 48354 7924 48356
rect 7868 48302 7870 48354
rect 7870 48302 7922 48354
rect 7922 48302 7924 48354
rect 7868 48300 7924 48302
rect 6412 46620 6468 46676
rect 5852 45778 5908 45780
rect 5852 45726 5854 45778
rect 5854 45726 5906 45778
rect 5906 45726 5908 45778
rect 5852 45724 5908 45726
rect 5292 44044 5348 44100
rect 5628 43708 5684 43764
rect 5516 43538 5572 43540
rect 5516 43486 5518 43538
rect 5518 43486 5570 43538
rect 5570 43486 5572 43538
rect 5516 43484 5572 43486
rect 3724 41916 3780 41972
rect 3164 41858 3220 41860
rect 3164 41806 3166 41858
rect 3166 41806 3218 41858
rect 3218 41806 3220 41858
rect 3164 41804 3220 41806
rect 2492 40572 2548 40628
rect 4060 41970 4116 41972
rect 4060 41918 4062 41970
rect 4062 41918 4114 41970
rect 4114 41918 4116 41970
rect 4060 41916 4116 41918
rect 6412 45164 6468 45220
rect 6524 45724 6580 45780
rect 5964 44380 6020 44436
rect 5628 43372 5684 43428
rect 5852 43314 5908 43316
rect 5852 43262 5854 43314
rect 5854 43262 5906 43314
rect 5906 43262 5908 43314
rect 5852 43260 5908 43262
rect 7532 46620 7588 46676
rect 6636 43538 6692 43540
rect 6636 43486 6638 43538
rect 6638 43486 6690 43538
rect 6690 43486 6692 43538
rect 6636 43484 6692 43486
rect 7308 44380 7364 44436
rect 8092 48242 8148 48244
rect 8092 48190 8094 48242
rect 8094 48190 8146 48242
rect 8146 48190 8148 48242
rect 8092 48188 8148 48190
rect 8652 48242 8708 48244
rect 8652 48190 8654 48242
rect 8654 48190 8706 48242
rect 8706 48190 8708 48242
rect 8652 48188 8708 48190
rect 8764 48130 8820 48132
rect 8764 48078 8766 48130
rect 8766 48078 8818 48130
rect 8818 48078 8820 48130
rect 8764 48076 8820 48078
rect 8988 48018 9044 48020
rect 8988 47966 8990 48018
rect 8990 47966 9042 48018
rect 9042 47966 9044 48018
rect 8988 47964 9044 47966
rect 8876 47570 8932 47572
rect 8876 47518 8878 47570
rect 8878 47518 8930 47570
rect 8930 47518 8932 47570
rect 8876 47516 8932 47518
rect 5628 42642 5684 42644
rect 5628 42590 5630 42642
rect 5630 42590 5682 42642
rect 5682 42590 5684 42642
rect 5628 42588 5684 42590
rect 4732 41970 4788 41972
rect 4732 41918 4734 41970
rect 4734 41918 4786 41970
rect 4786 41918 4788 41970
rect 4732 41916 4788 41918
rect 3948 41858 4004 41860
rect 3948 41806 3950 41858
rect 3950 41806 4002 41858
rect 4002 41806 4004 41858
rect 3948 41804 4004 41806
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5292 41970 5348 41972
rect 5292 41918 5294 41970
rect 5294 41918 5346 41970
rect 5346 41918 5348 41970
rect 5292 41916 5348 41918
rect 5964 41916 6020 41972
rect 4508 40626 4564 40628
rect 4508 40574 4510 40626
rect 4510 40574 4562 40626
rect 4562 40574 4564 40626
rect 4508 40572 4564 40574
rect 4844 40348 4900 40404
rect 4620 40290 4676 40292
rect 4620 40238 4622 40290
rect 4622 40238 4674 40290
rect 4674 40238 4676 40290
rect 4620 40236 4676 40238
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5628 41356 5684 41412
rect 6188 41186 6244 41188
rect 6188 41134 6190 41186
rect 6190 41134 6242 41186
rect 6242 41134 6244 41186
rect 6188 41132 6244 41134
rect 5852 41020 5908 41076
rect 5516 40236 5572 40292
rect 5964 40236 6020 40292
rect 3388 39228 3444 39284
rect 1820 38050 1876 38052
rect 1820 37998 1822 38050
rect 1822 37998 1874 38050
rect 1874 37998 1876 38050
rect 1820 37996 1876 37998
rect 2492 37938 2548 37940
rect 2492 37886 2494 37938
rect 2494 37886 2546 37938
rect 2546 37886 2548 37938
rect 2492 37884 2548 37886
rect 3500 37884 3556 37940
rect 3724 37436 3780 37492
rect 3388 37266 3444 37268
rect 3388 37214 3390 37266
rect 3390 37214 3442 37266
rect 3442 37214 3444 37266
rect 3388 37212 3444 37214
rect 4284 39394 4340 39396
rect 4284 39342 4286 39394
rect 4286 39342 4338 39394
rect 4338 39342 4340 39394
rect 4284 39340 4340 39342
rect 4732 39228 4788 39284
rect 4844 38892 4900 38948
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4620 38162 4676 38164
rect 4620 38110 4622 38162
rect 4622 38110 4674 38162
rect 4674 38110 4676 38162
rect 4620 38108 4676 38110
rect 4620 37436 4676 37492
rect 5068 37826 5124 37828
rect 5068 37774 5070 37826
rect 5070 37774 5122 37826
rect 5122 37774 5124 37826
rect 5068 37772 5124 37774
rect 5180 39340 5236 39396
rect 6412 42588 6468 42644
rect 8652 45218 8708 45220
rect 8652 45166 8654 45218
rect 8654 45166 8706 45218
rect 8706 45166 8708 45218
rect 8652 45164 8708 45166
rect 8764 44492 8820 44548
rect 8540 44434 8596 44436
rect 8540 44382 8542 44434
rect 8542 44382 8594 44434
rect 8594 44382 8596 44434
rect 8540 44380 8596 44382
rect 8988 43820 9044 43876
rect 7420 43596 7476 43652
rect 9100 43484 9156 43540
rect 7532 43260 7588 43316
rect 6860 41410 6916 41412
rect 6860 41358 6862 41410
rect 6862 41358 6914 41410
rect 6914 41358 6916 41410
rect 6860 41356 6916 41358
rect 6972 41186 7028 41188
rect 6972 41134 6974 41186
rect 6974 41134 7026 41186
rect 7026 41134 7028 41186
rect 6972 41132 7028 41134
rect 6636 41020 6692 41076
rect 7084 41074 7140 41076
rect 7084 41022 7086 41074
rect 7086 41022 7138 41074
rect 7138 41022 7140 41074
rect 7084 41020 7140 41022
rect 6524 40460 6580 40516
rect 6412 40348 6468 40404
rect 6076 39394 6132 39396
rect 6076 39342 6078 39394
rect 6078 39342 6130 39394
rect 6130 39342 6132 39394
rect 6076 39340 6132 39342
rect 5292 38946 5348 38948
rect 5292 38894 5294 38946
rect 5294 38894 5346 38946
rect 5346 38894 5348 38946
rect 5292 38892 5348 38894
rect 5516 38892 5572 38948
rect 6188 38892 6244 38948
rect 6524 39004 6580 39060
rect 6860 39340 6916 39396
rect 5180 37490 5236 37492
rect 5180 37438 5182 37490
rect 5182 37438 5234 37490
rect 5234 37438 5236 37490
rect 5180 37436 5236 37438
rect 6860 38780 6916 38836
rect 6972 39228 7028 39284
rect 8652 43260 8708 43316
rect 8876 42028 8932 42084
rect 8764 41970 8820 41972
rect 8764 41918 8766 41970
rect 8766 41918 8818 41970
rect 8818 41918 8820 41970
rect 8764 41916 8820 41918
rect 9100 41916 9156 41972
rect 8988 40626 9044 40628
rect 8988 40574 8990 40626
rect 8990 40574 9042 40626
rect 9042 40574 9044 40626
rect 8988 40572 9044 40574
rect 7756 40514 7812 40516
rect 7756 40462 7758 40514
rect 7758 40462 7810 40514
rect 7810 40462 7812 40514
rect 7756 40460 7812 40462
rect 7532 39004 7588 39060
rect 7420 38834 7476 38836
rect 7420 38782 7422 38834
rect 7422 38782 7474 38834
rect 7474 38782 7476 38834
rect 7420 38780 7476 38782
rect 8764 38780 8820 38836
rect 5516 38108 5572 38164
rect 5964 37772 6020 37828
rect 3836 37212 3892 37268
rect 4284 37266 4340 37268
rect 4284 37214 4286 37266
rect 4286 37214 4338 37266
rect 4338 37214 4340 37266
rect 4284 37212 4340 37214
rect 8428 37772 8484 37828
rect 6524 37212 6580 37268
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4284 29260 4340 29316
rect 5740 29260 5796 29316
rect 8876 37772 8932 37828
rect 9212 37826 9268 37828
rect 9212 37774 9214 37826
rect 9214 37774 9266 37826
rect 9266 37774 9268 37826
rect 9212 37772 9268 37774
rect 11676 51996 11732 52052
rect 12796 52892 12852 52948
rect 12460 52220 12516 52276
rect 12572 52332 12628 52388
rect 11340 51154 11396 51156
rect 11340 51102 11342 51154
rect 11342 51102 11394 51154
rect 11394 51102 11396 51154
rect 11340 51100 11396 51102
rect 10892 50428 10948 50484
rect 11788 50482 11844 50484
rect 11788 50430 11790 50482
rect 11790 50430 11842 50482
rect 11842 50430 11844 50482
rect 11788 50428 11844 50430
rect 11228 49644 11284 49700
rect 11676 49698 11732 49700
rect 11676 49646 11678 49698
rect 11678 49646 11730 49698
rect 11730 49646 11732 49698
rect 11676 49644 11732 49646
rect 9772 48860 9828 48916
rect 9772 48242 9828 48244
rect 9772 48190 9774 48242
rect 9774 48190 9826 48242
rect 9826 48190 9828 48242
rect 9772 48188 9828 48190
rect 11788 48972 11844 49028
rect 9884 48076 9940 48132
rect 11340 48412 11396 48468
rect 10892 48188 10948 48244
rect 9660 47516 9716 47572
rect 9996 48018 10052 48020
rect 9996 47966 9998 48018
rect 9998 47966 10050 48018
rect 10050 47966 10052 48018
rect 9996 47964 10052 47966
rect 11676 48300 11732 48356
rect 10556 46060 10612 46116
rect 10108 44546 10164 44548
rect 10108 44494 10110 44546
rect 10110 44494 10162 44546
rect 10162 44494 10164 44546
rect 10108 44492 10164 44494
rect 10556 45164 10612 45220
rect 10892 46060 10948 46116
rect 11564 46674 11620 46676
rect 11564 46622 11566 46674
rect 11566 46622 11618 46674
rect 11618 46622 11620 46674
rect 11564 46620 11620 46622
rect 12012 51154 12068 51156
rect 12012 51102 12014 51154
rect 12014 51102 12066 51154
rect 12066 51102 12068 51154
rect 12012 51100 12068 51102
rect 12908 50652 12964 50708
rect 13132 52108 13188 52164
rect 13468 53954 13524 53956
rect 13468 53902 13470 53954
rect 13470 53902 13522 53954
rect 13522 53902 13524 53954
rect 13468 53900 13524 53902
rect 13580 53842 13636 53844
rect 13580 53790 13582 53842
rect 13582 53790 13634 53842
rect 13634 53790 13636 53842
rect 13580 53788 13636 53790
rect 13468 52780 13524 52836
rect 12572 50594 12628 50596
rect 12572 50542 12574 50594
rect 12574 50542 12626 50594
rect 12626 50542 12628 50594
rect 12572 50540 12628 50542
rect 12348 50482 12404 50484
rect 12348 50430 12350 50482
rect 12350 50430 12402 50482
rect 12402 50430 12404 50482
rect 12348 50428 12404 50430
rect 12572 50316 12628 50372
rect 12236 49922 12292 49924
rect 12236 49870 12238 49922
rect 12238 49870 12290 49922
rect 12290 49870 12292 49922
rect 12236 49868 12292 49870
rect 11900 48860 11956 48916
rect 12124 48972 12180 49028
rect 12348 48018 12404 48020
rect 12348 47966 12350 48018
rect 12350 47966 12402 48018
rect 12402 47966 12404 48018
rect 12348 47964 12404 47966
rect 12124 47516 12180 47572
rect 11788 46284 11844 46340
rect 11228 45948 11284 46004
rect 10668 44828 10724 44884
rect 11004 44492 11060 44548
rect 10220 44434 10276 44436
rect 10220 44382 10222 44434
rect 10222 44382 10274 44434
rect 10274 44382 10276 44434
rect 10220 44380 10276 44382
rect 10332 43820 10388 43876
rect 9548 43596 9604 43652
rect 10220 43372 10276 43428
rect 10220 43036 10276 43092
rect 9660 41916 9716 41972
rect 9548 40572 9604 40628
rect 9660 38332 9716 38388
rect 10332 40514 10388 40516
rect 10332 40462 10334 40514
rect 10334 40462 10386 40514
rect 10386 40462 10388 40514
rect 10332 40460 10388 40462
rect 10108 37996 10164 38052
rect 11116 45052 11172 45108
rect 10668 44322 10724 44324
rect 10668 44270 10670 44322
rect 10670 44270 10722 44322
rect 10722 44270 10724 44322
rect 10668 44268 10724 44270
rect 11228 44940 11284 44996
rect 10892 43650 10948 43652
rect 10892 43598 10894 43650
rect 10894 43598 10946 43650
rect 10946 43598 10948 43650
rect 10892 43596 10948 43598
rect 11116 43820 11172 43876
rect 11788 44994 11844 44996
rect 11788 44942 11790 44994
rect 11790 44942 11842 44994
rect 11842 44942 11844 44994
rect 11788 44940 11844 44942
rect 11452 44492 11508 44548
rect 11788 44434 11844 44436
rect 11788 44382 11790 44434
rect 11790 44382 11842 44434
rect 11842 44382 11844 44434
rect 11788 44380 11844 44382
rect 11228 43650 11284 43652
rect 11228 43598 11230 43650
rect 11230 43598 11282 43650
rect 11282 43598 11284 43650
rect 11228 43596 11284 43598
rect 11676 44044 11732 44100
rect 11452 43148 11508 43204
rect 11788 43820 11844 43876
rect 11676 43314 11732 43316
rect 11676 43262 11678 43314
rect 11678 43262 11730 43314
rect 11730 43262 11732 43314
rect 11676 43260 11732 43262
rect 11452 41916 11508 41972
rect 13692 52444 13748 52500
rect 13804 52162 13860 52164
rect 13804 52110 13806 52162
rect 13806 52110 13858 52162
rect 13858 52110 13860 52162
rect 13804 52108 13860 52110
rect 13916 52780 13972 52836
rect 14812 52332 14868 52388
rect 16268 54236 16324 54292
rect 16492 53900 16548 53956
rect 16828 53506 16884 53508
rect 16828 53454 16830 53506
rect 16830 53454 16882 53506
rect 16882 53454 16884 53506
rect 16828 53452 16884 53454
rect 13692 50988 13748 51044
rect 13468 50652 13524 50708
rect 13132 49868 13188 49924
rect 12908 49756 12964 49812
rect 13244 48748 13300 48804
rect 12908 48188 12964 48244
rect 12684 47740 12740 47796
rect 14028 51378 14084 51380
rect 14028 51326 14030 51378
rect 14030 51326 14082 51378
rect 14082 51326 14084 51378
rect 14028 51324 14084 51326
rect 14364 51324 14420 51380
rect 14476 51436 14532 51492
rect 14364 50540 14420 50596
rect 13916 50316 13972 50372
rect 13804 49756 13860 49812
rect 13916 49644 13972 49700
rect 13356 47964 13412 48020
rect 13580 47682 13636 47684
rect 13580 47630 13582 47682
rect 13582 47630 13634 47682
rect 13634 47630 13636 47682
rect 13580 47628 13636 47630
rect 12572 47292 12628 47348
rect 13468 47068 13524 47124
rect 12908 46956 12964 47012
rect 12460 46060 12516 46116
rect 13580 46956 13636 47012
rect 13132 46674 13188 46676
rect 13132 46622 13134 46674
rect 13134 46622 13186 46674
rect 13186 46622 13188 46674
rect 13132 46620 13188 46622
rect 13356 46620 13412 46676
rect 12012 45106 12068 45108
rect 12012 45054 12014 45106
rect 12014 45054 12066 45106
rect 12066 45054 12068 45106
rect 12012 45052 12068 45054
rect 12572 45052 12628 45108
rect 12572 44492 12628 44548
rect 12908 44940 12964 44996
rect 12012 44044 12068 44100
rect 12348 44098 12404 44100
rect 12348 44046 12350 44098
rect 12350 44046 12402 44098
rect 12402 44046 12404 44098
rect 12348 44044 12404 44046
rect 13468 44380 13524 44436
rect 13244 44156 13300 44212
rect 13020 43932 13076 43988
rect 12684 43148 12740 43204
rect 13132 43538 13188 43540
rect 13132 43486 13134 43538
rect 13134 43486 13186 43538
rect 13186 43486 13188 43538
rect 13132 43484 13188 43486
rect 12796 42754 12852 42756
rect 12796 42702 12798 42754
rect 12798 42702 12850 42754
rect 12850 42702 12852 42754
rect 12796 42700 12852 42702
rect 12012 42530 12068 42532
rect 12012 42478 12014 42530
rect 12014 42478 12066 42530
rect 12066 42478 12068 42530
rect 12012 42476 12068 42478
rect 13356 43596 13412 43652
rect 13356 42476 13412 42532
rect 14140 47740 14196 47796
rect 13916 47180 13972 47236
rect 13692 46508 13748 46564
rect 14140 47346 14196 47348
rect 14140 47294 14142 47346
rect 14142 47294 14194 47346
rect 14194 47294 14196 47346
rect 14140 47292 14196 47294
rect 14140 47068 14196 47124
rect 14364 49810 14420 49812
rect 14364 49758 14366 49810
rect 14366 49758 14418 49810
rect 14418 49758 14420 49810
rect 14364 49756 14420 49758
rect 14364 46956 14420 47012
rect 15708 52220 15764 52276
rect 15484 52162 15540 52164
rect 15484 52110 15486 52162
rect 15486 52110 15538 52162
rect 15538 52110 15540 52162
rect 15484 52108 15540 52110
rect 15372 51490 15428 51492
rect 15372 51438 15374 51490
rect 15374 51438 15426 51490
rect 15426 51438 15428 51490
rect 15372 51436 15428 51438
rect 15596 51378 15652 51380
rect 15596 51326 15598 51378
rect 15598 51326 15650 51378
rect 15650 51326 15652 51378
rect 15596 51324 15652 51326
rect 15260 51212 15316 51268
rect 15148 50764 15204 50820
rect 15036 50594 15092 50596
rect 15036 50542 15038 50594
rect 15038 50542 15090 50594
rect 15090 50542 15092 50594
rect 15036 50540 15092 50542
rect 14924 50482 14980 50484
rect 14924 50430 14926 50482
rect 14926 50430 14978 50482
rect 14978 50430 14980 50482
rect 14924 50428 14980 50430
rect 14812 50316 14868 50372
rect 14812 49586 14868 49588
rect 14812 49534 14814 49586
rect 14814 49534 14866 49586
rect 14866 49534 14868 49586
rect 14812 49532 14868 49534
rect 15932 52444 15988 52500
rect 16156 51324 16212 51380
rect 16044 51266 16100 51268
rect 16044 51214 16046 51266
rect 16046 51214 16098 51266
rect 16098 51214 16100 51266
rect 16044 51212 16100 51214
rect 14924 48860 14980 48916
rect 15148 48412 15204 48468
rect 15260 48748 15316 48804
rect 14700 48242 14756 48244
rect 14700 48190 14702 48242
rect 14702 48190 14754 48242
rect 14754 48190 14756 48242
rect 14700 48188 14756 48190
rect 14588 47740 14644 47796
rect 14476 46508 14532 46564
rect 14588 46844 14644 46900
rect 14476 45388 14532 45444
rect 14700 45724 14756 45780
rect 14364 45106 14420 45108
rect 14364 45054 14366 45106
rect 14366 45054 14418 45106
rect 14418 45054 14420 45106
rect 14364 45052 14420 45054
rect 13692 44322 13748 44324
rect 13692 44270 13694 44322
rect 13694 44270 13746 44322
rect 13746 44270 13748 44322
rect 13692 44268 13748 44270
rect 13804 44098 13860 44100
rect 13804 44046 13806 44098
rect 13806 44046 13858 44098
rect 13858 44046 13860 44098
rect 13804 44044 13860 44046
rect 14476 44322 14532 44324
rect 14476 44270 14478 44322
rect 14478 44270 14530 44322
rect 14530 44270 14532 44322
rect 14476 44268 14532 44270
rect 14140 44156 14196 44212
rect 14364 44156 14420 44212
rect 14028 43708 14084 43764
rect 13692 43538 13748 43540
rect 13692 43486 13694 43538
rect 13694 43486 13746 43538
rect 13746 43486 13748 43538
rect 13692 43484 13748 43486
rect 13692 43148 13748 43204
rect 14476 43932 14532 43988
rect 14700 43820 14756 43876
rect 15148 46172 15204 46228
rect 15036 46002 15092 46004
rect 15036 45950 15038 46002
rect 15038 45950 15090 46002
rect 15090 45950 15092 46002
rect 15036 45948 15092 45950
rect 15036 45388 15092 45444
rect 15820 49586 15876 49588
rect 15820 49534 15822 49586
rect 15822 49534 15874 49586
rect 15874 49534 15876 49586
rect 15820 49532 15876 49534
rect 15596 48354 15652 48356
rect 15596 48302 15598 48354
rect 15598 48302 15650 48354
rect 15650 48302 15652 48354
rect 15596 48300 15652 48302
rect 15484 45948 15540 46004
rect 14924 44210 14980 44212
rect 14924 44158 14926 44210
rect 14926 44158 14978 44210
rect 14978 44158 14980 44210
rect 14924 44156 14980 44158
rect 15484 44210 15540 44212
rect 15484 44158 15486 44210
rect 15486 44158 15538 44210
rect 15538 44158 15540 44210
rect 15484 44156 15540 44158
rect 14028 42812 14084 42868
rect 14812 42812 14868 42868
rect 12236 41970 12292 41972
rect 12236 41918 12238 41970
rect 12238 41918 12290 41970
rect 12290 41918 12292 41970
rect 12236 41916 12292 41918
rect 13468 41804 13524 41860
rect 13356 41580 13412 41636
rect 11452 39730 11508 39732
rect 11452 39678 11454 39730
rect 11454 39678 11506 39730
rect 11506 39678 11508 39730
rect 11452 39676 11508 39678
rect 12572 40962 12628 40964
rect 12572 40910 12574 40962
rect 12574 40910 12626 40962
rect 12626 40910 12628 40962
rect 12572 40908 12628 40910
rect 12236 39676 12292 39732
rect 13132 40348 13188 40404
rect 12684 39730 12740 39732
rect 12684 39678 12686 39730
rect 12686 39678 12738 39730
rect 12738 39678 12740 39730
rect 12684 39676 12740 39678
rect 11900 39004 11956 39060
rect 11788 37938 11844 37940
rect 11788 37886 11790 37938
rect 11790 37886 11842 37938
rect 11842 37886 11844 37938
rect 11788 37884 11844 37886
rect 13020 39506 13076 39508
rect 13020 39454 13022 39506
rect 13022 39454 13074 39506
rect 13074 39454 13076 39506
rect 13020 39452 13076 39454
rect 12684 38332 12740 38388
rect 11116 37266 11172 37268
rect 11116 37214 11118 37266
rect 11118 37214 11170 37266
rect 11170 37214 11172 37266
rect 11116 37212 11172 37214
rect 12572 37212 12628 37268
rect 13244 35308 13300 35364
rect 12684 35084 12740 35140
rect 10556 34860 10612 34916
rect 9436 32732 9492 32788
rect 11788 33068 11844 33124
rect 13804 42028 13860 42084
rect 13580 40460 13636 40516
rect 14140 42754 14196 42756
rect 14140 42702 14142 42754
rect 14142 42702 14194 42754
rect 14194 42702 14196 42754
rect 14140 42700 14196 42702
rect 14364 42194 14420 42196
rect 14364 42142 14366 42194
rect 14366 42142 14418 42194
rect 14418 42142 14420 42194
rect 14364 42140 14420 42142
rect 14476 42082 14532 42084
rect 14476 42030 14478 42082
rect 14478 42030 14530 42082
rect 14530 42030 14532 42082
rect 14476 42028 14532 42030
rect 14924 42082 14980 42084
rect 14924 42030 14926 42082
rect 14926 42030 14978 42082
rect 14978 42030 14980 42082
rect 14924 42028 14980 42030
rect 15148 43820 15204 43876
rect 13916 41580 13972 41636
rect 14252 41298 14308 41300
rect 14252 41246 14254 41298
rect 14254 41246 14306 41298
rect 14306 41246 14308 41298
rect 14252 41244 14308 41246
rect 14364 40684 14420 40740
rect 13916 40626 13972 40628
rect 13916 40574 13918 40626
rect 13918 40574 13970 40626
rect 13970 40574 13972 40626
rect 13916 40572 13972 40574
rect 14812 41746 14868 41748
rect 14812 41694 14814 41746
rect 14814 41694 14866 41746
rect 14866 41694 14868 41746
rect 14812 41692 14868 41694
rect 14924 41020 14980 41076
rect 14812 40684 14868 40740
rect 13916 40402 13972 40404
rect 13916 40350 13918 40402
rect 13918 40350 13970 40402
rect 13970 40350 13972 40402
rect 13916 40348 13972 40350
rect 13692 39900 13748 39956
rect 13916 39340 13972 39396
rect 13804 38946 13860 38948
rect 13804 38894 13806 38946
rect 13806 38894 13858 38946
rect 13858 38894 13860 38946
rect 13804 38892 13860 38894
rect 13692 37212 13748 37268
rect 14588 39340 14644 39396
rect 14700 39228 14756 39284
rect 15260 43596 15316 43652
rect 15708 46956 15764 47012
rect 15820 46450 15876 46452
rect 15820 46398 15822 46450
rect 15822 46398 15874 46450
rect 15874 46398 15876 46450
rect 15820 46396 15876 46398
rect 16828 51100 16884 51156
rect 16604 50764 16660 50820
rect 16492 49868 16548 49924
rect 16380 49810 16436 49812
rect 16380 49758 16382 49810
rect 16382 49758 16434 49810
rect 16434 49758 16436 49810
rect 16380 49756 16436 49758
rect 16604 49026 16660 49028
rect 16604 48974 16606 49026
rect 16606 48974 16658 49026
rect 16658 48974 16660 49026
rect 16604 48972 16660 48974
rect 16604 48748 16660 48804
rect 16492 47628 16548 47684
rect 16492 47292 16548 47348
rect 16044 46956 16100 47012
rect 15932 46172 15988 46228
rect 15708 45778 15764 45780
rect 15708 45726 15710 45778
rect 15710 45726 15762 45778
rect 15762 45726 15764 45778
rect 15708 45724 15764 45726
rect 16044 45666 16100 45668
rect 16044 45614 16046 45666
rect 16046 45614 16098 45666
rect 16098 45614 16100 45666
rect 16044 45612 16100 45614
rect 16268 46786 16324 46788
rect 16268 46734 16270 46786
rect 16270 46734 16322 46786
rect 16322 46734 16324 46786
rect 16268 46732 16324 46734
rect 16380 46508 16436 46564
rect 16828 48636 16884 48692
rect 16828 47852 16884 47908
rect 16716 47404 16772 47460
rect 16716 47180 16772 47236
rect 16716 46732 16772 46788
rect 16604 46284 16660 46340
rect 17948 55468 18004 55524
rect 18508 55410 18564 55412
rect 18508 55358 18510 55410
rect 18510 55358 18562 55410
rect 18562 55358 18564 55410
rect 18508 55356 18564 55358
rect 17612 55244 17668 55300
rect 17388 54460 17444 54516
rect 17164 53954 17220 53956
rect 17164 53902 17166 53954
rect 17166 53902 17218 53954
rect 17218 53902 17220 53954
rect 17164 53900 17220 53902
rect 18284 55244 18340 55300
rect 17836 55020 17892 55076
rect 17948 54684 18004 54740
rect 17500 54236 17556 54292
rect 18284 54236 18340 54292
rect 17836 53452 17892 53508
rect 17724 52834 17780 52836
rect 17724 52782 17726 52834
rect 17726 52782 17778 52834
rect 17778 52782 17780 52834
rect 17724 52780 17780 52782
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19180 55522 19236 55524
rect 19180 55470 19182 55522
rect 19182 55470 19234 55522
rect 19234 55470 19236 55522
rect 19180 55468 19236 55470
rect 19852 55356 19908 55412
rect 18956 55244 19012 55300
rect 20188 55244 20244 55300
rect 19628 55132 19684 55188
rect 18844 55074 18900 55076
rect 18844 55022 18846 55074
rect 18846 55022 18898 55074
rect 18898 55022 18900 55074
rect 18844 55020 18900 55022
rect 19180 54738 19236 54740
rect 19180 54686 19182 54738
rect 19182 54686 19234 54738
rect 19234 54686 19236 54738
rect 19180 54684 19236 54686
rect 18620 53900 18676 53956
rect 18732 52834 18788 52836
rect 18732 52782 18734 52834
rect 18734 52782 18786 52834
rect 18786 52782 18788 52834
rect 18732 52780 18788 52782
rect 17948 52108 18004 52164
rect 17388 51490 17444 51492
rect 17388 51438 17390 51490
rect 17390 51438 17442 51490
rect 17442 51438 17444 51490
rect 17388 51436 17444 51438
rect 17612 51266 17668 51268
rect 17612 51214 17614 51266
rect 17614 51214 17666 51266
rect 17666 51214 17668 51266
rect 17612 51212 17668 51214
rect 17276 49868 17332 49924
rect 17164 49026 17220 49028
rect 17164 48974 17166 49026
rect 17166 48974 17218 49026
rect 17218 48974 17220 49026
rect 17164 48972 17220 48974
rect 17500 48466 17556 48468
rect 17500 48414 17502 48466
rect 17502 48414 17554 48466
rect 17554 48414 17556 48466
rect 17500 48412 17556 48414
rect 17276 48242 17332 48244
rect 17276 48190 17278 48242
rect 17278 48190 17330 48242
rect 17330 48190 17332 48242
rect 17276 48188 17332 48190
rect 17164 46956 17220 47012
rect 16492 46060 16548 46116
rect 17164 46114 17220 46116
rect 17164 46062 17166 46114
rect 17166 46062 17218 46114
rect 17218 46062 17220 46114
rect 17164 46060 17220 46062
rect 17052 45778 17108 45780
rect 17052 45726 17054 45778
rect 17054 45726 17106 45778
rect 17106 45726 17108 45778
rect 17052 45724 17108 45726
rect 15260 42140 15316 42196
rect 15372 42364 15428 42420
rect 15260 41692 15316 41748
rect 15596 41356 15652 41412
rect 15372 41132 15428 41188
rect 15484 41020 15540 41076
rect 15372 40908 15428 40964
rect 15260 40572 15316 40628
rect 15148 39228 15204 39284
rect 17164 45276 17220 45332
rect 17276 45052 17332 45108
rect 15932 44210 15988 44212
rect 15932 44158 15934 44210
rect 15934 44158 15986 44210
rect 15986 44158 15988 44210
rect 15932 44156 15988 44158
rect 16380 44828 16436 44884
rect 16268 43538 16324 43540
rect 16268 43486 16270 43538
rect 16270 43486 16322 43538
rect 16322 43486 16324 43538
rect 16268 43484 16324 43486
rect 16044 42978 16100 42980
rect 16044 42926 16046 42978
rect 16046 42926 16098 42978
rect 16098 42926 16100 42978
rect 16044 42924 16100 42926
rect 16268 42754 16324 42756
rect 16268 42702 16270 42754
rect 16270 42702 16322 42754
rect 16322 42702 16324 42754
rect 16268 42700 16324 42702
rect 16156 42588 16212 42644
rect 16044 42364 16100 42420
rect 17836 48412 17892 48468
rect 17948 48076 18004 48132
rect 17836 47852 17892 47908
rect 17724 46732 17780 46788
rect 17948 46674 18004 46676
rect 17948 46622 17950 46674
rect 17950 46622 18002 46674
rect 18002 46622 18004 46674
rect 17948 46620 18004 46622
rect 17388 44716 17444 44772
rect 17724 45890 17780 45892
rect 17724 45838 17726 45890
rect 17726 45838 17778 45890
rect 17778 45838 17780 45890
rect 17724 45836 17780 45838
rect 16716 43260 16772 43316
rect 16828 44604 16884 44660
rect 16604 42812 16660 42868
rect 16716 42588 16772 42644
rect 16268 41970 16324 41972
rect 16268 41918 16270 41970
rect 16270 41918 16322 41970
rect 16322 41918 16324 41970
rect 16268 41916 16324 41918
rect 16380 41858 16436 41860
rect 16380 41806 16382 41858
rect 16382 41806 16434 41858
rect 16434 41806 16436 41858
rect 16380 41804 16436 41806
rect 16268 41580 16324 41636
rect 16044 41356 16100 41412
rect 16156 41298 16212 41300
rect 16156 41246 16158 41298
rect 16158 41246 16210 41298
rect 16210 41246 16212 41298
rect 16156 41244 16212 41246
rect 15708 41020 15764 41076
rect 16156 41020 16212 41076
rect 15484 40460 15540 40516
rect 15372 40236 15428 40292
rect 15708 40626 15764 40628
rect 15708 40574 15710 40626
rect 15710 40574 15762 40626
rect 15762 40574 15764 40626
rect 15708 40572 15764 40574
rect 15596 40124 15652 40180
rect 15372 39842 15428 39844
rect 15372 39790 15374 39842
rect 15374 39790 15426 39842
rect 15426 39790 15428 39842
rect 15372 39788 15428 39790
rect 17276 44492 17332 44548
rect 17052 44434 17108 44436
rect 17052 44382 17054 44434
rect 17054 44382 17106 44434
rect 17106 44382 17108 44434
rect 17052 44380 17108 44382
rect 17612 45052 17668 45108
rect 17388 43708 17444 43764
rect 16940 43538 16996 43540
rect 16940 43486 16942 43538
rect 16942 43486 16994 43538
rect 16994 43486 16996 43538
rect 16940 43484 16996 43486
rect 17164 43372 17220 43428
rect 17500 43426 17556 43428
rect 17500 43374 17502 43426
rect 17502 43374 17554 43426
rect 17554 43374 17556 43426
rect 17500 43372 17556 43374
rect 17276 43260 17332 43316
rect 17724 44604 17780 44660
rect 17724 43820 17780 43876
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19516 54514 19572 54516
rect 19516 54462 19518 54514
rect 19518 54462 19570 54514
rect 19570 54462 19572 54514
rect 19516 54460 19572 54462
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19180 52946 19236 52948
rect 19180 52894 19182 52946
rect 19182 52894 19234 52946
rect 19234 52894 19236 52946
rect 19180 52892 19236 52894
rect 19852 52946 19908 52948
rect 19852 52894 19854 52946
rect 19854 52894 19906 52946
rect 19906 52894 19908 52946
rect 19852 52892 19908 52894
rect 19292 52834 19348 52836
rect 19292 52782 19294 52834
rect 19294 52782 19346 52834
rect 19346 52782 19348 52834
rect 19292 52780 19348 52782
rect 18956 52220 19012 52276
rect 18732 52162 18788 52164
rect 18732 52110 18734 52162
rect 18734 52110 18786 52162
rect 18786 52110 18788 52162
rect 18732 52108 18788 52110
rect 18284 51660 18340 51716
rect 18284 51490 18340 51492
rect 18284 51438 18286 51490
rect 18286 51438 18338 51490
rect 18338 51438 18340 51490
rect 18284 51436 18340 51438
rect 18620 51436 18676 51492
rect 18396 51100 18452 51156
rect 18284 50428 18340 50484
rect 18172 49756 18228 49812
rect 18620 50316 18676 50372
rect 18732 49980 18788 50036
rect 18508 49084 18564 49140
rect 18172 47852 18228 47908
rect 18396 48188 18452 48244
rect 18396 47516 18452 47572
rect 18508 47458 18564 47460
rect 18508 47406 18510 47458
rect 18510 47406 18562 47458
rect 18562 47406 18564 47458
rect 18508 47404 18564 47406
rect 18732 46284 18788 46340
rect 19068 51660 19124 51716
rect 18956 51154 19012 51156
rect 18956 51102 18958 51154
rect 18958 51102 19010 51154
rect 19010 51102 19012 51154
rect 18956 51100 19012 51102
rect 18956 50876 19012 50932
rect 19180 50482 19236 50484
rect 19180 50430 19182 50482
rect 19182 50430 19234 50482
rect 19234 50430 19236 50482
rect 19180 50428 19236 50430
rect 19068 50316 19124 50372
rect 19740 52162 19796 52164
rect 19740 52110 19742 52162
rect 19742 52110 19794 52162
rect 19794 52110 19796 52162
rect 19740 52108 19796 52110
rect 20636 52892 20692 52948
rect 21532 53676 21588 53732
rect 22204 53730 22260 53732
rect 22204 53678 22206 53730
rect 22206 53678 22258 53730
rect 22258 53678 22260 53730
rect 22204 53676 22260 53678
rect 20972 53564 21028 53620
rect 23100 54514 23156 54516
rect 23100 54462 23102 54514
rect 23102 54462 23154 54514
rect 23154 54462 23156 54514
rect 23100 54460 23156 54462
rect 24332 54514 24388 54516
rect 24332 54462 24334 54514
rect 24334 54462 24386 54514
rect 24386 54462 24388 54514
rect 24332 54460 24388 54462
rect 23884 54348 23940 54404
rect 22428 53004 22484 53060
rect 22204 52892 22260 52948
rect 20860 52834 20916 52836
rect 20860 52782 20862 52834
rect 20862 52782 20914 52834
rect 20914 52782 20916 52834
rect 20860 52780 20916 52782
rect 20748 52444 20804 52500
rect 20188 52274 20244 52276
rect 20188 52222 20190 52274
rect 20190 52222 20242 52274
rect 20242 52222 20244 52274
rect 20188 52220 20244 52222
rect 20748 52220 20804 52276
rect 20076 52108 20132 52164
rect 20972 52108 21028 52164
rect 20636 52050 20692 52052
rect 20636 51998 20638 52050
rect 20638 51998 20690 52050
rect 20690 51998 20692 52050
rect 20636 51996 20692 51998
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19628 50988 19684 51044
rect 19404 50764 19460 50820
rect 19404 50428 19460 50484
rect 20076 51266 20132 51268
rect 20076 51214 20078 51266
rect 20078 51214 20130 51266
rect 20130 51214 20132 51266
rect 20076 51212 20132 51214
rect 19852 50876 19908 50932
rect 20188 50988 20244 51044
rect 19740 50428 19796 50484
rect 19964 50482 20020 50484
rect 19964 50430 19966 50482
rect 19966 50430 20018 50482
rect 20018 50430 20020 50482
rect 19964 50428 20020 50430
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19516 49810 19572 49812
rect 19516 49758 19518 49810
rect 19518 49758 19570 49810
rect 19570 49758 19572 49810
rect 19516 49756 19572 49758
rect 19628 49698 19684 49700
rect 19628 49646 19630 49698
rect 19630 49646 19682 49698
rect 19682 49646 19684 49698
rect 19628 49644 19684 49646
rect 19964 49138 20020 49140
rect 19964 49086 19966 49138
rect 19966 49086 20018 49138
rect 20018 49086 20020 49138
rect 19964 49084 20020 49086
rect 19404 48466 19460 48468
rect 19404 48414 19406 48466
rect 19406 48414 19458 48466
rect 19458 48414 19460 48466
rect 19404 48412 19460 48414
rect 19628 48860 19684 48916
rect 20188 48860 20244 48916
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20524 49420 20580 49476
rect 20412 48412 20468 48468
rect 20636 49084 20692 49140
rect 19516 47628 19572 47684
rect 18956 46620 19012 46676
rect 18060 46060 18116 46116
rect 19628 47458 19684 47460
rect 19628 47406 19630 47458
rect 19630 47406 19682 47458
rect 19682 47406 19684 47458
rect 19628 47404 19684 47406
rect 20412 47404 20468 47460
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19740 46898 19796 46900
rect 19740 46846 19742 46898
rect 19742 46846 19794 46898
rect 19794 46846 19796 46898
rect 19740 46844 19796 46846
rect 19068 46060 19124 46116
rect 19292 46620 19348 46676
rect 19292 46060 19348 46116
rect 17948 45052 18004 45108
rect 18284 45778 18340 45780
rect 18284 45726 18286 45778
rect 18286 45726 18338 45778
rect 18338 45726 18340 45778
rect 18284 45724 18340 45726
rect 17948 44882 18004 44884
rect 17948 44830 17950 44882
rect 17950 44830 18002 44882
rect 18002 44830 18004 44882
rect 17948 44828 18004 44830
rect 18172 44380 18228 44436
rect 17948 44322 18004 44324
rect 17948 44270 17950 44322
rect 17950 44270 18002 44322
rect 18002 44270 18004 44322
rect 17948 44268 18004 44270
rect 18060 43484 18116 43540
rect 17052 42866 17108 42868
rect 17052 42814 17054 42866
rect 17054 42814 17106 42866
rect 17106 42814 17108 42866
rect 17052 42812 17108 42814
rect 17164 42642 17220 42644
rect 17164 42590 17166 42642
rect 17166 42590 17218 42642
rect 17218 42590 17220 42642
rect 17164 42588 17220 42590
rect 16940 42252 16996 42308
rect 16940 41970 16996 41972
rect 16940 41918 16942 41970
rect 16942 41918 16994 41970
rect 16994 41918 16996 41970
rect 16940 41916 16996 41918
rect 17724 42754 17780 42756
rect 17724 42702 17726 42754
rect 17726 42702 17778 42754
rect 17778 42702 17780 42754
rect 17724 42700 17780 42702
rect 17500 42588 17556 42644
rect 17388 42140 17444 42196
rect 16268 40908 16324 40964
rect 16828 40684 16884 40740
rect 15484 39618 15540 39620
rect 15484 39566 15486 39618
rect 15486 39566 15538 39618
rect 15538 39566 15540 39618
rect 15484 39564 15540 39566
rect 15372 39228 15428 39284
rect 15260 39116 15316 39172
rect 14140 38780 14196 38836
rect 14028 37436 14084 37492
rect 13804 36652 13860 36708
rect 13804 36370 13860 36372
rect 13804 36318 13806 36370
rect 13806 36318 13858 36370
rect 13858 36318 13860 36370
rect 13804 36316 13860 36318
rect 14028 36482 14084 36484
rect 14028 36430 14030 36482
rect 14030 36430 14082 36482
rect 14082 36430 14084 36482
rect 14028 36428 14084 36430
rect 14028 35308 14084 35364
rect 13580 35084 13636 35140
rect 14364 37436 14420 37492
rect 14364 37266 14420 37268
rect 14364 37214 14366 37266
rect 14366 37214 14418 37266
rect 14418 37214 14420 37266
rect 14364 37212 14420 37214
rect 15372 38946 15428 38948
rect 15372 38894 15374 38946
rect 15374 38894 15426 38946
rect 15426 38894 15428 38946
rect 15372 38892 15428 38894
rect 15148 38780 15204 38836
rect 15708 39116 15764 39172
rect 14700 38220 14756 38276
rect 15596 38332 15652 38388
rect 14812 37938 14868 37940
rect 14812 37886 14814 37938
rect 14814 37886 14866 37938
rect 14866 37886 14868 37938
rect 14812 37884 14868 37886
rect 15036 37324 15092 37380
rect 15372 37378 15428 37380
rect 15372 37326 15374 37378
rect 15374 37326 15426 37378
rect 15426 37326 15428 37378
rect 15372 37324 15428 37326
rect 15036 36988 15092 37044
rect 16044 38892 16100 38948
rect 16492 39564 16548 39620
rect 17052 40572 17108 40628
rect 16492 39116 16548 39172
rect 16268 39058 16324 39060
rect 16268 39006 16270 39058
rect 16270 39006 16322 39058
rect 16322 39006 16324 39058
rect 16268 39004 16324 39006
rect 16380 38668 16436 38724
rect 15708 37100 15764 37156
rect 15820 38050 15876 38052
rect 15820 37998 15822 38050
rect 15822 37998 15874 38050
rect 15874 37998 15876 38050
rect 15820 37996 15876 37998
rect 16044 37660 16100 37716
rect 16492 38556 16548 38612
rect 15820 36988 15876 37044
rect 15932 36876 15988 36932
rect 15820 36652 15876 36708
rect 15260 36482 15316 36484
rect 15260 36430 15262 36482
rect 15262 36430 15314 36482
rect 15314 36430 15316 36482
rect 15260 36428 15316 36430
rect 15036 35196 15092 35252
rect 14140 33740 14196 33796
rect 13356 32620 13412 32676
rect 12460 32562 12516 32564
rect 12460 32510 12462 32562
rect 12462 32510 12514 32562
rect 12514 32510 12516 32562
rect 12460 32508 12516 32510
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 8316 29260 8372 29316
rect 7868 28642 7924 28644
rect 7868 28590 7870 28642
rect 7870 28590 7922 28642
rect 7922 28590 7924 28642
rect 7868 28588 7924 28590
rect 4732 27746 4788 27748
rect 4732 27694 4734 27746
rect 4734 27694 4786 27746
rect 4786 27694 4788 27746
rect 4732 27692 4788 27694
rect 5628 27692 5684 27748
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 5964 27580 6020 27636
rect 7308 27634 7364 27636
rect 7308 27582 7310 27634
rect 7310 27582 7362 27634
rect 7362 27582 7364 27634
rect 7308 27580 7364 27582
rect 6972 27132 7028 27188
rect 7084 26572 7140 26628
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 7420 25676 7476 25732
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 7084 23996 7140 24052
rect 8204 27132 8260 27188
rect 8988 29314 9044 29316
rect 8988 29262 8990 29314
rect 8990 29262 9042 29314
rect 9042 29262 9044 29314
rect 8988 29260 9044 29262
rect 8540 28588 8596 28644
rect 8652 28530 8708 28532
rect 8652 28478 8654 28530
rect 8654 28478 8706 28530
rect 8706 28478 8708 28530
rect 8652 28476 8708 28478
rect 10892 28476 10948 28532
rect 8316 26572 8372 26628
rect 8092 25228 8148 25284
rect 7532 23996 7588 24052
rect 7308 23884 7364 23940
rect 4620 23324 4676 23380
rect 3276 23154 3332 23156
rect 3276 23102 3278 23154
rect 3278 23102 3330 23154
rect 3330 23102 3332 23154
rect 3276 23100 3332 23102
rect 5068 23100 5124 23156
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 2716 22540 2772 22596
rect 4620 21868 4676 21924
rect 6524 23378 6580 23380
rect 6524 23326 6526 23378
rect 6526 23326 6578 23378
rect 6578 23326 6580 23378
rect 6524 23324 6580 23326
rect 6412 23100 6468 23156
rect 5740 22594 5796 22596
rect 5740 22542 5742 22594
rect 5742 22542 5794 22594
rect 5794 22542 5796 22594
rect 5740 22540 5796 22542
rect 6076 22540 6132 22596
rect 6860 22540 6916 22596
rect 4620 21308 4676 21364
rect 6860 22370 6916 22372
rect 6860 22318 6862 22370
rect 6862 22318 6914 22370
rect 6914 22318 6916 22370
rect 6860 22316 6916 22318
rect 6076 21868 6132 21924
rect 6860 21980 6916 22036
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 2716 20690 2772 20692
rect 2716 20638 2718 20690
rect 2718 20638 2770 20690
rect 2770 20638 2772 20690
rect 2716 20636 2772 20638
rect 3836 20690 3892 20692
rect 3836 20638 3838 20690
rect 3838 20638 3890 20690
rect 3890 20638 3892 20690
rect 3836 20636 3892 20638
rect 4732 20690 4788 20692
rect 4732 20638 4734 20690
rect 4734 20638 4786 20690
rect 4786 20638 4788 20690
rect 4732 20636 4788 20638
rect 4956 20412 5012 20468
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 2828 18396 2884 18452
rect 6748 20636 6804 20692
rect 6860 19852 6916 19908
rect 5068 18956 5124 19012
rect 4956 18284 5012 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 3612 17836 3668 17892
rect 5740 19010 5796 19012
rect 5740 18958 5742 19010
rect 5742 18958 5794 19010
rect 5794 18958 5796 19010
rect 5740 18956 5796 18958
rect 6860 18620 6916 18676
rect 5628 18450 5684 18452
rect 5628 18398 5630 18450
rect 5630 18398 5682 18450
rect 5682 18398 5684 18450
rect 5628 18396 5684 18398
rect 5964 18450 6020 18452
rect 5964 18398 5966 18450
rect 5966 18398 6018 18450
rect 6018 18398 6020 18450
rect 5964 18396 6020 18398
rect 5740 17890 5796 17892
rect 5740 17838 5742 17890
rect 5742 17838 5794 17890
rect 5794 17838 5796 17890
rect 5740 17836 5796 17838
rect 6748 18508 6804 18564
rect 6412 17724 6468 17780
rect 2716 16604 2772 16660
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4620 16268 4676 16324
rect 7756 23884 7812 23940
rect 7644 22370 7700 22372
rect 7644 22318 7646 22370
rect 7646 22318 7698 22370
rect 7698 22318 7700 22370
rect 7644 22316 7700 22318
rect 7980 22876 8036 22932
rect 7532 21868 7588 21924
rect 7420 21196 7476 21252
rect 7084 17724 7140 17780
rect 6412 17500 6468 17556
rect 6972 16940 7028 16996
rect 6076 16882 6132 16884
rect 6076 16830 6078 16882
rect 6078 16830 6130 16882
rect 6130 16830 6132 16882
rect 6076 16828 6132 16830
rect 5964 16716 6020 16772
rect 5740 16604 5796 16660
rect 6076 16322 6132 16324
rect 6076 16270 6078 16322
rect 6078 16270 6130 16322
rect 6130 16270 6132 16322
rect 6076 16268 6132 16270
rect 2380 15260 2436 15316
rect 2940 15314 2996 15316
rect 2940 15262 2942 15314
rect 2942 15262 2994 15314
rect 2994 15262 2996 15314
rect 2940 15260 2996 15262
rect 5068 15260 5124 15316
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5068 14476 5124 14532
rect 5964 14530 6020 14532
rect 5964 14478 5966 14530
rect 5966 14478 6018 14530
rect 6018 14478 6020 14530
rect 5964 14476 6020 14478
rect 4172 14418 4228 14420
rect 4172 14366 4174 14418
rect 4174 14366 4226 14418
rect 4226 14366 4228 14418
rect 4172 14364 4228 14366
rect 6188 14364 6244 14420
rect 2492 13804 2548 13860
rect 3724 13858 3780 13860
rect 3724 13806 3726 13858
rect 3726 13806 3778 13858
rect 3778 13806 3780 13858
rect 3724 13804 3780 13806
rect 3276 13132 3332 13188
rect 5292 13634 5348 13636
rect 5292 13582 5294 13634
rect 5294 13582 5346 13634
rect 5346 13582 5348 13634
rect 5292 13580 5348 13582
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5740 13186 5796 13188
rect 5740 13134 5742 13186
rect 5742 13134 5794 13186
rect 5794 13134 5796 13186
rect 5740 13132 5796 13134
rect 6412 13020 6468 13076
rect 4956 12908 5012 12964
rect 6076 12962 6132 12964
rect 6076 12910 6078 12962
rect 6078 12910 6130 12962
rect 6130 12910 6132 12962
rect 6076 12908 6132 12910
rect 6860 15932 6916 15988
rect 6972 15314 7028 15316
rect 6972 15262 6974 15314
rect 6974 15262 7026 15314
rect 7026 15262 7028 15314
rect 6972 15260 7028 15262
rect 7308 19068 7364 19124
rect 7644 21308 7700 21364
rect 7868 21474 7924 21476
rect 7868 21422 7870 21474
rect 7870 21422 7922 21474
rect 7922 21422 7924 21474
rect 7868 21420 7924 21422
rect 8876 25564 8932 25620
rect 8652 24050 8708 24052
rect 8652 23998 8654 24050
rect 8654 23998 8706 24050
rect 8706 23998 8708 24050
rect 8652 23996 8708 23998
rect 9212 24050 9268 24052
rect 9212 23998 9214 24050
rect 9214 23998 9266 24050
rect 9266 23998 9268 24050
rect 9212 23996 9268 23998
rect 8988 22764 9044 22820
rect 8652 22594 8708 22596
rect 8652 22542 8654 22594
rect 8654 22542 8706 22594
rect 8706 22542 8708 22594
rect 8652 22540 8708 22542
rect 8764 21756 8820 21812
rect 8876 21644 8932 21700
rect 8540 21586 8596 21588
rect 8540 21534 8542 21586
rect 8542 21534 8594 21586
rect 8594 21534 8596 21586
rect 8540 21532 8596 21534
rect 7980 21026 8036 21028
rect 7980 20974 7982 21026
rect 7982 20974 8034 21026
rect 8034 20974 8036 21026
rect 7980 20972 8036 20974
rect 7756 20412 7812 20468
rect 7644 19906 7700 19908
rect 7644 19854 7646 19906
rect 7646 19854 7698 19906
rect 7698 19854 7700 19906
rect 7644 19852 7700 19854
rect 7532 19740 7588 19796
rect 7980 19740 8036 19796
rect 8092 18956 8148 19012
rect 8652 21474 8708 21476
rect 8652 21422 8654 21474
rect 8654 21422 8706 21474
rect 8706 21422 8708 21474
rect 8652 21420 8708 21422
rect 8540 21026 8596 21028
rect 8540 20974 8542 21026
rect 8542 20974 8594 21026
rect 8594 20974 8596 21026
rect 8540 20972 8596 20974
rect 8204 19292 8260 19348
rect 8540 20802 8596 20804
rect 8540 20750 8542 20802
rect 8542 20750 8594 20802
rect 8594 20750 8596 20802
rect 8540 20748 8596 20750
rect 8316 19122 8372 19124
rect 8316 19070 8318 19122
rect 8318 19070 8370 19122
rect 8370 19070 8372 19122
rect 8316 19068 8372 19070
rect 7980 18508 8036 18564
rect 8988 20972 9044 21028
rect 8876 20860 8932 20916
rect 8988 19964 9044 20020
rect 8652 19068 8708 19124
rect 7868 17554 7924 17556
rect 7868 17502 7870 17554
rect 7870 17502 7922 17554
rect 7922 17502 7924 17554
rect 7868 17500 7924 17502
rect 8092 17554 8148 17556
rect 8092 17502 8094 17554
rect 8094 17502 8146 17554
rect 8146 17502 8148 17554
rect 8092 17500 8148 17502
rect 8876 18396 8932 18452
rect 9324 22764 9380 22820
rect 10220 27020 10276 27076
rect 10780 27074 10836 27076
rect 10780 27022 10782 27074
rect 10782 27022 10834 27074
rect 10834 27022 10836 27074
rect 10780 27020 10836 27022
rect 10108 26572 10164 26628
rect 11116 27186 11172 27188
rect 11116 27134 11118 27186
rect 11118 27134 11170 27186
rect 11170 27134 11172 27186
rect 11116 27132 11172 27134
rect 13580 32508 13636 32564
rect 13132 31836 13188 31892
rect 13916 31890 13972 31892
rect 13916 31838 13918 31890
rect 13918 31838 13970 31890
rect 13970 31838 13972 31890
rect 13916 31836 13972 31838
rect 13804 31778 13860 31780
rect 13804 31726 13806 31778
rect 13806 31726 13858 31778
rect 13858 31726 13860 31778
rect 13804 31724 13860 31726
rect 13468 31612 13524 31668
rect 13244 31218 13300 31220
rect 13244 31166 13246 31218
rect 13246 31166 13298 31218
rect 13298 31166 13300 31218
rect 13244 31164 13300 31166
rect 14140 31164 14196 31220
rect 12236 29426 12292 29428
rect 12236 29374 12238 29426
rect 12238 29374 12290 29426
rect 12290 29374 12292 29426
rect 12236 29372 12292 29374
rect 13468 29372 13524 29428
rect 12908 28588 12964 28644
rect 13468 28642 13524 28644
rect 13468 28590 13470 28642
rect 13470 28590 13522 28642
rect 13522 28590 13524 28642
rect 13468 28588 13524 28590
rect 13804 28588 13860 28644
rect 11116 26460 11172 26516
rect 9660 26236 9716 26292
rect 9884 25618 9940 25620
rect 9884 25566 9886 25618
rect 9886 25566 9938 25618
rect 9938 25566 9940 25618
rect 9884 25564 9940 25566
rect 10332 25282 10388 25284
rect 10332 25230 10334 25282
rect 10334 25230 10386 25282
rect 10386 25230 10388 25282
rect 10332 25228 10388 25230
rect 10668 25340 10724 25396
rect 11452 25676 11508 25732
rect 11228 25564 11284 25620
rect 11452 25228 11508 25284
rect 11564 25340 11620 25396
rect 9660 23154 9716 23156
rect 9660 23102 9662 23154
rect 9662 23102 9714 23154
rect 9714 23102 9716 23154
rect 9660 23100 9716 23102
rect 9884 21756 9940 21812
rect 9772 21586 9828 21588
rect 9772 21534 9774 21586
rect 9774 21534 9826 21586
rect 9826 21534 9828 21586
rect 9772 21532 9828 21534
rect 11900 25394 11956 25396
rect 11900 25342 11902 25394
rect 11902 25342 11954 25394
rect 11954 25342 11956 25394
rect 11900 25340 11956 25342
rect 10108 21644 10164 21700
rect 11228 21698 11284 21700
rect 11228 21646 11230 21698
rect 11230 21646 11282 21698
rect 11282 21646 11284 21698
rect 11228 21644 11284 21646
rect 11900 21698 11956 21700
rect 11900 21646 11902 21698
rect 11902 21646 11954 21698
rect 11954 21646 11956 21698
rect 11900 21644 11956 21646
rect 9660 21474 9716 21476
rect 9660 21422 9662 21474
rect 9662 21422 9714 21474
rect 9714 21422 9716 21474
rect 9660 21420 9716 21422
rect 11564 21308 11620 21364
rect 9548 19906 9604 19908
rect 9548 19854 9550 19906
rect 9550 19854 9602 19906
rect 9602 19854 9604 19906
rect 9548 19852 9604 19854
rect 11564 19794 11620 19796
rect 11564 19742 11566 19794
rect 11566 19742 11618 19794
rect 11618 19742 11620 19794
rect 11564 19740 11620 19742
rect 10108 19010 10164 19012
rect 10108 18958 10110 19010
rect 10110 18958 10162 19010
rect 10162 18958 10164 19010
rect 10108 18956 10164 18958
rect 9548 18620 9604 18676
rect 9100 18396 9156 18452
rect 9436 18508 9492 18564
rect 8988 17554 9044 17556
rect 8988 17502 8990 17554
rect 8990 17502 9042 17554
rect 9042 17502 9044 17554
rect 8988 17500 9044 17502
rect 9212 17500 9268 17556
rect 8316 17442 8372 17444
rect 8316 17390 8318 17442
rect 8318 17390 8370 17442
rect 8370 17390 8372 17442
rect 8316 17388 8372 17390
rect 9212 17276 9268 17332
rect 7308 16828 7364 16884
rect 7644 16828 7700 16884
rect 7420 16770 7476 16772
rect 7420 16718 7422 16770
rect 7422 16718 7474 16770
rect 7474 16718 7476 16770
rect 7420 16716 7476 16718
rect 7868 16940 7924 16996
rect 9324 16492 9380 16548
rect 7420 15986 7476 15988
rect 7420 15934 7422 15986
rect 7422 15934 7474 15986
rect 7474 15934 7476 15986
rect 7420 15932 7476 15934
rect 7756 15986 7812 15988
rect 7756 15934 7758 15986
rect 7758 15934 7810 15986
rect 7810 15934 7812 15986
rect 7756 15932 7812 15934
rect 7644 15484 7700 15540
rect 7084 14530 7140 14532
rect 7084 14478 7086 14530
rect 7086 14478 7138 14530
rect 7138 14478 7140 14530
rect 7084 14476 7140 14478
rect 4060 12348 4116 12404
rect 4620 12572 4676 12628
rect 5404 12572 5460 12628
rect 5068 12402 5124 12404
rect 5068 12350 5070 12402
rect 5070 12350 5122 12402
rect 5122 12350 5124 12402
rect 5068 12348 5124 12350
rect 6076 12290 6132 12292
rect 6076 12238 6078 12290
rect 6078 12238 6130 12290
rect 6130 12238 6132 12290
rect 6076 12236 6132 12238
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 8204 14476 8260 14532
rect 8316 15820 8372 15876
rect 8540 15260 8596 15316
rect 8204 13580 8260 13636
rect 8988 14364 9044 14420
rect 9100 13970 9156 13972
rect 9100 13918 9102 13970
rect 9102 13918 9154 13970
rect 9154 13918 9156 13970
rect 9100 13916 9156 13918
rect 8540 13356 8596 13412
rect 7196 12236 7252 12292
rect 8204 13244 8260 13300
rect 7420 11564 7476 11620
rect 1820 11452 1876 11508
rect 4844 11506 4900 11508
rect 4844 11454 4846 11506
rect 4846 11454 4898 11506
rect 4898 11454 4900 11506
rect 4844 11452 4900 11454
rect 5628 11452 5684 11508
rect 6076 11452 6132 11508
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 8876 13580 8932 13636
rect 6636 9660 6692 9716
rect 7308 9714 7364 9716
rect 7308 9662 7310 9714
rect 7310 9662 7362 9714
rect 7362 9662 7364 9714
rect 7308 9660 7364 9662
rect 8316 12236 8372 12292
rect 8540 11564 8596 11620
rect 9660 18172 9716 18228
rect 9996 18450 10052 18452
rect 9996 18398 9998 18450
rect 9998 18398 10050 18450
rect 10050 18398 10052 18450
rect 9996 18396 10052 18398
rect 10220 18396 10276 18452
rect 9548 17724 9604 17780
rect 10444 18060 10500 18116
rect 10668 17554 10724 17556
rect 10668 17502 10670 17554
rect 10670 17502 10722 17554
rect 10722 17502 10724 17554
rect 10668 17500 10724 17502
rect 9772 16492 9828 16548
rect 10332 16828 10388 16884
rect 10332 15260 10388 15316
rect 10444 15932 10500 15988
rect 10892 15932 10948 15988
rect 11116 18396 11172 18452
rect 11116 17948 11172 18004
rect 11452 18396 11508 18452
rect 15372 34972 15428 35028
rect 16156 36652 16212 36708
rect 16604 38220 16660 38276
rect 17052 39506 17108 39508
rect 17052 39454 17054 39506
rect 17054 39454 17106 39506
rect 17106 39454 17108 39506
rect 17052 39452 17108 39454
rect 17724 42476 17780 42532
rect 17164 38556 17220 38612
rect 17612 40236 17668 40292
rect 17948 42812 18004 42868
rect 18284 44322 18340 44324
rect 18284 44270 18286 44322
rect 18286 44270 18338 44322
rect 18338 44270 18340 44322
rect 18284 44268 18340 44270
rect 18844 45164 18900 45220
rect 19516 46284 19572 46340
rect 18620 44940 18676 44996
rect 18956 44268 19012 44324
rect 19068 45052 19124 45108
rect 19068 44716 19124 44772
rect 18284 43820 18340 43876
rect 18844 44044 18900 44100
rect 18060 42364 18116 42420
rect 17948 42028 18004 42084
rect 18172 41970 18228 41972
rect 18172 41918 18174 41970
rect 18174 41918 18226 41970
rect 18226 41918 18228 41970
rect 18172 41916 18228 41918
rect 18396 43596 18452 43652
rect 18620 43314 18676 43316
rect 18620 43262 18622 43314
rect 18622 43262 18674 43314
rect 18674 43262 18676 43314
rect 18620 43260 18676 43262
rect 18508 42642 18564 42644
rect 18508 42590 18510 42642
rect 18510 42590 18562 42642
rect 18562 42590 18564 42642
rect 18508 42588 18564 42590
rect 19404 45500 19460 45556
rect 19292 44828 19348 44884
rect 19292 43932 19348 43988
rect 19404 43820 19460 43876
rect 19292 43762 19348 43764
rect 19292 43710 19294 43762
rect 19294 43710 19346 43762
rect 19346 43710 19348 43762
rect 19292 43708 19348 43710
rect 20748 48188 20804 48244
rect 22764 51996 22820 52052
rect 22316 51602 22372 51604
rect 22316 51550 22318 51602
rect 22318 51550 22370 51602
rect 22370 51550 22372 51602
rect 22316 51548 22372 51550
rect 22092 51266 22148 51268
rect 22092 51214 22094 51266
rect 22094 51214 22146 51266
rect 22146 51214 22148 51266
rect 22092 51212 22148 51214
rect 21980 50540 22036 50596
rect 22092 49868 22148 49924
rect 21196 49586 21252 49588
rect 21196 49534 21198 49586
rect 21198 49534 21250 49586
rect 21250 49534 21252 49586
rect 21196 49532 21252 49534
rect 21084 49420 21140 49476
rect 20972 48972 21028 49028
rect 21868 49586 21924 49588
rect 21868 49534 21870 49586
rect 21870 49534 21922 49586
rect 21922 49534 21924 49586
rect 21868 49532 21924 49534
rect 22428 49756 22484 49812
rect 21420 49084 21476 49140
rect 25116 54908 25172 54964
rect 24668 54348 24724 54404
rect 22988 52108 23044 52164
rect 23100 51996 23156 52052
rect 22876 51660 22932 51716
rect 23100 51490 23156 51492
rect 23100 51438 23102 51490
rect 23102 51438 23154 51490
rect 23154 51438 23156 51490
rect 23100 51436 23156 51438
rect 22876 50482 22932 50484
rect 22876 50430 22878 50482
rect 22878 50430 22930 50482
rect 22930 50430 22932 50482
rect 22876 50428 22932 50430
rect 23548 53618 23604 53620
rect 23548 53566 23550 53618
rect 23550 53566 23602 53618
rect 23602 53566 23604 53618
rect 23548 53564 23604 53566
rect 23772 53116 23828 53172
rect 24220 53116 24276 53172
rect 23548 52946 23604 52948
rect 23548 52894 23550 52946
rect 23550 52894 23602 52946
rect 23602 52894 23604 52946
rect 23548 52892 23604 52894
rect 23996 52946 24052 52948
rect 23996 52894 23998 52946
rect 23998 52894 24050 52946
rect 24050 52894 24052 52946
rect 23996 52892 24052 52894
rect 24556 53004 24612 53060
rect 25004 53004 25060 53060
rect 23548 52162 23604 52164
rect 23548 52110 23550 52162
rect 23550 52110 23602 52162
rect 23602 52110 23604 52162
rect 23548 52108 23604 52110
rect 23660 51602 23716 51604
rect 23660 51550 23662 51602
rect 23662 51550 23714 51602
rect 23714 51550 23716 51602
rect 23660 51548 23716 51550
rect 23436 50764 23492 50820
rect 22876 49868 22932 49924
rect 23100 49810 23156 49812
rect 23100 49758 23102 49810
rect 23102 49758 23154 49810
rect 23154 49758 23156 49810
rect 23100 49756 23156 49758
rect 22988 49698 23044 49700
rect 22988 49646 22990 49698
rect 22990 49646 23042 49698
rect 23042 49646 23044 49698
rect 22988 49644 23044 49646
rect 22988 49196 23044 49252
rect 21308 48860 21364 48916
rect 20748 47068 20804 47124
rect 20748 46898 20804 46900
rect 20748 46846 20750 46898
rect 20750 46846 20802 46898
rect 20802 46846 20804 46898
rect 20748 46844 20804 46846
rect 20860 46620 20916 46676
rect 20300 45778 20356 45780
rect 20300 45726 20302 45778
rect 20302 45726 20354 45778
rect 20354 45726 20356 45778
rect 20300 45724 20356 45726
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 20300 44994 20356 44996
rect 20300 44942 20302 44994
rect 20302 44942 20354 44994
rect 20354 44942 20356 44994
rect 20300 44940 20356 44942
rect 19852 44604 19908 44660
rect 20076 44268 20132 44324
rect 19740 44044 19796 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19964 43596 20020 43652
rect 19180 42364 19236 42420
rect 18844 42252 18900 42308
rect 18508 42082 18564 42084
rect 18508 42030 18510 42082
rect 18510 42030 18562 42082
rect 18562 42030 18564 42082
rect 18508 42028 18564 42030
rect 17948 41186 18004 41188
rect 17948 41134 17950 41186
rect 17950 41134 18002 41186
rect 18002 41134 18004 41186
rect 17948 41132 18004 41134
rect 18956 41916 19012 41972
rect 17724 39788 17780 39844
rect 17836 40012 17892 40068
rect 17500 39452 17556 39508
rect 17724 39004 17780 39060
rect 17500 38780 17556 38836
rect 17276 38332 17332 38388
rect 17388 38444 17444 38500
rect 15820 35868 15876 35924
rect 15932 36316 15988 36372
rect 15932 35756 15988 35812
rect 16492 36316 16548 36372
rect 16044 35698 16100 35700
rect 16044 35646 16046 35698
rect 16046 35646 16098 35698
rect 16098 35646 16100 35698
rect 16044 35644 16100 35646
rect 14812 33906 14868 33908
rect 14812 33854 14814 33906
rect 14814 33854 14866 33906
rect 14866 33854 14868 33906
rect 14812 33852 14868 33854
rect 16716 36540 16772 36596
rect 17388 37772 17444 37828
rect 17948 39004 18004 39060
rect 17836 38556 17892 38612
rect 17612 38162 17668 38164
rect 17612 38110 17614 38162
rect 17614 38110 17666 38162
rect 17666 38110 17668 38162
rect 17612 38108 17668 38110
rect 17836 37378 17892 37380
rect 17836 37326 17838 37378
rect 17838 37326 17890 37378
rect 17890 37326 17892 37378
rect 17836 37324 17892 37326
rect 17836 36988 17892 37044
rect 16716 35644 16772 35700
rect 16604 35420 16660 35476
rect 17388 35922 17444 35924
rect 17388 35870 17390 35922
rect 17390 35870 17442 35922
rect 17442 35870 17444 35922
rect 17388 35868 17444 35870
rect 17164 35196 17220 35252
rect 17276 35308 17332 35364
rect 15820 33180 15876 33236
rect 16380 33180 16436 33236
rect 15708 32508 15764 32564
rect 14812 31890 14868 31892
rect 14812 31838 14814 31890
rect 14814 31838 14866 31890
rect 14866 31838 14868 31890
rect 14812 31836 14868 31838
rect 15596 31890 15652 31892
rect 15596 31838 15598 31890
rect 15598 31838 15650 31890
rect 15650 31838 15652 31890
rect 15596 31836 15652 31838
rect 17724 34076 17780 34132
rect 18284 40572 18340 40628
rect 18508 40290 18564 40292
rect 18508 40238 18510 40290
rect 18510 40238 18562 40290
rect 18562 40238 18564 40290
rect 18508 40236 18564 40238
rect 18284 40178 18340 40180
rect 18284 40126 18286 40178
rect 18286 40126 18338 40178
rect 18338 40126 18340 40178
rect 18284 40124 18340 40126
rect 18284 39788 18340 39844
rect 18732 40572 18788 40628
rect 18620 39564 18676 39620
rect 19404 43484 19460 43540
rect 19852 42754 19908 42756
rect 19852 42702 19854 42754
rect 19854 42702 19906 42754
rect 19906 42702 19908 42754
rect 19852 42700 19908 42702
rect 19404 42476 19460 42532
rect 19292 42252 19348 42308
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19292 42082 19348 42084
rect 19292 42030 19294 42082
rect 19294 42030 19346 42082
rect 19346 42030 19348 42082
rect 19292 42028 19348 42030
rect 19068 40962 19124 40964
rect 19068 40910 19070 40962
rect 19070 40910 19122 40962
rect 19122 40910 19124 40962
rect 19068 40908 19124 40910
rect 19404 40572 19460 40628
rect 20188 42028 20244 42084
rect 19964 41858 20020 41860
rect 19964 41806 19966 41858
rect 19966 41806 20018 41858
rect 20018 41806 20020 41858
rect 19964 41804 20020 41806
rect 19964 41580 20020 41636
rect 20300 41970 20356 41972
rect 20300 41918 20302 41970
rect 20302 41918 20354 41970
rect 20354 41918 20356 41970
rect 20300 41916 20356 41918
rect 19516 40460 19572 40516
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 18620 39116 18676 39172
rect 18284 38722 18340 38724
rect 18284 38670 18286 38722
rect 18286 38670 18338 38722
rect 18338 38670 18340 38722
rect 18284 38668 18340 38670
rect 18508 38108 18564 38164
rect 17948 35868 18004 35924
rect 18396 37100 18452 37156
rect 19740 40572 19796 40628
rect 19180 40178 19236 40180
rect 19180 40126 19182 40178
rect 19182 40126 19234 40178
rect 19234 40126 19236 40178
rect 19180 40124 19236 40126
rect 19292 40012 19348 40068
rect 19292 39116 19348 39172
rect 20636 45948 20692 46004
rect 20524 44268 20580 44324
rect 20636 44044 20692 44100
rect 20636 43484 20692 43540
rect 20860 43372 20916 43428
rect 20524 43148 20580 43204
rect 20524 41804 20580 41860
rect 20188 40236 20244 40292
rect 20748 41746 20804 41748
rect 20748 41694 20750 41746
rect 20750 41694 20802 41746
rect 20802 41694 20804 41746
rect 20748 41692 20804 41694
rect 21420 48130 21476 48132
rect 21420 48078 21422 48130
rect 21422 48078 21474 48130
rect 21474 48078 21476 48130
rect 21420 48076 21476 48078
rect 21308 47458 21364 47460
rect 21308 47406 21310 47458
rect 21310 47406 21362 47458
rect 21362 47406 21364 47458
rect 21308 47404 21364 47406
rect 21196 47068 21252 47124
rect 21756 47404 21812 47460
rect 21532 47068 21588 47124
rect 21196 43708 21252 43764
rect 20636 40236 20692 40292
rect 21084 42140 21140 42196
rect 19964 39452 20020 39508
rect 20524 39452 20580 39508
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19740 39004 19796 39060
rect 20524 38892 20580 38948
rect 20300 38834 20356 38836
rect 20300 38782 20302 38834
rect 20302 38782 20354 38834
rect 20354 38782 20356 38834
rect 20300 38780 20356 38782
rect 19964 38444 20020 38500
rect 18732 37660 18788 37716
rect 18732 37212 18788 37268
rect 19068 37266 19124 37268
rect 19068 37214 19070 37266
rect 19070 37214 19122 37266
rect 19122 37214 19124 37266
rect 19068 37212 19124 37214
rect 18732 36988 18788 37044
rect 19628 37826 19684 37828
rect 19628 37774 19630 37826
rect 19630 37774 19682 37826
rect 19682 37774 19684 37826
rect 19628 37772 19684 37774
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20076 37436 20132 37492
rect 20300 37324 20356 37380
rect 19628 37100 19684 37156
rect 19852 37154 19908 37156
rect 19852 37102 19854 37154
rect 19854 37102 19906 37154
rect 19906 37102 19908 37154
rect 19852 37100 19908 37102
rect 19404 36988 19460 37044
rect 19180 36764 19236 36820
rect 19292 36876 19348 36932
rect 18620 35922 18676 35924
rect 18620 35870 18622 35922
rect 18622 35870 18674 35922
rect 18674 35870 18676 35922
rect 18620 35868 18676 35870
rect 18508 35084 18564 35140
rect 18620 35420 18676 35476
rect 18956 36204 19012 36260
rect 19068 35810 19124 35812
rect 19068 35758 19070 35810
rect 19070 35758 19122 35810
rect 19122 35758 19124 35810
rect 19068 35756 19124 35758
rect 20188 36988 20244 37044
rect 19516 36258 19572 36260
rect 19516 36206 19518 36258
rect 19518 36206 19570 36258
rect 19570 36206 19572 36258
rect 19516 36204 19572 36206
rect 19836 36090 19892 36092
rect 19516 35980 19572 36036
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 18956 35138 19012 35140
rect 18956 35086 18958 35138
rect 18958 35086 19010 35138
rect 19010 35086 19012 35138
rect 18956 35084 19012 35086
rect 18732 35026 18788 35028
rect 18732 34974 18734 35026
rect 18734 34974 18786 35026
rect 18786 34974 18788 35026
rect 18732 34972 18788 34974
rect 18844 34860 18900 34916
rect 17948 33964 18004 34020
rect 18620 34076 18676 34132
rect 17612 33852 17668 33908
rect 16828 33234 16884 33236
rect 16828 33182 16830 33234
rect 16830 33182 16882 33234
rect 16882 33182 16884 33234
rect 16828 33180 16884 33182
rect 15932 31724 15988 31780
rect 15596 31554 15652 31556
rect 15596 31502 15598 31554
rect 15598 31502 15650 31554
rect 15650 31502 15652 31554
rect 15596 31500 15652 31502
rect 15932 31388 15988 31444
rect 14588 31164 14644 31220
rect 16492 31500 16548 31556
rect 16380 30828 16436 30884
rect 16156 30716 16212 30772
rect 16492 30716 16548 30772
rect 15708 30098 15764 30100
rect 15708 30046 15710 30098
rect 15710 30046 15762 30098
rect 15762 30046 15764 30098
rect 15708 30044 15764 30046
rect 16044 29986 16100 29988
rect 16044 29934 16046 29986
rect 16046 29934 16098 29986
rect 16098 29934 16100 29986
rect 16044 29932 16100 29934
rect 17388 30882 17444 30884
rect 17388 30830 17390 30882
rect 17390 30830 17442 30882
rect 17442 30830 17444 30882
rect 17388 30828 17444 30830
rect 17948 33122 18004 33124
rect 17948 33070 17950 33122
rect 17950 33070 18002 33122
rect 18002 33070 18004 33122
rect 17948 33068 18004 33070
rect 17836 31724 17892 31780
rect 17724 31388 17780 31444
rect 17836 31164 17892 31220
rect 17948 30828 18004 30884
rect 16604 30098 16660 30100
rect 16604 30046 16606 30098
rect 16606 30046 16658 30098
rect 16658 30046 16660 30098
rect 16604 30044 16660 30046
rect 16156 29820 16212 29876
rect 15932 29484 15988 29540
rect 12348 26290 12404 26292
rect 12348 26238 12350 26290
rect 12350 26238 12402 26290
rect 12402 26238 12404 26290
rect 12348 26236 12404 26238
rect 12236 25676 12292 25732
rect 12796 25676 12852 25732
rect 12124 25340 12180 25396
rect 12908 25340 12964 25396
rect 13916 26460 13972 26516
rect 13916 25564 13972 25620
rect 14140 25394 14196 25396
rect 14140 25342 14142 25394
rect 14142 25342 14194 25394
rect 14194 25342 14196 25394
rect 14140 25340 14196 25342
rect 14700 25394 14756 25396
rect 14700 25342 14702 25394
rect 14702 25342 14754 25394
rect 14754 25342 14756 25394
rect 14700 25340 14756 25342
rect 15260 25340 15316 25396
rect 15484 29314 15540 29316
rect 15484 29262 15486 29314
rect 15486 29262 15538 29314
rect 15538 29262 15540 29314
rect 15484 29260 15540 29262
rect 16828 29260 16884 29316
rect 15484 28588 15540 28644
rect 17388 29932 17444 29988
rect 17948 29820 18004 29876
rect 18284 33068 18340 33124
rect 18396 31724 18452 31780
rect 18396 31388 18452 31444
rect 18284 30882 18340 30884
rect 18284 30830 18286 30882
rect 18286 30830 18338 30882
rect 18338 30830 18340 30882
rect 18284 30828 18340 30830
rect 18732 33628 18788 33684
rect 20300 36092 20356 36148
rect 20188 35868 20244 35924
rect 19628 35196 19684 35252
rect 18956 34188 19012 34244
rect 19068 34076 19124 34132
rect 18956 33740 19012 33796
rect 19292 33740 19348 33796
rect 19404 33628 19460 33684
rect 18732 31666 18788 31668
rect 18732 31614 18734 31666
rect 18734 31614 18786 31666
rect 18786 31614 18788 31666
rect 18732 31612 18788 31614
rect 18732 31164 18788 31220
rect 19068 30882 19124 30884
rect 19068 30830 19070 30882
rect 19070 30830 19122 30882
rect 19122 30830 19124 30882
rect 19068 30828 19124 30830
rect 18732 30770 18788 30772
rect 18732 30718 18734 30770
rect 18734 30718 18786 30770
rect 18786 30718 18788 30770
rect 18732 30716 18788 30718
rect 18060 29708 18116 29764
rect 18396 30156 18452 30212
rect 18060 29538 18116 29540
rect 18060 29486 18062 29538
rect 18062 29486 18114 29538
rect 18114 29486 18116 29538
rect 18060 29484 18116 29486
rect 17164 29036 17220 29092
rect 17836 29036 17892 29092
rect 16828 28028 16884 28084
rect 17500 28082 17556 28084
rect 17500 28030 17502 28082
rect 17502 28030 17554 28082
rect 17554 28030 17556 28082
rect 17500 28028 17556 28030
rect 17164 27580 17220 27636
rect 15484 25564 15540 25620
rect 16156 25116 16212 25172
rect 16268 24892 16324 24948
rect 15820 24722 15876 24724
rect 15820 24670 15822 24722
rect 15822 24670 15874 24722
rect 15874 24670 15876 24722
rect 15820 24668 15876 24670
rect 16268 24722 16324 24724
rect 16268 24670 16270 24722
rect 16270 24670 16322 24722
rect 16322 24670 16324 24722
rect 16268 24668 16324 24670
rect 12348 23212 12404 23268
rect 13692 23436 13748 23492
rect 12572 23042 12628 23044
rect 12572 22990 12574 23042
rect 12574 22990 12626 23042
rect 12626 22990 12628 23042
rect 12572 22988 12628 22990
rect 12236 21586 12292 21588
rect 12236 21534 12238 21586
rect 12238 21534 12290 21586
rect 12290 21534 12292 21586
rect 12236 21532 12292 21534
rect 12348 21420 12404 21476
rect 12348 20636 12404 20692
rect 13916 23212 13972 23268
rect 13804 22988 13860 23044
rect 13468 22876 13524 22932
rect 12908 22204 12964 22260
rect 12572 21532 12628 21588
rect 13468 22204 13524 22260
rect 13804 22540 13860 22596
rect 12796 21196 12852 21252
rect 12908 20802 12964 20804
rect 12908 20750 12910 20802
rect 12910 20750 12962 20802
rect 12962 20750 12964 20802
rect 12908 20748 12964 20750
rect 13580 20748 13636 20804
rect 12572 20636 12628 20692
rect 11900 17836 11956 17892
rect 11116 16828 11172 16884
rect 12684 20524 12740 20580
rect 12796 19404 12852 19460
rect 12460 18396 12516 18452
rect 12572 17890 12628 17892
rect 12572 17838 12574 17890
rect 12574 17838 12626 17890
rect 12626 17838 12628 17890
rect 12572 17836 12628 17838
rect 11676 16268 11732 16324
rect 11564 15874 11620 15876
rect 11564 15822 11566 15874
rect 11566 15822 11618 15874
rect 11618 15822 11620 15874
rect 11564 15820 11620 15822
rect 9884 14642 9940 14644
rect 9884 14590 9886 14642
rect 9886 14590 9938 14642
rect 9938 14590 9940 14642
rect 9884 14588 9940 14590
rect 10892 14642 10948 14644
rect 10892 14590 10894 14642
rect 10894 14590 10946 14642
rect 10946 14590 10948 14642
rect 10892 14588 10948 14590
rect 10220 14418 10276 14420
rect 10220 14366 10222 14418
rect 10222 14366 10274 14418
rect 10274 14366 10276 14418
rect 10220 14364 10276 14366
rect 11228 14252 11284 14308
rect 10668 13634 10724 13636
rect 10668 13582 10670 13634
rect 10670 13582 10722 13634
rect 10722 13582 10724 13634
rect 10668 13580 10724 13582
rect 9996 13356 10052 13412
rect 9772 13244 9828 13300
rect 12796 18450 12852 18452
rect 12796 18398 12798 18450
rect 12798 18398 12850 18450
rect 12850 18398 12852 18450
rect 12796 18396 12852 18398
rect 13356 18508 13412 18564
rect 12908 18284 12964 18340
rect 12908 17724 12964 17780
rect 12460 16828 12516 16884
rect 12124 16268 12180 16324
rect 12012 15426 12068 15428
rect 12012 15374 12014 15426
rect 12014 15374 12066 15426
rect 12066 15374 12068 15426
rect 12012 15372 12068 15374
rect 12460 15986 12516 15988
rect 12460 15934 12462 15986
rect 12462 15934 12514 15986
rect 12514 15934 12516 15986
rect 12460 15932 12516 15934
rect 13020 16882 13076 16884
rect 13020 16830 13022 16882
rect 13022 16830 13074 16882
rect 13074 16830 13076 16882
rect 13020 16828 13076 16830
rect 12908 16604 12964 16660
rect 11900 14588 11956 14644
rect 11788 13916 11844 13972
rect 11228 13020 11284 13076
rect 11340 13468 11396 13524
rect 8876 11452 8932 11508
rect 9548 11452 9604 11508
rect 8540 11228 8596 11284
rect 8988 9660 9044 9716
rect 7644 8876 7700 8932
rect 8988 8930 9044 8932
rect 8988 8878 8990 8930
rect 8990 8878 9042 8930
rect 9042 8878 9044 8930
rect 8988 8876 9044 8878
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 10892 12684 10948 12740
rect 10220 12178 10276 12180
rect 10220 12126 10222 12178
rect 10222 12126 10274 12178
rect 10274 12126 10276 12178
rect 10220 12124 10276 12126
rect 11676 13132 11732 13188
rect 12012 12908 12068 12964
rect 12236 13804 12292 13860
rect 11340 12572 11396 12628
rect 9772 8316 9828 8372
rect 11900 9714 11956 9716
rect 11900 9662 11902 9714
rect 11902 9662 11954 9714
rect 11954 9662 11956 9714
rect 11900 9660 11956 9662
rect 12460 13356 12516 13412
rect 12572 13132 12628 13188
rect 12348 12178 12404 12180
rect 12348 12126 12350 12178
rect 12350 12126 12402 12178
rect 12402 12126 12404 12178
rect 12348 12124 12404 12126
rect 12796 15538 12852 15540
rect 12796 15486 12798 15538
rect 12798 15486 12850 15538
rect 12850 15486 12852 15538
rect 12796 15484 12852 15486
rect 12796 15260 12852 15316
rect 12796 14028 12852 14084
rect 12908 14476 12964 14532
rect 13244 18172 13300 18228
rect 13692 19740 13748 19796
rect 13580 18562 13636 18564
rect 13580 18510 13582 18562
rect 13582 18510 13634 18562
rect 13634 18510 13636 18562
rect 13580 18508 13636 18510
rect 13468 17948 13524 18004
rect 13132 13916 13188 13972
rect 13356 16156 13412 16212
rect 14252 22540 14308 22596
rect 14476 21532 14532 21588
rect 14700 21420 14756 21476
rect 14364 21026 14420 21028
rect 14364 20974 14366 21026
rect 14366 20974 14418 21026
rect 14418 20974 14420 21026
rect 14364 20972 14420 20974
rect 14364 20802 14420 20804
rect 14364 20750 14366 20802
rect 14366 20750 14418 20802
rect 14418 20750 14420 20802
rect 14364 20748 14420 20750
rect 15148 22764 15204 22820
rect 15484 22988 15540 23044
rect 15372 22258 15428 22260
rect 15372 22206 15374 22258
rect 15374 22206 15426 22258
rect 15426 22206 15428 22258
rect 15372 22204 15428 22206
rect 15260 21474 15316 21476
rect 15260 21422 15262 21474
rect 15262 21422 15314 21474
rect 15314 21422 15316 21474
rect 15260 21420 15316 21422
rect 15260 20748 15316 20804
rect 14700 20524 14756 20580
rect 13804 18956 13860 19012
rect 14588 19964 14644 20020
rect 14812 20188 14868 20244
rect 14476 19404 14532 19460
rect 15036 20018 15092 20020
rect 15036 19966 15038 20018
rect 15038 19966 15090 20018
rect 15090 19966 15092 20018
rect 15036 19964 15092 19966
rect 14924 19740 14980 19796
rect 15036 19234 15092 19236
rect 15036 19182 15038 19234
rect 15038 19182 15090 19234
rect 15090 19182 15092 19234
rect 15036 19180 15092 19182
rect 13916 17164 13972 17220
rect 14476 18284 14532 18340
rect 13916 16828 13972 16884
rect 13804 16380 13860 16436
rect 13580 16044 13636 16100
rect 14364 17388 14420 17444
rect 14140 16044 14196 16100
rect 14252 16828 14308 16884
rect 14700 17666 14756 17668
rect 14700 17614 14702 17666
rect 14702 17614 14754 17666
rect 14754 17614 14756 17666
rect 14700 17612 14756 17614
rect 15148 17666 15204 17668
rect 15148 17614 15150 17666
rect 15150 17614 15202 17666
rect 15202 17614 15204 17666
rect 15148 17612 15204 17614
rect 16156 22764 16212 22820
rect 15932 21980 15988 22036
rect 15484 20076 15540 20132
rect 15372 17778 15428 17780
rect 15372 17726 15374 17778
rect 15374 17726 15426 17778
rect 15426 17726 15428 17778
rect 15372 17724 15428 17726
rect 14588 16716 14644 16772
rect 14700 17388 14756 17444
rect 14924 17164 14980 17220
rect 14812 16994 14868 16996
rect 14812 16942 14814 16994
rect 14814 16942 14866 16994
rect 14866 16942 14868 16994
rect 14812 16940 14868 16942
rect 14364 16658 14420 16660
rect 14364 16606 14366 16658
rect 14366 16606 14418 16658
rect 14418 16606 14420 16658
rect 14364 16604 14420 16606
rect 14588 16380 14644 16436
rect 14364 15932 14420 15988
rect 14812 16098 14868 16100
rect 14812 16046 14814 16098
rect 14814 16046 14866 16098
rect 14866 16046 14868 16098
rect 14812 16044 14868 16046
rect 14364 15708 14420 15764
rect 13468 15538 13524 15540
rect 13468 15486 13470 15538
rect 13470 15486 13522 15538
rect 13522 15486 13524 15538
rect 13468 15484 13524 15486
rect 13356 15372 13412 15428
rect 12908 12796 12964 12852
rect 12460 12012 12516 12068
rect 12460 11788 12516 11844
rect 12684 12066 12740 12068
rect 12684 12014 12686 12066
rect 12686 12014 12738 12066
rect 12738 12014 12740 12066
rect 12684 12012 12740 12014
rect 13804 14530 13860 14532
rect 13804 14478 13806 14530
rect 13806 14478 13858 14530
rect 13858 14478 13860 14530
rect 13804 14476 13860 14478
rect 13580 14306 13636 14308
rect 13580 14254 13582 14306
rect 13582 14254 13634 14306
rect 13634 14254 13636 14306
rect 13580 14252 13636 14254
rect 13468 14028 13524 14084
rect 13804 13970 13860 13972
rect 13804 13918 13806 13970
rect 13806 13918 13858 13970
rect 13858 13918 13860 13970
rect 13804 13916 13860 13918
rect 14140 14418 14196 14420
rect 14140 14366 14142 14418
rect 14142 14366 14194 14418
rect 14194 14366 14196 14418
rect 14140 14364 14196 14366
rect 13916 13804 13972 13860
rect 14140 13522 14196 13524
rect 14140 13470 14142 13522
rect 14142 13470 14194 13522
rect 14194 13470 14196 13522
rect 14140 13468 14196 13470
rect 13916 12962 13972 12964
rect 13916 12910 13918 12962
rect 13918 12910 13970 12962
rect 13970 12910 13972 12962
rect 13916 12908 13972 12910
rect 13580 12738 13636 12740
rect 13580 12686 13582 12738
rect 13582 12686 13634 12738
rect 13634 12686 13636 12738
rect 13580 12684 13636 12686
rect 14140 12850 14196 12852
rect 14140 12798 14142 12850
rect 14142 12798 14194 12850
rect 14194 12798 14196 12850
rect 14140 12796 14196 12798
rect 14924 14364 14980 14420
rect 14476 13858 14532 13860
rect 14476 13806 14478 13858
rect 14478 13806 14530 13858
rect 14530 13806 14532 13858
rect 14476 13804 14532 13806
rect 14700 12908 14756 12964
rect 13916 11788 13972 11844
rect 14812 11564 14868 11620
rect 15148 16716 15204 16772
rect 15260 15986 15316 15988
rect 15260 15934 15262 15986
rect 15262 15934 15314 15986
rect 15314 15934 15316 15986
rect 15260 15932 15316 15934
rect 15148 15820 15204 15876
rect 15148 15596 15204 15652
rect 15708 20018 15764 20020
rect 15708 19966 15710 20018
rect 15710 19966 15762 20018
rect 15762 19966 15764 20018
rect 15708 19964 15764 19966
rect 15932 19794 15988 19796
rect 15932 19742 15934 19794
rect 15934 19742 15986 19794
rect 15986 19742 15988 19794
rect 15932 19740 15988 19742
rect 16716 23042 16772 23044
rect 16716 22990 16718 23042
rect 16718 22990 16770 23042
rect 16770 22990 16772 23042
rect 16716 22988 16772 22990
rect 16716 21420 16772 21476
rect 16940 21420 16996 21476
rect 16604 20018 16660 20020
rect 16604 19966 16606 20018
rect 16606 19966 16658 20018
rect 16658 19966 16660 20018
rect 16604 19964 16660 19966
rect 16492 19404 16548 19460
rect 15708 19234 15764 19236
rect 15708 19182 15710 19234
rect 15710 19182 15762 19234
rect 15762 19182 15764 19234
rect 15708 19180 15764 19182
rect 15596 17948 15652 18004
rect 16156 18284 16212 18340
rect 16044 17948 16100 18004
rect 15596 17666 15652 17668
rect 15596 17614 15598 17666
rect 15598 17614 15650 17666
rect 15650 17614 15652 17666
rect 15596 17612 15652 17614
rect 15484 16882 15540 16884
rect 15484 16830 15486 16882
rect 15486 16830 15538 16882
rect 15538 16830 15540 16882
rect 15484 16828 15540 16830
rect 15820 16156 15876 16212
rect 16156 17778 16212 17780
rect 16156 17726 16158 17778
rect 16158 17726 16210 17778
rect 16210 17726 16212 17778
rect 16156 17724 16212 17726
rect 16156 17276 16212 17332
rect 16716 19180 16772 19236
rect 16604 17612 16660 17668
rect 16492 17052 16548 17108
rect 16940 17836 16996 17892
rect 16604 16940 16660 16996
rect 16828 16716 16884 16772
rect 16716 16604 16772 16660
rect 16044 16268 16100 16324
rect 16380 16268 16436 16324
rect 16828 16044 16884 16100
rect 15596 15202 15652 15204
rect 15596 15150 15598 15202
rect 15598 15150 15650 15202
rect 15650 15150 15652 15202
rect 15596 15148 15652 15150
rect 11900 8204 11956 8260
rect 12572 10668 12628 10724
rect 14588 11340 14644 11396
rect 14028 11282 14084 11284
rect 14028 11230 14030 11282
rect 14030 11230 14082 11282
rect 14082 11230 14084 11282
rect 14028 11228 14084 11230
rect 12908 8652 12964 8708
rect 12236 8092 12292 8148
rect 12572 8204 12628 8260
rect 13132 8204 13188 8260
rect 15036 9884 15092 9940
rect 15148 9324 15204 9380
rect 13692 8652 13748 8708
rect 14700 8818 14756 8820
rect 14700 8766 14702 8818
rect 14702 8766 14754 8818
rect 14754 8766 14756 8818
rect 14700 8764 14756 8766
rect 13580 8370 13636 8372
rect 13580 8318 13582 8370
rect 13582 8318 13634 8370
rect 13634 8318 13636 8370
rect 13580 8316 13636 8318
rect 11452 7196 11508 7252
rect 10108 6690 10164 6692
rect 10108 6638 10110 6690
rect 10110 6638 10162 6690
rect 10162 6638 10164 6690
rect 10108 6636 10164 6638
rect 12236 7250 12292 7252
rect 12236 7198 12238 7250
rect 12238 7198 12290 7250
rect 12290 7198 12292 7250
rect 12236 7196 12292 7198
rect 12236 6636 12292 6692
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 12908 7532 12964 7588
rect 13356 7586 13412 7588
rect 13356 7534 13358 7586
rect 13358 7534 13410 7586
rect 13410 7534 13412 7586
rect 13356 7532 13412 7534
rect 13244 7474 13300 7476
rect 13244 7422 13246 7474
rect 13246 7422 13298 7474
rect 13298 7422 13300 7474
rect 13244 7420 13300 7422
rect 12684 6636 12740 6692
rect 14140 8146 14196 8148
rect 14140 8094 14142 8146
rect 14142 8094 14194 8146
rect 14194 8094 14196 8146
rect 14140 8092 14196 8094
rect 13916 7532 13972 7588
rect 14700 7532 14756 7588
rect 14812 8092 14868 8148
rect 14812 7420 14868 7476
rect 16492 15820 16548 15876
rect 16380 15596 16436 15652
rect 15932 14700 15988 14756
rect 19516 30210 19572 30212
rect 19516 30158 19518 30210
rect 19518 30158 19570 30210
rect 19570 30158 19572 30210
rect 19516 30156 19572 30158
rect 18620 29036 18676 29092
rect 18844 29708 18900 29764
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19740 33068 19796 33124
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20748 38780 20804 38836
rect 20748 38108 20804 38164
rect 20860 39788 20916 39844
rect 21756 46674 21812 46676
rect 21756 46622 21758 46674
rect 21758 46622 21810 46674
rect 21810 46622 21812 46674
rect 21756 46620 21812 46622
rect 21756 46002 21812 46004
rect 21756 45950 21758 46002
rect 21758 45950 21810 46002
rect 21810 45950 21812 46002
rect 21756 45948 21812 45950
rect 21644 45836 21700 45892
rect 21308 42700 21364 42756
rect 21532 41970 21588 41972
rect 21532 41918 21534 41970
rect 21534 41918 21586 41970
rect 21586 41918 21588 41970
rect 21532 41916 21588 41918
rect 23212 48914 23268 48916
rect 23212 48862 23214 48914
rect 23214 48862 23266 48914
rect 23266 48862 23268 48914
rect 23212 48860 23268 48862
rect 23884 50540 23940 50596
rect 23660 49868 23716 49924
rect 24108 50428 24164 50484
rect 24556 52274 24612 52276
rect 24556 52222 24558 52274
rect 24558 52222 24610 52274
rect 24610 52222 24612 52274
rect 24556 52220 24612 52222
rect 25228 54348 25284 54404
rect 27804 55916 27860 55972
rect 26124 54908 26180 54964
rect 25788 54402 25844 54404
rect 25788 54350 25790 54402
rect 25790 54350 25842 54402
rect 25842 54350 25844 54402
rect 25788 54348 25844 54350
rect 29596 56252 29652 56308
rect 30716 56252 30772 56308
rect 29932 55970 29988 55972
rect 29932 55918 29934 55970
rect 29934 55918 29986 55970
rect 29986 55918 29988 55970
rect 29932 55916 29988 55918
rect 28252 54684 28308 54740
rect 29260 54738 29316 54740
rect 29260 54686 29262 54738
rect 29262 54686 29314 54738
rect 29314 54686 29316 54738
rect 29260 54684 29316 54686
rect 29148 54348 29204 54404
rect 29708 54402 29764 54404
rect 29708 54350 29710 54402
rect 29710 54350 29762 54402
rect 29762 54350 29764 54402
rect 29708 54348 29764 54350
rect 26460 54012 26516 54068
rect 28252 53900 28308 53956
rect 25340 53004 25396 53060
rect 25228 52220 25284 52276
rect 24332 51436 24388 51492
rect 25228 51660 25284 51716
rect 24444 51212 24500 51268
rect 25564 52722 25620 52724
rect 25564 52670 25566 52722
rect 25566 52670 25618 52722
rect 25618 52670 25620 52722
rect 25564 52668 25620 52670
rect 27132 52668 27188 52724
rect 25564 52444 25620 52500
rect 25452 50482 25508 50484
rect 25452 50430 25454 50482
rect 25454 50430 25506 50482
rect 25506 50430 25508 50482
rect 25452 50428 25508 50430
rect 24108 49196 24164 49252
rect 23884 48914 23940 48916
rect 23884 48862 23886 48914
rect 23886 48862 23938 48914
rect 23938 48862 23940 48914
rect 23884 48860 23940 48862
rect 22652 48300 22708 48356
rect 22540 47346 22596 47348
rect 22540 47294 22542 47346
rect 22542 47294 22594 47346
rect 22594 47294 22596 47346
rect 22540 47292 22596 47294
rect 23772 48354 23828 48356
rect 23772 48302 23774 48354
rect 23774 48302 23826 48354
rect 23826 48302 23828 48354
rect 23772 48300 23828 48302
rect 23100 48188 23156 48244
rect 22764 48130 22820 48132
rect 22764 48078 22766 48130
rect 22766 48078 22818 48130
rect 22818 48078 22820 48130
rect 22764 48076 22820 48078
rect 22988 48018 23044 48020
rect 22988 47966 22990 48018
rect 22990 47966 23042 48018
rect 23042 47966 23044 48018
rect 22988 47964 23044 47966
rect 22764 47740 22820 47796
rect 23548 48076 23604 48132
rect 22316 46508 22372 46564
rect 21980 46060 22036 46116
rect 22092 44940 22148 44996
rect 22204 43708 22260 43764
rect 21868 43372 21924 43428
rect 21868 43036 21924 43092
rect 22428 43762 22484 43764
rect 22428 43710 22430 43762
rect 22430 43710 22482 43762
rect 22482 43710 22484 43762
rect 22428 43708 22484 43710
rect 23100 46844 23156 46900
rect 21980 42028 22036 42084
rect 21644 41580 21700 41636
rect 21868 41916 21924 41972
rect 21308 41132 21364 41188
rect 21756 41020 21812 41076
rect 21644 40962 21700 40964
rect 21644 40910 21646 40962
rect 21646 40910 21698 40962
rect 21698 40910 21700 40962
rect 21644 40908 21700 40910
rect 21420 40236 21476 40292
rect 21084 39452 21140 39508
rect 20860 39004 20916 39060
rect 22092 42476 22148 42532
rect 21980 41186 22036 41188
rect 21980 41134 21982 41186
rect 21982 41134 22034 41186
rect 22034 41134 22036 41186
rect 21980 41132 22036 41134
rect 22204 42364 22260 42420
rect 22316 42140 22372 42196
rect 23212 46172 23268 46228
rect 22988 45890 23044 45892
rect 22988 45838 22990 45890
rect 22990 45838 23042 45890
rect 23042 45838 23044 45890
rect 22988 45836 23044 45838
rect 22988 45500 23044 45556
rect 23436 47068 23492 47124
rect 23660 47964 23716 48020
rect 25004 48860 25060 48916
rect 24668 48412 24724 48468
rect 24332 48242 24388 48244
rect 24332 48190 24334 48242
rect 24334 48190 24386 48242
rect 24386 48190 24388 48242
rect 24332 48188 24388 48190
rect 24332 47628 24388 47684
rect 24108 47234 24164 47236
rect 24108 47182 24110 47234
rect 24110 47182 24162 47234
rect 24162 47182 24164 47234
rect 24108 47180 24164 47182
rect 24556 47234 24612 47236
rect 24556 47182 24558 47234
rect 24558 47182 24610 47234
rect 24610 47182 24612 47234
rect 24556 47180 24612 47182
rect 23436 45052 23492 45108
rect 22988 44044 23044 44100
rect 24108 46898 24164 46900
rect 24108 46846 24110 46898
rect 24110 46846 24162 46898
rect 24162 46846 24164 46898
rect 24108 46844 24164 46846
rect 24220 46002 24276 46004
rect 24220 45950 24222 46002
rect 24222 45950 24274 46002
rect 24274 45950 24276 46002
rect 24220 45948 24276 45950
rect 23884 45500 23940 45556
rect 23996 45164 24052 45220
rect 23884 45106 23940 45108
rect 23884 45054 23886 45106
rect 23886 45054 23938 45106
rect 23938 45054 23940 45106
rect 23884 45052 23940 45054
rect 23212 43538 23268 43540
rect 23212 43486 23214 43538
rect 23214 43486 23266 43538
rect 23266 43486 23268 43538
rect 23212 43484 23268 43486
rect 23212 42642 23268 42644
rect 23212 42590 23214 42642
rect 23214 42590 23266 42642
rect 23266 42590 23268 42642
rect 23212 42588 23268 42590
rect 22204 41244 22260 41300
rect 22540 41468 22596 41524
rect 22652 41356 22708 41412
rect 23548 42924 23604 42980
rect 23100 41244 23156 41300
rect 22876 41132 22932 41188
rect 23324 41916 23380 41972
rect 23772 42812 23828 42868
rect 23660 42588 23716 42644
rect 23548 41746 23604 41748
rect 23548 41694 23550 41746
rect 23550 41694 23602 41746
rect 23602 41694 23604 41746
rect 23548 41692 23604 41694
rect 23660 41580 23716 41636
rect 23324 41298 23380 41300
rect 23324 41246 23326 41298
rect 23326 41246 23378 41298
rect 23378 41246 23380 41298
rect 23324 41244 23380 41246
rect 23436 41074 23492 41076
rect 23436 41022 23438 41074
rect 23438 41022 23490 41074
rect 23490 41022 23492 41074
rect 23436 41020 23492 41022
rect 24668 45388 24724 45444
rect 24332 45276 24388 45332
rect 24220 44268 24276 44324
rect 24220 43650 24276 43652
rect 24220 43598 24222 43650
rect 24222 43598 24274 43650
rect 24274 43598 24276 43650
rect 24220 43596 24276 43598
rect 24220 43372 24276 43428
rect 24108 42924 24164 42980
rect 24556 43426 24612 43428
rect 24556 43374 24558 43426
rect 24558 43374 24610 43426
rect 24610 43374 24612 43426
rect 24556 43372 24612 43374
rect 24668 43036 24724 43092
rect 25116 48748 25172 48804
rect 25116 46844 25172 46900
rect 25004 46396 25060 46452
rect 25004 44434 25060 44436
rect 25004 44382 25006 44434
rect 25006 44382 25058 44434
rect 25058 44382 25060 44434
rect 25004 44380 25060 44382
rect 25116 43148 25172 43204
rect 24444 42588 24500 42644
rect 24108 41244 24164 41300
rect 22092 40908 22148 40964
rect 21868 39788 21924 39844
rect 21308 39676 21364 39732
rect 21868 39452 21924 39508
rect 21756 38834 21812 38836
rect 21756 38782 21758 38834
rect 21758 38782 21810 38834
rect 21810 38782 21812 38834
rect 21756 38780 21812 38782
rect 21756 38556 21812 38612
rect 21756 38162 21812 38164
rect 21756 38110 21758 38162
rect 21758 38110 21810 38162
rect 21810 38110 21812 38162
rect 21756 38108 21812 38110
rect 22092 40236 22148 40292
rect 21420 37324 21476 37380
rect 21308 37212 21364 37268
rect 21644 37266 21700 37268
rect 21644 37214 21646 37266
rect 21646 37214 21698 37266
rect 21698 37214 21700 37266
rect 21644 37212 21700 37214
rect 20636 37100 20692 37156
rect 20636 36764 20692 36820
rect 20524 36482 20580 36484
rect 20524 36430 20526 36482
rect 20526 36430 20578 36482
rect 20578 36430 20580 36482
rect 20524 36428 20580 36430
rect 21756 36428 21812 36484
rect 21308 36092 21364 36148
rect 20748 35868 20804 35924
rect 20748 35308 20804 35364
rect 20412 33964 20468 34020
rect 20412 33740 20468 33796
rect 21308 34914 21364 34916
rect 21308 34862 21310 34914
rect 21310 34862 21362 34914
rect 21362 34862 21364 34914
rect 21308 34860 21364 34862
rect 20748 34802 20804 34804
rect 20748 34750 20750 34802
rect 20750 34750 20802 34802
rect 20802 34750 20804 34802
rect 20748 34748 20804 34750
rect 22428 40572 22484 40628
rect 22316 40514 22372 40516
rect 22316 40462 22318 40514
rect 22318 40462 22370 40514
rect 22370 40462 22372 40514
rect 22316 40460 22372 40462
rect 22876 40348 22932 40404
rect 22428 39618 22484 39620
rect 22428 39566 22430 39618
rect 22430 39566 22482 39618
rect 22482 39566 22484 39618
rect 22428 39564 22484 39566
rect 22540 39228 22596 39284
rect 22428 37266 22484 37268
rect 22428 37214 22430 37266
rect 22430 37214 22482 37266
rect 22482 37214 22484 37266
rect 22428 37212 22484 37214
rect 22204 36428 22260 36484
rect 22428 36316 22484 36372
rect 22204 35980 22260 36036
rect 21980 34802 22036 34804
rect 21980 34750 21982 34802
rect 21982 34750 22034 34802
rect 22034 34750 22036 34802
rect 21980 34748 22036 34750
rect 20860 34130 20916 34132
rect 20860 34078 20862 34130
rect 20862 34078 20914 34130
rect 20914 34078 20916 34130
rect 20860 34076 20916 34078
rect 21308 34018 21364 34020
rect 21308 33966 21310 34018
rect 21310 33966 21362 34018
rect 21362 33966 21364 34018
rect 21308 33964 21364 33966
rect 20524 33628 20580 33684
rect 21756 33628 21812 33684
rect 20524 33122 20580 33124
rect 20524 33070 20526 33122
rect 20526 33070 20578 33122
rect 20578 33070 20580 33122
rect 20524 33068 20580 33070
rect 21420 32956 21476 33012
rect 20524 31778 20580 31780
rect 20524 31726 20526 31778
rect 20526 31726 20578 31778
rect 20578 31726 20580 31778
rect 20524 31724 20580 31726
rect 20412 31666 20468 31668
rect 20412 31614 20414 31666
rect 20414 31614 20466 31666
rect 20466 31614 20468 31666
rect 20412 31612 20468 31614
rect 20748 31666 20804 31668
rect 20748 31614 20750 31666
rect 20750 31614 20802 31666
rect 20802 31614 20804 31666
rect 20748 31612 20804 31614
rect 20076 31500 20132 31556
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 21308 31500 21364 31556
rect 21308 30828 21364 30884
rect 21644 30210 21700 30212
rect 21644 30158 21646 30210
rect 21646 30158 21698 30210
rect 21698 30158 21700 30210
rect 21644 30156 21700 30158
rect 20076 29932 20132 29988
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 22428 35420 22484 35476
rect 23884 40124 23940 40180
rect 23548 39730 23604 39732
rect 23548 39678 23550 39730
rect 23550 39678 23602 39730
rect 23602 39678 23604 39730
rect 23548 39676 23604 39678
rect 22988 39340 23044 39396
rect 23100 39228 23156 39284
rect 22988 38668 23044 38724
rect 22988 38332 23044 38388
rect 22988 38162 23044 38164
rect 22988 38110 22990 38162
rect 22990 38110 23042 38162
rect 23042 38110 23044 38162
rect 22988 38108 23044 38110
rect 22988 37490 23044 37492
rect 22988 37438 22990 37490
rect 22990 37438 23042 37490
rect 23042 37438 23044 37490
rect 22988 37436 23044 37438
rect 22876 35980 22932 36036
rect 23996 38444 24052 38500
rect 23996 37938 24052 37940
rect 23996 37886 23998 37938
rect 23998 37886 24050 37938
rect 24050 37886 24052 37938
rect 23996 37884 24052 37886
rect 24108 37436 24164 37492
rect 23324 36988 23380 37044
rect 22988 35868 23044 35924
rect 23212 35980 23268 36036
rect 23324 35644 23380 35700
rect 25004 40908 25060 40964
rect 24668 40626 24724 40628
rect 24668 40574 24670 40626
rect 24670 40574 24722 40626
rect 24722 40574 24724 40626
rect 24668 40572 24724 40574
rect 25340 47628 25396 47684
rect 25452 47068 25508 47124
rect 25340 46674 25396 46676
rect 25340 46622 25342 46674
rect 25342 46622 25394 46674
rect 25394 46622 25396 46674
rect 25340 46620 25396 46622
rect 27356 51266 27412 51268
rect 27356 51214 27358 51266
rect 27358 51214 27410 51266
rect 27410 51214 27412 51266
rect 27356 51212 27412 51214
rect 26908 50428 26964 50484
rect 26796 48636 26852 48692
rect 25676 48524 25732 48580
rect 25788 48412 25844 48468
rect 26460 48412 26516 48468
rect 26012 48242 26068 48244
rect 26012 48190 26014 48242
rect 26014 48190 26066 48242
rect 26066 48190 26068 48242
rect 26012 48188 26068 48190
rect 26684 48076 26740 48132
rect 25676 47682 25732 47684
rect 25676 47630 25678 47682
rect 25678 47630 25730 47682
rect 25730 47630 25732 47682
rect 25676 47628 25732 47630
rect 26684 47628 26740 47684
rect 25676 47180 25732 47236
rect 26012 47292 26068 47348
rect 25564 45500 25620 45556
rect 25676 45388 25732 45444
rect 25900 45612 25956 45668
rect 26236 47068 26292 47124
rect 26012 45500 26068 45556
rect 26572 46060 26628 46116
rect 26796 46450 26852 46452
rect 26796 46398 26798 46450
rect 26798 46398 26850 46450
rect 26850 46398 26852 46450
rect 26796 46396 26852 46398
rect 28588 51548 28644 51604
rect 27580 49084 27636 49140
rect 27244 47740 27300 47796
rect 27356 48636 27412 48692
rect 27244 47570 27300 47572
rect 27244 47518 27246 47570
rect 27246 47518 27298 47570
rect 27298 47518 27300 47570
rect 27244 47516 27300 47518
rect 28476 49084 28532 49140
rect 27804 49026 27860 49028
rect 27804 48974 27806 49026
rect 27806 48974 27858 49026
rect 27858 48974 27860 49026
rect 27804 48972 27860 48974
rect 27580 48524 27636 48580
rect 28252 48802 28308 48804
rect 28252 48750 28254 48802
rect 28254 48750 28306 48802
rect 28306 48750 28308 48802
rect 28252 48748 28308 48750
rect 27916 48076 27972 48132
rect 28364 48076 28420 48132
rect 27692 47458 27748 47460
rect 27692 47406 27694 47458
rect 27694 47406 27746 47458
rect 27746 47406 27748 47458
rect 27692 47404 27748 47406
rect 27692 47180 27748 47236
rect 28028 47292 28084 47348
rect 27132 46844 27188 46900
rect 27020 46060 27076 46116
rect 26348 45276 26404 45332
rect 25900 44044 25956 44100
rect 26236 43932 26292 43988
rect 25788 43820 25844 43876
rect 26796 45164 26852 45220
rect 26684 45106 26740 45108
rect 26684 45054 26686 45106
rect 26686 45054 26738 45106
rect 26738 45054 26740 45106
rect 26684 45052 26740 45054
rect 27468 46060 27524 46116
rect 27580 46396 27636 46452
rect 27244 45666 27300 45668
rect 27244 45614 27246 45666
rect 27246 45614 27298 45666
rect 27298 45614 27300 45666
rect 27244 45612 27300 45614
rect 27692 45724 27748 45780
rect 27020 45388 27076 45444
rect 27244 44828 27300 44884
rect 26908 44604 26964 44660
rect 27356 44322 27412 44324
rect 27356 44270 27358 44322
rect 27358 44270 27410 44322
rect 27410 44270 27412 44322
rect 27356 44268 27412 44270
rect 25452 43596 25508 43652
rect 25340 43260 25396 43316
rect 25788 43260 25844 43316
rect 25452 42754 25508 42756
rect 25452 42702 25454 42754
rect 25454 42702 25506 42754
rect 25506 42702 25508 42754
rect 25452 42700 25508 42702
rect 25676 43148 25732 43204
rect 25340 40962 25396 40964
rect 25340 40910 25342 40962
rect 25342 40910 25394 40962
rect 25394 40910 25396 40962
rect 25340 40908 25396 40910
rect 24668 38444 24724 38500
rect 25340 39618 25396 39620
rect 25340 39566 25342 39618
rect 25342 39566 25394 39618
rect 25394 39566 25396 39618
rect 25340 39564 25396 39566
rect 25452 38556 25508 38612
rect 22764 35196 22820 35252
rect 21868 32956 21924 33012
rect 22428 32956 22484 33012
rect 22316 32508 22372 32564
rect 21868 31890 21924 31892
rect 21868 31838 21870 31890
rect 21870 31838 21922 31890
rect 21922 31838 21924 31890
rect 21868 31836 21924 31838
rect 22540 31724 22596 31780
rect 21980 31612 22036 31668
rect 21868 30380 21924 30436
rect 18396 28530 18452 28532
rect 18396 28478 18398 28530
rect 18398 28478 18450 28530
rect 18450 28478 18452 28530
rect 18396 28476 18452 28478
rect 18620 27692 18676 27748
rect 17276 23772 17332 23828
rect 17500 23324 17556 23380
rect 17724 23772 17780 23828
rect 18172 25228 18228 25284
rect 18732 25282 18788 25284
rect 18732 25230 18734 25282
rect 18734 25230 18786 25282
rect 18786 25230 18788 25282
rect 18732 25228 18788 25230
rect 18396 25116 18452 25172
rect 19180 28476 19236 28532
rect 19068 28364 19124 28420
rect 18956 27634 19012 27636
rect 18956 27582 18958 27634
rect 18958 27582 19010 27634
rect 19010 27582 19012 27634
rect 18956 27580 19012 27582
rect 21756 29596 21812 29652
rect 21868 29708 21924 29764
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19740 27692 19796 27748
rect 22428 30380 22484 30436
rect 22316 30156 22372 30212
rect 22988 30156 23044 30212
rect 22876 30098 22932 30100
rect 22876 30046 22878 30098
rect 22878 30046 22930 30098
rect 22930 30046 22932 30098
rect 22876 30044 22932 30046
rect 21420 28418 21476 28420
rect 21420 28366 21422 28418
rect 21422 28366 21474 28418
rect 21474 28366 21476 28418
rect 21420 28364 21476 28366
rect 21756 28364 21812 28420
rect 21532 27468 21588 27524
rect 20524 27074 20580 27076
rect 20524 27022 20526 27074
rect 20526 27022 20578 27074
rect 20578 27022 20580 27074
rect 20524 27020 20580 27022
rect 20076 26796 20132 26852
rect 18508 24834 18564 24836
rect 18508 24782 18510 24834
rect 18510 24782 18562 24834
rect 18562 24782 18564 24834
rect 18508 24780 18564 24782
rect 17724 22316 17780 22372
rect 17948 24444 18004 24500
rect 18284 23436 18340 23492
rect 18172 23324 18228 23380
rect 18060 23154 18116 23156
rect 18060 23102 18062 23154
rect 18062 23102 18114 23154
rect 18114 23102 18116 23154
rect 18060 23100 18116 23102
rect 17948 22204 18004 22260
rect 18284 21980 18340 22036
rect 17500 21474 17556 21476
rect 17500 21422 17502 21474
rect 17502 21422 17554 21474
rect 17554 21422 17556 21474
rect 17500 21420 17556 21422
rect 17612 21196 17668 21252
rect 17388 20972 17444 21028
rect 18060 21196 18116 21252
rect 17612 20188 17668 20244
rect 17836 20972 17892 21028
rect 17388 19964 17444 20020
rect 17612 19740 17668 19796
rect 17500 18396 17556 18452
rect 17948 18338 18004 18340
rect 17948 18286 17950 18338
rect 17950 18286 18002 18338
rect 18002 18286 18004 18338
rect 17948 18284 18004 18286
rect 17388 16492 17444 16548
rect 17500 16940 17556 16996
rect 18060 17724 18116 17780
rect 18172 20972 18228 21028
rect 19516 26684 19572 26740
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19516 26124 19572 26180
rect 19068 25116 19124 25172
rect 18956 24444 19012 24500
rect 18732 23826 18788 23828
rect 18732 23774 18734 23826
rect 18734 23774 18786 23826
rect 18786 23774 18788 23826
rect 18732 23772 18788 23774
rect 18620 23324 18676 23380
rect 18396 21644 18452 21700
rect 18508 21196 18564 21252
rect 19292 23660 19348 23716
rect 20636 26460 20692 26516
rect 20300 25340 20356 25396
rect 19964 25228 20020 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19628 24444 19684 24500
rect 19516 23324 19572 23380
rect 19628 23772 19684 23828
rect 18732 22370 18788 22372
rect 18732 22318 18734 22370
rect 18734 22318 18786 22370
rect 18786 22318 18788 22370
rect 18732 22316 18788 22318
rect 19068 22258 19124 22260
rect 19068 22206 19070 22258
rect 19070 22206 19122 22258
rect 19122 22206 19124 22258
rect 19068 22204 19124 22206
rect 18956 21084 19012 21140
rect 18284 20412 18340 20468
rect 18172 18060 18228 18116
rect 17836 16940 17892 16996
rect 17948 16828 18004 16884
rect 17612 16716 17668 16772
rect 18284 18396 18340 18452
rect 18396 18338 18452 18340
rect 18396 18286 18398 18338
rect 18398 18286 18450 18338
rect 18450 18286 18452 18338
rect 18396 18284 18452 18286
rect 18172 16716 18228 16772
rect 18284 16268 18340 16324
rect 17164 15874 17220 15876
rect 17164 15822 17166 15874
rect 17166 15822 17218 15874
rect 17218 15822 17220 15874
rect 17164 15820 17220 15822
rect 17052 15596 17108 15652
rect 18060 16098 18116 16100
rect 18060 16046 18062 16098
rect 18062 16046 18114 16098
rect 18114 16046 18116 16098
rect 18060 16044 18116 16046
rect 16828 14700 16884 14756
rect 19516 23100 19572 23156
rect 19964 23660 20020 23716
rect 20748 25228 20804 25284
rect 20748 24946 20804 24948
rect 20748 24894 20750 24946
rect 20750 24894 20802 24946
rect 20802 24894 20804 24946
rect 20748 24892 20804 24894
rect 21196 26124 21252 26180
rect 21196 25228 21252 25284
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19852 23324 19908 23380
rect 20188 23324 20244 23380
rect 20300 23660 20356 23716
rect 20076 23266 20132 23268
rect 20076 23214 20078 23266
rect 20078 23214 20130 23266
rect 20130 23214 20132 23266
rect 20076 23212 20132 23214
rect 20300 23212 20356 23268
rect 20412 23436 20468 23492
rect 19852 22428 19908 22484
rect 20748 23324 20804 23380
rect 22764 28588 22820 28644
rect 22092 27468 22148 27524
rect 22988 27746 23044 27748
rect 22988 27694 22990 27746
rect 22990 27694 23042 27746
rect 23042 27694 23044 27746
rect 22988 27692 23044 27694
rect 22540 27468 22596 27524
rect 21644 26460 21700 26516
rect 22540 27074 22596 27076
rect 22540 27022 22542 27074
rect 22542 27022 22594 27074
rect 22594 27022 22596 27074
rect 22540 27020 22596 27022
rect 23884 35698 23940 35700
rect 23884 35646 23886 35698
rect 23886 35646 23938 35698
rect 23938 35646 23940 35698
rect 23884 35644 23940 35646
rect 23772 35084 23828 35140
rect 25788 41244 25844 41300
rect 25676 39788 25732 39844
rect 24556 36988 24612 37044
rect 26012 43036 26068 43092
rect 26348 43484 26404 43540
rect 26684 43932 26740 43988
rect 26572 43820 26628 43876
rect 26124 42700 26180 42756
rect 26460 42754 26516 42756
rect 26460 42702 26462 42754
rect 26462 42702 26514 42754
rect 26514 42702 26516 42754
rect 26460 42700 26516 42702
rect 26236 42642 26292 42644
rect 26236 42590 26238 42642
rect 26238 42590 26290 42642
rect 26290 42590 26292 42642
rect 26236 42588 26292 42590
rect 26012 42530 26068 42532
rect 26012 42478 26014 42530
rect 26014 42478 26066 42530
rect 26066 42478 26068 42530
rect 26012 42476 26068 42478
rect 26012 41580 26068 41636
rect 26236 41356 26292 41412
rect 26236 40572 26292 40628
rect 26572 41132 26628 41188
rect 26460 40348 26516 40404
rect 27356 43932 27412 43988
rect 26796 43820 26852 43876
rect 26908 43708 26964 43764
rect 26796 43260 26852 43316
rect 27020 43650 27076 43652
rect 27020 43598 27022 43650
rect 27022 43598 27074 43650
rect 27074 43598 27076 43650
rect 27020 43596 27076 43598
rect 27132 43426 27188 43428
rect 27132 43374 27134 43426
rect 27134 43374 27186 43426
rect 27186 43374 27188 43426
rect 27132 43372 27188 43374
rect 29484 49084 29540 49140
rect 29148 49026 29204 49028
rect 29148 48974 29150 49026
rect 29150 48974 29202 49026
rect 29202 48974 29204 49026
rect 29148 48972 29204 48974
rect 30940 56252 30996 56308
rect 32284 57036 32340 57092
rect 32620 56252 32676 56308
rect 30380 53564 30436 53620
rect 30940 54348 30996 54404
rect 32060 54402 32116 54404
rect 32060 54350 32062 54402
rect 32062 54350 32114 54402
rect 32114 54350 32116 54402
rect 32060 54348 32116 54350
rect 33628 56924 33684 56980
rect 34076 56252 34132 56308
rect 34188 57036 34244 57092
rect 32508 54402 32564 54404
rect 32508 54350 32510 54402
rect 32510 54350 32562 54402
rect 32562 54350 32564 54402
rect 32508 54348 32564 54350
rect 33852 56028 33908 56084
rect 34972 57036 35028 57092
rect 35308 56306 35364 56308
rect 35308 56254 35310 56306
rect 35310 56254 35362 56306
rect 35362 56254 35364 56306
rect 35308 56252 35364 56254
rect 35980 56082 36036 56084
rect 35980 56030 35982 56082
rect 35982 56030 36034 56082
rect 36034 56030 36036 56082
rect 35980 56028 36036 56030
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35308 55468 35364 55524
rect 36428 56924 36484 56980
rect 37660 56700 37716 56756
rect 37996 57036 38052 57092
rect 36764 56252 36820 56308
rect 37548 55468 37604 55524
rect 36316 55356 36372 55412
rect 37436 55410 37492 55412
rect 37436 55358 37438 55410
rect 37438 55358 37490 55410
rect 37490 55358 37492 55410
rect 37436 55356 37492 55358
rect 33180 53116 33236 53172
rect 32284 52946 32340 52948
rect 32284 52894 32286 52946
rect 32286 52894 32338 52946
rect 32338 52894 32340 52946
rect 32284 52892 32340 52894
rect 33516 54012 33572 54068
rect 31164 51996 31220 52052
rect 30492 51548 30548 51604
rect 31836 51602 31892 51604
rect 31836 51550 31838 51602
rect 31838 51550 31890 51602
rect 31890 51550 31892 51602
rect 31836 51548 31892 51550
rect 34188 54348 34244 54404
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 39004 56812 39060 56868
rect 39116 56306 39172 56308
rect 39116 56254 39118 56306
rect 39118 56254 39170 56306
rect 39170 56254 39172 56306
rect 39116 56252 39172 56254
rect 39116 54290 39172 54292
rect 39116 54238 39118 54290
rect 39118 54238 39170 54290
rect 39170 54238 39172 54290
rect 39116 54236 39172 54238
rect 34076 53340 34132 53396
rect 33964 53170 34020 53172
rect 33964 53118 33966 53170
rect 33966 53118 34018 53170
rect 34018 53118 34020 53170
rect 33964 53116 34020 53118
rect 34748 53564 34804 53620
rect 34524 53228 34580 53284
rect 34188 51490 34244 51492
rect 34188 51438 34190 51490
rect 34190 51438 34242 51490
rect 34242 51438 34244 51490
rect 34188 51436 34244 51438
rect 34412 51378 34468 51380
rect 34412 51326 34414 51378
rect 34414 51326 34466 51378
rect 34466 51326 34468 51378
rect 34412 51324 34468 51326
rect 30492 49698 30548 49700
rect 30492 49646 30494 49698
rect 30494 49646 30546 49698
rect 30546 49646 30548 49698
rect 30492 49644 30548 49646
rect 30156 49196 30212 49252
rect 30380 49084 30436 49140
rect 28924 48860 28980 48916
rect 29372 48748 29428 48804
rect 28700 48242 28756 48244
rect 28700 48190 28702 48242
rect 28702 48190 28754 48242
rect 28754 48190 28756 48242
rect 28700 48188 28756 48190
rect 28700 47852 28756 47908
rect 28028 46674 28084 46676
rect 28028 46622 28030 46674
rect 28030 46622 28082 46674
rect 28082 46622 28084 46674
rect 28028 46620 28084 46622
rect 28476 47180 28532 47236
rect 28588 46786 28644 46788
rect 28588 46734 28590 46786
rect 28590 46734 28642 46786
rect 28642 46734 28644 46786
rect 28588 46732 28644 46734
rect 29708 48802 29764 48804
rect 29708 48750 29710 48802
rect 29710 48750 29762 48802
rect 29762 48750 29764 48802
rect 29708 48748 29764 48750
rect 30716 49868 30772 49924
rect 31164 49868 31220 49924
rect 30828 49644 30884 49700
rect 29148 48130 29204 48132
rect 29148 48078 29150 48130
rect 29150 48078 29202 48130
rect 29202 48078 29204 48130
rect 29148 48076 29204 48078
rect 29260 47964 29316 48020
rect 29036 47458 29092 47460
rect 29036 47406 29038 47458
rect 29038 47406 29090 47458
rect 29090 47406 29092 47458
rect 29036 47404 29092 47406
rect 28924 46956 28980 47012
rect 29260 46786 29316 46788
rect 29260 46734 29262 46786
rect 29262 46734 29314 46786
rect 29314 46734 29316 46786
rect 29260 46732 29316 46734
rect 28028 45890 28084 45892
rect 28028 45838 28030 45890
rect 28030 45838 28082 45890
rect 28082 45838 28084 45890
rect 28028 45836 28084 45838
rect 28140 45948 28196 46004
rect 27804 43932 27860 43988
rect 27916 43708 27972 43764
rect 28252 45388 28308 45444
rect 29484 46844 29540 46900
rect 29484 46508 29540 46564
rect 29708 47740 29764 47796
rect 29820 47516 29876 47572
rect 30940 48412 30996 48468
rect 29708 46898 29764 46900
rect 29708 46846 29710 46898
rect 29710 46846 29762 46898
rect 29762 46846 29764 46898
rect 29708 46844 29764 46846
rect 30156 46898 30212 46900
rect 30156 46846 30158 46898
rect 30158 46846 30210 46898
rect 30210 46846 30212 46898
rect 30156 46844 30212 46846
rect 29596 46732 29652 46788
rect 28364 44380 28420 44436
rect 29372 45388 29428 45444
rect 29148 45276 29204 45332
rect 28476 44828 28532 44884
rect 28252 44322 28308 44324
rect 28252 44270 28254 44322
rect 28254 44270 28306 44322
rect 28306 44270 28308 44322
rect 28252 44268 28308 44270
rect 28588 44492 28644 44548
rect 28140 43820 28196 43876
rect 29260 45052 29316 45108
rect 30828 46844 30884 46900
rect 30940 46786 30996 46788
rect 30940 46734 30942 46786
rect 30942 46734 30994 46786
rect 30994 46734 30996 46786
rect 30940 46732 30996 46734
rect 33964 51212 34020 51268
rect 34412 50652 34468 50708
rect 34300 50540 34356 50596
rect 32172 49922 32228 49924
rect 32172 49870 32174 49922
rect 32174 49870 32226 49922
rect 32226 49870 32228 49922
rect 32172 49868 32228 49870
rect 34860 51996 34916 52052
rect 35196 53564 35252 53620
rect 35308 53004 35364 53060
rect 35308 52668 35364 52724
rect 35420 52780 35476 52836
rect 35868 53228 35924 53284
rect 38556 53842 38612 53844
rect 38556 53790 38558 53842
rect 38558 53790 38610 53842
rect 38610 53790 38612 53842
rect 38556 53788 38612 53790
rect 37884 53676 37940 53732
rect 38332 53676 38388 53732
rect 37996 53564 38052 53620
rect 37212 52946 37268 52948
rect 37212 52894 37214 52946
rect 37214 52894 37266 52946
rect 37266 52894 37268 52946
rect 37212 52892 37268 52894
rect 37884 52892 37940 52948
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35644 52444 35700 52500
rect 35532 52220 35588 52276
rect 35308 51884 35364 51940
rect 34972 51212 35028 51268
rect 36316 52668 36372 52724
rect 36204 52332 36260 52388
rect 35756 52050 35812 52052
rect 35756 51998 35758 52050
rect 35758 51998 35810 52050
rect 35810 51998 35812 52050
rect 35756 51996 35812 51998
rect 36316 52220 36372 52276
rect 36316 51996 36372 52052
rect 35532 51548 35588 51604
rect 35420 51490 35476 51492
rect 35420 51438 35422 51490
rect 35422 51438 35474 51490
rect 35474 51438 35476 51490
rect 35420 51436 35476 51438
rect 34748 51100 34804 51156
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35084 50428 35140 50484
rect 31276 49698 31332 49700
rect 31276 49646 31278 49698
rect 31278 49646 31330 49698
rect 31330 49646 31332 49698
rect 31276 49644 31332 49646
rect 31276 49026 31332 49028
rect 31276 48974 31278 49026
rect 31278 48974 31330 49026
rect 31330 48974 31332 49026
rect 31276 48972 31332 48974
rect 35420 50594 35476 50596
rect 35420 50542 35422 50594
rect 35422 50542 35474 50594
rect 35474 50542 35476 50594
rect 35420 50540 35476 50542
rect 34860 49810 34916 49812
rect 34860 49758 34862 49810
rect 34862 49758 34914 49810
rect 34914 49758 34916 49810
rect 34860 49756 34916 49758
rect 35644 51378 35700 51380
rect 35644 51326 35646 51378
rect 35646 51326 35698 51378
rect 35698 51326 35700 51378
rect 35644 51324 35700 51326
rect 35644 50988 35700 51044
rect 35644 49756 35700 49812
rect 34300 49420 34356 49476
rect 33964 48972 34020 49028
rect 31948 48914 32004 48916
rect 31948 48862 31950 48914
rect 31950 48862 32002 48914
rect 32002 48862 32004 48914
rect 31948 48860 32004 48862
rect 33404 48860 33460 48916
rect 33180 48300 33236 48356
rect 31836 48188 31892 48244
rect 32508 48242 32564 48244
rect 32508 48190 32510 48242
rect 32510 48190 32562 48242
rect 32562 48190 32564 48242
rect 32508 48188 32564 48190
rect 33068 47852 33124 47908
rect 31388 47404 31444 47460
rect 32732 47458 32788 47460
rect 32732 47406 32734 47458
rect 32734 47406 32786 47458
rect 32786 47406 32788 47458
rect 32732 47404 32788 47406
rect 33292 48242 33348 48244
rect 33292 48190 33294 48242
rect 33294 48190 33346 48242
rect 33346 48190 33348 48242
rect 33292 48188 33348 48190
rect 33292 47068 33348 47124
rect 31164 46786 31220 46788
rect 31164 46734 31166 46786
rect 31166 46734 31218 46786
rect 31218 46734 31220 46786
rect 31164 46732 31220 46734
rect 32508 46956 32564 47012
rect 31052 46620 31108 46676
rect 31276 46674 31332 46676
rect 31276 46622 31278 46674
rect 31278 46622 31330 46674
rect 31330 46622 31332 46674
rect 31276 46620 31332 46622
rect 30156 45778 30212 45780
rect 30156 45726 30158 45778
rect 30158 45726 30210 45778
rect 30210 45726 30212 45778
rect 30156 45724 30212 45726
rect 30044 45164 30100 45220
rect 29820 45052 29876 45108
rect 29596 44492 29652 44548
rect 28140 43596 28196 43652
rect 27468 43036 27524 43092
rect 27356 42924 27412 42980
rect 27132 42700 27188 42756
rect 27132 42082 27188 42084
rect 27132 42030 27134 42082
rect 27134 42030 27186 42082
rect 27186 42030 27188 42082
rect 27132 42028 27188 42030
rect 26796 41804 26852 41860
rect 27580 42588 27636 42644
rect 27916 42812 27972 42868
rect 27468 42194 27524 42196
rect 27468 42142 27470 42194
rect 27470 42142 27522 42194
rect 27522 42142 27524 42194
rect 27468 42140 27524 42142
rect 27244 41804 27300 41860
rect 27692 41858 27748 41860
rect 27692 41806 27694 41858
rect 27694 41806 27746 41858
rect 27746 41806 27748 41858
rect 27692 41804 27748 41806
rect 28028 42364 28084 42420
rect 26684 40124 26740 40180
rect 27580 41410 27636 41412
rect 27580 41358 27582 41410
rect 27582 41358 27634 41410
rect 27634 41358 27636 41410
rect 27580 41356 27636 41358
rect 26908 40236 26964 40292
rect 26908 39900 26964 39956
rect 26572 39618 26628 39620
rect 26572 39566 26574 39618
rect 26574 39566 26626 39618
rect 26626 39566 26628 39618
rect 26572 39564 26628 39566
rect 26012 39506 26068 39508
rect 26012 39454 26014 39506
rect 26014 39454 26066 39506
rect 26066 39454 26068 39506
rect 26012 39452 26068 39454
rect 26684 39004 26740 39060
rect 26012 38556 26068 38612
rect 25900 37884 25956 37940
rect 24444 35756 24500 35812
rect 24892 35868 24948 35924
rect 24556 35084 24612 35140
rect 23772 34188 23828 34244
rect 24668 34300 24724 34356
rect 24332 33906 24388 33908
rect 24332 33854 24334 33906
rect 24334 33854 24386 33906
rect 24386 33854 24388 33906
rect 24332 33852 24388 33854
rect 23324 32956 23380 33012
rect 23324 30380 23380 30436
rect 24892 33068 24948 33124
rect 23660 32956 23716 33012
rect 24444 32956 24500 33012
rect 23660 32562 23716 32564
rect 23660 32510 23662 32562
rect 23662 32510 23714 32562
rect 23714 32510 23716 32562
rect 23660 32508 23716 32510
rect 25004 31666 25060 31668
rect 25004 31614 25006 31666
rect 25006 31614 25058 31666
rect 25058 31614 25060 31666
rect 25004 31612 25060 31614
rect 24668 31218 24724 31220
rect 24668 31166 24670 31218
rect 24670 31166 24722 31218
rect 24722 31166 24724 31218
rect 24668 31164 24724 31166
rect 23436 29708 23492 29764
rect 24108 30044 24164 30100
rect 23436 28642 23492 28644
rect 23436 28590 23438 28642
rect 23438 28590 23490 28642
rect 23490 28590 23492 28642
rect 23436 28588 23492 28590
rect 23436 27692 23492 27748
rect 21756 26796 21812 26852
rect 21644 26012 21700 26068
rect 21420 25228 21476 25284
rect 22428 26572 22484 26628
rect 22652 26850 22708 26852
rect 22652 26798 22654 26850
rect 22654 26798 22706 26850
rect 22706 26798 22708 26850
rect 22652 26796 22708 26798
rect 23212 26572 23268 26628
rect 22540 26402 22596 26404
rect 22540 26350 22542 26402
rect 22542 26350 22594 26402
rect 22594 26350 22596 26402
rect 22540 26348 22596 26350
rect 23100 26290 23156 26292
rect 23100 26238 23102 26290
rect 23102 26238 23154 26290
rect 23154 26238 23156 26290
rect 23100 26236 23156 26238
rect 22988 26012 23044 26068
rect 22540 25340 22596 25396
rect 21980 25282 22036 25284
rect 21980 25230 21982 25282
rect 21982 25230 22034 25282
rect 22034 25230 22036 25282
rect 21980 25228 22036 25230
rect 23996 27858 24052 27860
rect 23996 27806 23998 27858
rect 23998 27806 24050 27858
rect 24050 27806 24052 27858
rect 23996 27804 24052 27806
rect 24668 29426 24724 29428
rect 24668 29374 24670 29426
rect 24670 29374 24722 29426
rect 24722 29374 24724 29426
rect 24668 29372 24724 29374
rect 24108 28588 24164 28644
rect 24332 28812 24388 28868
rect 23548 26460 23604 26516
rect 24668 29202 24724 29204
rect 24668 29150 24670 29202
rect 24670 29150 24722 29202
rect 24722 29150 24724 29202
rect 24668 29148 24724 29150
rect 25228 36764 25284 36820
rect 25564 37212 25620 37268
rect 25900 36316 25956 36372
rect 25564 35922 25620 35924
rect 25564 35870 25566 35922
rect 25566 35870 25618 35922
rect 25618 35870 25620 35922
rect 25564 35868 25620 35870
rect 25228 35196 25284 35252
rect 26124 35698 26180 35700
rect 26124 35646 26126 35698
rect 26126 35646 26178 35698
rect 26178 35646 26180 35698
rect 26124 35644 26180 35646
rect 26012 35532 26068 35588
rect 25452 34354 25508 34356
rect 25452 34302 25454 34354
rect 25454 34302 25506 34354
rect 25506 34302 25508 34354
rect 25452 34300 25508 34302
rect 25340 34076 25396 34132
rect 26460 34130 26516 34132
rect 26460 34078 26462 34130
rect 26462 34078 26514 34130
rect 26514 34078 26516 34130
rect 26460 34076 26516 34078
rect 26012 33906 26068 33908
rect 26012 33854 26014 33906
rect 26014 33854 26066 33906
rect 26066 33854 26068 33906
rect 26012 33852 26068 33854
rect 26012 31666 26068 31668
rect 26012 31614 26014 31666
rect 26014 31614 26066 31666
rect 26066 31614 26068 31666
rect 26012 31612 26068 31614
rect 25676 31500 25732 31556
rect 25228 30380 25284 30436
rect 26124 31500 26180 31556
rect 26124 30268 26180 30324
rect 25340 29932 25396 29988
rect 25228 28812 25284 28868
rect 25452 29372 25508 29428
rect 25228 28642 25284 28644
rect 25228 28590 25230 28642
rect 25230 28590 25282 28642
rect 25282 28590 25284 28642
rect 25228 28588 25284 28590
rect 25452 28588 25508 28644
rect 23884 26178 23940 26180
rect 23884 26126 23886 26178
rect 23886 26126 23938 26178
rect 23938 26126 23940 26178
rect 23884 26124 23940 26126
rect 23548 25564 23604 25620
rect 23996 25506 24052 25508
rect 23996 25454 23998 25506
rect 23998 25454 24050 25506
rect 24050 25454 24052 25506
rect 23996 25452 24052 25454
rect 24332 26290 24388 26292
rect 24332 26238 24334 26290
rect 24334 26238 24386 26290
rect 24386 26238 24388 26290
rect 24332 26236 24388 26238
rect 24892 26012 24948 26068
rect 24444 25564 24500 25620
rect 24332 25340 24388 25396
rect 23100 24834 23156 24836
rect 23100 24782 23102 24834
rect 23102 24782 23154 24834
rect 23154 24782 23156 24834
rect 23100 24780 23156 24782
rect 21532 23826 21588 23828
rect 21532 23774 21534 23826
rect 21534 23774 21586 23826
rect 21586 23774 21588 23826
rect 21532 23772 21588 23774
rect 21868 23772 21924 23828
rect 21308 23436 21364 23492
rect 21196 23324 21252 23380
rect 21756 23324 21812 23380
rect 20412 22316 20468 22372
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19964 21698 20020 21700
rect 19964 21646 19966 21698
rect 19966 21646 20018 21698
rect 20018 21646 20020 21698
rect 19964 21644 20020 21646
rect 18620 20578 18676 20580
rect 18620 20526 18622 20578
rect 18622 20526 18674 20578
rect 18674 20526 18676 20578
rect 18620 20524 18676 20526
rect 20188 21586 20244 21588
rect 20188 21534 20190 21586
rect 20190 21534 20242 21586
rect 20242 21534 20244 21586
rect 20188 21532 20244 21534
rect 20524 21868 20580 21924
rect 21532 21868 21588 21924
rect 20860 21586 20916 21588
rect 20860 21534 20862 21586
rect 20862 21534 20914 21586
rect 20914 21534 20916 21586
rect 20860 21532 20916 21534
rect 19964 20636 20020 20692
rect 20300 20748 20356 20804
rect 19628 20412 19684 20468
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20188 20076 20244 20132
rect 19404 19794 19460 19796
rect 19404 19742 19406 19794
rect 19406 19742 19458 19794
rect 19458 19742 19460 19794
rect 19404 19740 19460 19742
rect 18732 15708 18788 15764
rect 18508 14476 18564 14532
rect 16604 13580 16660 13636
rect 16380 12460 16436 12516
rect 15372 11564 15428 11620
rect 15372 10668 15428 10724
rect 15484 11340 15540 11396
rect 15708 11452 15764 11508
rect 17164 13020 17220 13076
rect 17388 12460 17444 12516
rect 18284 13634 18340 13636
rect 18284 13582 18286 13634
rect 18286 13582 18338 13634
rect 18338 13582 18340 13634
rect 18284 13580 18340 13582
rect 18620 12684 18676 12740
rect 18396 12178 18452 12180
rect 18396 12126 18398 12178
rect 18398 12126 18450 12178
rect 18450 12126 18452 12178
rect 18396 12124 18452 12126
rect 16604 11452 16660 11508
rect 17276 11452 17332 11508
rect 15484 9324 15540 9380
rect 15036 6578 15092 6580
rect 15036 6526 15038 6578
rect 15038 6526 15090 6578
rect 15090 6526 15092 6578
rect 15036 6524 15092 6526
rect 15260 6524 15316 6580
rect 16380 9938 16436 9940
rect 16380 9886 16382 9938
rect 16382 9886 16434 9938
rect 16434 9886 16436 9938
rect 16380 9884 16436 9886
rect 16940 9938 16996 9940
rect 16940 9886 16942 9938
rect 16942 9886 16994 9938
rect 16994 9886 16996 9938
rect 16940 9884 16996 9886
rect 17836 11452 17892 11508
rect 21308 20690 21364 20692
rect 21308 20638 21310 20690
rect 21310 20638 21362 20690
rect 21362 20638 21364 20690
rect 21308 20636 21364 20638
rect 20860 20188 20916 20244
rect 21084 20188 21140 20244
rect 20300 19404 20356 19460
rect 20412 19740 20468 19796
rect 21308 20130 21364 20132
rect 21308 20078 21310 20130
rect 21310 20078 21362 20130
rect 21362 20078 21364 20130
rect 21308 20076 21364 20078
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 21084 19292 21140 19348
rect 21196 18620 21252 18676
rect 18956 16716 19012 16772
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19852 16492 19908 16548
rect 21308 18396 21364 18452
rect 21196 18226 21252 18228
rect 21196 18174 21198 18226
rect 21198 18174 21250 18226
rect 21250 18174 21252 18226
rect 21196 18172 21252 18174
rect 21644 21308 21700 21364
rect 21868 21532 21924 21588
rect 22204 23266 22260 23268
rect 22204 23214 22206 23266
rect 22206 23214 22258 23266
rect 22258 23214 22260 23266
rect 22204 23212 22260 23214
rect 22316 21868 22372 21924
rect 22092 21308 22148 21364
rect 23100 23938 23156 23940
rect 23100 23886 23102 23938
rect 23102 23886 23154 23938
rect 23154 23886 23156 23938
rect 23100 23884 23156 23886
rect 22764 23772 22820 23828
rect 22540 23100 22596 23156
rect 22652 23436 22708 23492
rect 22876 23714 22932 23716
rect 22876 23662 22878 23714
rect 22878 23662 22930 23714
rect 22930 23662 22932 23714
rect 22876 23660 22932 23662
rect 23100 23324 23156 23380
rect 23548 24834 23604 24836
rect 23548 24782 23550 24834
rect 23550 24782 23602 24834
rect 23602 24782 23604 24834
rect 23548 24780 23604 24782
rect 23660 24498 23716 24500
rect 23660 24446 23662 24498
rect 23662 24446 23714 24498
rect 23714 24446 23716 24498
rect 23660 24444 23716 24446
rect 23324 23324 23380 23380
rect 23100 22482 23156 22484
rect 23100 22430 23102 22482
rect 23102 22430 23154 22482
rect 23154 22430 23156 22482
rect 23100 22428 23156 22430
rect 23324 21868 23380 21924
rect 23212 21698 23268 21700
rect 23212 21646 23214 21698
rect 23214 21646 23266 21698
rect 23266 21646 23268 21698
rect 23212 21644 23268 21646
rect 22204 20188 22260 20244
rect 22764 20188 22820 20244
rect 21980 20076 22036 20132
rect 22428 20130 22484 20132
rect 22428 20078 22430 20130
rect 22430 20078 22482 20130
rect 22482 20078 22484 20130
rect 22428 20076 22484 20078
rect 21756 19964 21812 20020
rect 21644 19292 21700 19348
rect 20972 16268 21028 16324
rect 20636 16156 20692 16212
rect 18956 15932 19012 15988
rect 19180 15708 19236 15764
rect 20412 15986 20468 15988
rect 20412 15934 20414 15986
rect 20414 15934 20466 15986
rect 20466 15934 20468 15986
rect 20412 15932 20468 15934
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19180 15372 19236 15428
rect 19852 15314 19908 15316
rect 19852 15262 19854 15314
rect 19854 15262 19906 15314
rect 19906 15262 19908 15314
rect 19852 15260 19908 15262
rect 20524 15426 20580 15428
rect 20524 15374 20526 15426
rect 20526 15374 20578 15426
rect 20578 15374 20580 15426
rect 20524 15372 20580 15374
rect 20076 14588 20132 14644
rect 21644 18450 21700 18452
rect 21644 18398 21646 18450
rect 21646 18398 21698 18450
rect 21698 18398 21700 18450
rect 21644 18396 21700 18398
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19628 13580 19684 13636
rect 19404 12684 19460 12740
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19292 11900 19348 11956
rect 18956 10834 19012 10836
rect 18956 10782 18958 10834
rect 18958 10782 19010 10834
rect 19010 10782 19012 10834
rect 18956 10780 19012 10782
rect 19068 10220 19124 10276
rect 16268 8764 16324 8820
rect 18060 8764 18116 8820
rect 17836 8204 17892 8260
rect 17724 8146 17780 8148
rect 17724 8094 17726 8146
rect 17726 8094 17778 8146
rect 17778 8094 17780 8146
rect 17724 8092 17780 8094
rect 16828 7474 16884 7476
rect 16828 7422 16830 7474
rect 16830 7422 16882 7474
rect 16882 7422 16884 7474
rect 16828 7420 16884 7422
rect 17500 7474 17556 7476
rect 17500 7422 17502 7474
rect 17502 7422 17554 7474
rect 17554 7422 17556 7474
rect 17500 7420 17556 7422
rect 17836 7474 17892 7476
rect 17836 7422 17838 7474
rect 17838 7422 17890 7474
rect 17890 7422 17892 7474
rect 17836 7420 17892 7422
rect 15708 6690 15764 6692
rect 15708 6638 15710 6690
rect 15710 6638 15762 6690
rect 15762 6638 15764 6690
rect 15708 6636 15764 6638
rect 16604 6636 16660 6692
rect 16044 6018 16100 6020
rect 16044 5966 16046 6018
rect 16046 5966 16098 6018
rect 16098 5966 16100 6018
rect 16044 5964 16100 5966
rect 16492 5906 16548 5908
rect 16492 5854 16494 5906
rect 16494 5854 16546 5906
rect 16546 5854 16548 5906
rect 16492 5852 16548 5854
rect 17612 5906 17668 5908
rect 17612 5854 17614 5906
rect 17614 5854 17666 5906
rect 17666 5854 17668 5906
rect 17612 5852 17668 5854
rect 18732 8818 18788 8820
rect 18732 8766 18734 8818
rect 18734 8766 18786 8818
rect 18786 8766 18788 8818
rect 18732 8764 18788 8766
rect 18284 8258 18340 8260
rect 18284 8206 18286 8258
rect 18286 8206 18338 8258
rect 18338 8206 18340 8258
rect 18284 8204 18340 8206
rect 19292 8876 19348 8932
rect 19180 8258 19236 8260
rect 19180 8206 19182 8258
rect 19182 8206 19234 8258
rect 19234 8206 19236 8258
rect 19180 8204 19236 8206
rect 18508 7980 18564 8036
rect 19180 7980 19236 8036
rect 19180 7698 19236 7700
rect 19180 7646 19182 7698
rect 19182 7646 19234 7698
rect 19234 7646 19236 7698
rect 19180 7644 19236 7646
rect 18508 7586 18564 7588
rect 18508 7534 18510 7586
rect 18510 7534 18562 7586
rect 18562 7534 18564 7586
rect 18508 7532 18564 7534
rect 20076 11900 20132 11956
rect 20860 13132 20916 13188
rect 20524 12124 20580 12180
rect 21644 17276 21700 17332
rect 21532 16940 21588 16996
rect 21196 16492 21252 16548
rect 21420 16156 21476 16212
rect 21980 19906 22036 19908
rect 21980 19854 21982 19906
rect 21982 19854 22034 19906
rect 22034 19854 22036 19906
rect 21980 19852 22036 19854
rect 22652 19852 22708 19908
rect 22204 19516 22260 19572
rect 22092 19122 22148 19124
rect 22092 19070 22094 19122
rect 22094 19070 22146 19122
rect 22146 19070 22148 19122
rect 22092 19068 22148 19070
rect 21980 18060 22036 18116
rect 21980 17276 22036 17332
rect 21868 17052 21924 17108
rect 21644 15314 21700 15316
rect 21644 15262 21646 15314
rect 21646 15262 21698 15314
rect 21698 15262 21700 15314
rect 21644 15260 21700 15262
rect 21308 14476 21364 14532
rect 21420 13580 21476 13636
rect 21196 13468 21252 13524
rect 21980 15148 22036 15204
rect 22092 14642 22148 14644
rect 22092 14590 22094 14642
rect 22094 14590 22146 14642
rect 22146 14590 22148 14642
rect 22092 14588 22148 14590
rect 21868 13468 21924 13524
rect 21868 13244 21924 13300
rect 20748 11900 20804 11956
rect 20300 11788 20356 11844
rect 19964 11452 20020 11508
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19628 9772 19684 9828
rect 20076 10332 20132 10388
rect 20636 11282 20692 11284
rect 20636 11230 20638 11282
rect 20638 11230 20690 11282
rect 20690 11230 20692 11282
rect 20636 11228 20692 11230
rect 20300 10780 20356 10836
rect 20188 9996 20244 10052
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20412 9826 20468 9828
rect 20412 9774 20414 9826
rect 20414 9774 20466 9826
rect 20466 9774 20468 9826
rect 20412 9772 20468 9774
rect 21532 10332 21588 10388
rect 20076 8930 20132 8932
rect 20076 8878 20078 8930
rect 20078 8878 20130 8930
rect 20130 8878 20132 8930
rect 20076 8876 20132 8878
rect 20076 7980 20132 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19404 7420 19460 7476
rect 21308 8930 21364 8932
rect 21308 8878 21310 8930
rect 21310 8878 21362 8930
rect 21362 8878 21364 8930
rect 21308 8876 21364 8878
rect 20412 8764 20468 8820
rect 21756 8428 21812 8484
rect 22092 13186 22148 13188
rect 22092 13134 22094 13186
rect 22094 13134 22146 13186
rect 22146 13134 22148 13186
rect 22092 13132 22148 13134
rect 21980 12572 22036 12628
rect 22652 17052 22708 17108
rect 22764 16380 22820 16436
rect 23324 21084 23380 21140
rect 24220 23884 24276 23940
rect 24668 24946 24724 24948
rect 24668 24894 24670 24946
rect 24670 24894 24722 24946
rect 24722 24894 24724 24946
rect 24668 24892 24724 24894
rect 24444 23660 24500 23716
rect 23996 23436 24052 23492
rect 24556 24780 24612 24836
rect 23996 22540 24052 22596
rect 24444 22540 24500 22596
rect 24892 23938 24948 23940
rect 24892 23886 24894 23938
rect 24894 23886 24946 23938
rect 24946 23886 24948 23938
rect 24892 23884 24948 23886
rect 24556 21756 24612 21812
rect 24668 21698 24724 21700
rect 24668 21646 24670 21698
rect 24670 21646 24722 21698
rect 24722 21646 24724 21698
rect 24668 21644 24724 21646
rect 23436 20300 23492 20356
rect 23212 20242 23268 20244
rect 23212 20190 23214 20242
rect 23214 20190 23266 20242
rect 23266 20190 23268 20242
rect 23212 20188 23268 20190
rect 22988 19964 23044 20020
rect 23436 20018 23492 20020
rect 23436 19966 23438 20018
rect 23438 19966 23490 20018
rect 23490 19966 23492 20018
rect 23436 19964 23492 19966
rect 23212 17836 23268 17892
rect 23548 17554 23604 17556
rect 23548 17502 23550 17554
rect 23550 17502 23602 17554
rect 23602 17502 23604 17554
rect 23548 17500 23604 17502
rect 23772 20130 23828 20132
rect 23772 20078 23774 20130
rect 23774 20078 23826 20130
rect 23826 20078 23828 20130
rect 23772 20076 23828 20078
rect 24220 19346 24276 19348
rect 24220 19294 24222 19346
rect 24222 19294 24274 19346
rect 24274 19294 24276 19346
rect 24220 19292 24276 19294
rect 24220 18732 24276 18788
rect 24892 21532 24948 21588
rect 25116 26290 25172 26292
rect 25116 26238 25118 26290
rect 25118 26238 25170 26290
rect 25170 26238 25172 26290
rect 25116 26236 25172 26238
rect 27916 39618 27972 39620
rect 27916 39566 27918 39618
rect 27918 39566 27970 39618
rect 27970 39566 27972 39618
rect 27916 39564 27972 39566
rect 28476 43538 28532 43540
rect 28476 43486 28478 43538
rect 28478 43486 28530 43538
rect 28530 43486 28532 43538
rect 28476 43484 28532 43486
rect 28924 43538 28980 43540
rect 28924 43486 28926 43538
rect 28926 43486 28978 43538
rect 28978 43486 28980 43538
rect 28924 43484 28980 43486
rect 28700 43372 28756 43428
rect 28588 43148 28644 43204
rect 28476 42642 28532 42644
rect 28476 42590 28478 42642
rect 28478 42590 28530 42642
rect 28530 42590 28532 42642
rect 28476 42588 28532 42590
rect 28364 42364 28420 42420
rect 28364 42194 28420 42196
rect 28364 42142 28366 42194
rect 28366 42142 28418 42194
rect 28418 42142 28420 42194
rect 28364 42140 28420 42142
rect 28812 43314 28868 43316
rect 28812 43262 28814 43314
rect 28814 43262 28866 43314
rect 28866 43262 28868 43314
rect 28812 43260 28868 43262
rect 30716 45500 30772 45556
rect 30940 45052 30996 45108
rect 32396 46786 32452 46788
rect 32396 46734 32398 46786
rect 32398 46734 32450 46786
rect 32450 46734 32452 46786
rect 32396 46732 32452 46734
rect 32060 46620 32116 46676
rect 31724 46508 31780 46564
rect 31164 45724 31220 45780
rect 31276 45276 31332 45332
rect 31724 45778 31780 45780
rect 31724 45726 31726 45778
rect 31726 45726 31778 45778
rect 31778 45726 31780 45778
rect 31724 45724 31780 45726
rect 31388 45218 31444 45220
rect 31388 45166 31390 45218
rect 31390 45166 31442 45218
rect 31442 45166 31444 45218
rect 31388 45164 31444 45166
rect 31276 44492 31332 44548
rect 29932 44098 29988 44100
rect 29932 44046 29934 44098
rect 29934 44046 29986 44098
rect 29986 44046 29988 44098
rect 29932 44044 29988 44046
rect 30044 43932 30100 43988
rect 29708 43596 29764 43652
rect 29148 42866 29204 42868
rect 29148 42814 29150 42866
rect 29150 42814 29202 42866
rect 29202 42814 29204 42866
rect 29148 42812 29204 42814
rect 29484 42700 29540 42756
rect 29708 42812 29764 42868
rect 28588 41692 28644 41748
rect 30156 43820 30212 43876
rect 29932 42364 29988 42420
rect 28588 40908 28644 40964
rect 28364 40236 28420 40292
rect 29148 40348 29204 40404
rect 28252 39506 28308 39508
rect 28252 39454 28254 39506
rect 28254 39454 28306 39506
rect 28306 39454 28308 39506
rect 28252 39452 28308 39454
rect 27692 39004 27748 39060
rect 28924 40012 28980 40068
rect 29036 40124 29092 40180
rect 28588 39842 28644 39844
rect 28588 39790 28590 39842
rect 28590 39790 28642 39842
rect 28642 39790 28644 39842
rect 28588 39788 28644 39790
rect 28924 39788 28980 39844
rect 28588 39618 28644 39620
rect 28588 39566 28590 39618
rect 28590 39566 28642 39618
rect 28642 39566 28644 39618
rect 28588 39564 28644 39566
rect 29148 40012 29204 40068
rect 29036 39058 29092 39060
rect 29036 39006 29038 39058
rect 29038 39006 29090 39058
rect 29090 39006 29092 39058
rect 29036 39004 29092 39006
rect 27020 38274 27076 38276
rect 27020 38222 27022 38274
rect 27022 38222 27074 38274
rect 27074 38222 27076 38274
rect 27020 38220 27076 38222
rect 27916 38332 27972 38388
rect 27244 37266 27300 37268
rect 27244 37214 27246 37266
rect 27246 37214 27298 37266
rect 27298 37214 27300 37266
rect 27244 37212 27300 37214
rect 26908 36988 26964 37044
rect 27356 36540 27412 36596
rect 28476 38332 28532 38388
rect 28588 38050 28644 38052
rect 28588 37998 28590 38050
rect 28590 37998 28642 38050
rect 28642 37998 28644 38050
rect 28588 37996 28644 37998
rect 28028 36876 28084 36932
rect 27692 36370 27748 36372
rect 27692 36318 27694 36370
rect 27694 36318 27746 36370
rect 27746 36318 27748 36370
rect 27692 36316 27748 36318
rect 27020 34748 27076 34804
rect 27132 34636 27188 34692
rect 28140 36594 28196 36596
rect 28140 36542 28142 36594
rect 28142 36542 28194 36594
rect 28194 36542 28196 36594
rect 28140 36540 28196 36542
rect 28588 36594 28644 36596
rect 28588 36542 28590 36594
rect 28590 36542 28642 36594
rect 28642 36542 28644 36594
rect 28588 36540 28644 36542
rect 28812 35868 28868 35924
rect 29596 41858 29652 41860
rect 29596 41806 29598 41858
rect 29598 41806 29650 41858
rect 29650 41806 29652 41858
rect 29596 41804 29652 41806
rect 30044 41692 30100 41748
rect 30604 43708 30660 43764
rect 30268 43484 30324 43540
rect 30268 41580 30324 41636
rect 30380 41916 30436 41972
rect 29484 41074 29540 41076
rect 29484 41022 29486 41074
rect 29486 41022 29538 41074
rect 29538 41022 29540 41074
rect 29484 41020 29540 41022
rect 29372 40402 29428 40404
rect 29372 40350 29374 40402
rect 29374 40350 29426 40402
rect 29426 40350 29428 40402
rect 29372 40348 29428 40350
rect 30268 40962 30324 40964
rect 30268 40910 30270 40962
rect 30270 40910 30322 40962
rect 30322 40910 30324 40962
rect 30268 40908 30324 40910
rect 29596 40236 29652 40292
rect 29820 40290 29876 40292
rect 29820 40238 29822 40290
rect 29822 40238 29874 40290
rect 29874 40238 29876 40290
rect 29820 40236 29876 40238
rect 29708 39394 29764 39396
rect 29708 39342 29710 39394
rect 29710 39342 29762 39394
rect 29762 39342 29764 39394
rect 29708 39340 29764 39342
rect 30156 39004 30212 39060
rect 30604 41580 30660 41636
rect 31052 44098 31108 44100
rect 31052 44046 31054 44098
rect 31054 44046 31106 44098
rect 31106 44046 31108 44098
rect 31052 44044 31108 44046
rect 31276 44322 31332 44324
rect 31276 44270 31278 44322
rect 31278 44270 31330 44322
rect 31330 44270 31332 44322
rect 31276 44268 31332 44270
rect 31612 44604 31668 44660
rect 32284 45218 32340 45220
rect 32284 45166 32286 45218
rect 32286 45166 32338 45218
rect 32338 45166 32340 45218
rect 32284 45164 32340 45166
rect 33068 46956 33124 47012
rect 31164 43148 31220 43204
rect 32508 44604 32564 44660
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 34748 48914 34804 48916
rect 34748 48862 34750 48914
rect 34750 48862 34802 48914
rect 34802 48862 34804 48914
rect 34748 48860 34804 48862
rect 34972 48914 35028 48916
rect 34972 48862 34974 48914
rect 34974 48862 35026 48914
rect 35026 48862 35028 48914
rect 34972 48860 35028 48862
rect 34076 48300 34132 48356
rect 33404 46172 33460 46228
rect 33628 47068 33684 47124
rect 33292 45724 33348 45780
rect 32956 44492 33012 44548
rect 33404 44828 33460 44884
rect 32844 44434 32900 44436
rect 32844 44382 32846 44434
rect 32846 44382 32898 44434
rect 32898 44382 32900 44434
rect 32844 44380 32900 44382
rect 32172 43708 32228 43764
rect 32396 44268 32452 44324
rect 31388 42364 31444 42420
rect 31276 42194 31332 42196
rect 31276 42142 31278 42194
rect 31278 42142 31330 42194
rect 31330 42142 31332 42194
rect 31276 42140 31332 42142
rect 30828 42028 30884 42084
rect 30940 41970 30996 41972
rect 30940 41918 30942 41970
rect 30942 41918 30994 41970
rect 30994 41918 30996 41970
rect 30940 41916 30996 41918
rect 30828 41356 30884 41412
rect 30604 40348 30660 40404
rect 32284 42194 32340 42196
rect 32284 42142 32286 42194
rect 32286 42142 32338 42194
rect 32338 42142 32340 42194
rect 32284 42140 32340 42142
rect 32060 42082 32116 42084
rect 32060 42030 32062 42082
rect 32062 42030 32114 42082
rect 32114 42030 32116 42082
rect 32060 42028 32116 42030
rect 31948 41916 32004 41972
rect 32172 41692 32228 41748
rect 31948 41468 32004 41524
rect 31836 41356 31892 41412
rect 32060 41244 32116 41300
rect 32284 40626 32340 40628
rect 32284 40574 32286 40626
rect 32286 40574 32338 40626
rect 32338 40574 32340 40626
rect 32284 40572 32340 40574
rect 31948 39788 32004 39844
rect 33404 44268 33460 44324
rect 33516 44492 33572 44548
rect 33404 44044 33460 44100
rect 32620 42028 32676 42084
rect 33068 41916 33124 41972
rect 33292 41916 33348 41972
rect 33068 41746 33124 41748
rect 33068 41694 33070 41746
rect 33070 41694 33122 41746
rect 33122 41694 33124 41746
rect 33068 41692 33124 41694
rect 33516 41916 33572 41972
rect 33516 41132 33572 41188
rect 32508 40236 32564 40292
rect 30828 38722 30884 38724
rect 30828 38670 30830 38722
rect 30830 38670 30882 38722
rect 30882 38670 30884 38722
rect 30828 38668 30884 38670
rect 29484 38050 29540 38052
rect 29484 37998 29486 38050
rect 29486 37998 29538 38050
rect 29538 37998 29540 38050
rect 29484 37996 29540 37998
rect 29484 36540 29540 36596
rect 29260 35922 29316 35924
rect 29260 35870 29262 35922
rect 29262 35870 29314 35922
rect 29314 35870 29316 35922
rect 29260 35868 29316 35870
rect 27916 35586 27972 35588
rect 27916 35534 27918 35586
rect 27918 35534 27970 35586
rect 27970 35534 27972 35586
rect 27916 35532 27972 35534
rect 30268 38050 30324 38052
rect 30268 37998 30270 38050
rect 30270 37998 30322 38050
rect 30322 37998 30324 38050
rect 30268 37996 30324 37998
rect 29820 37938 29876 37940
rect 29820 37886 29822 37938
rect 29822 37886 29874 37938
rect 29874 37886 29876 37938
rect 29820 37884 29876 37886
rect 30492 37266 30548 37268
rect 30492 37214 30494 37266
rect 30494 37214 30546 37266
rect 30546 37214 30548 37266
rect 30492 37212 30548 37214
rect 30044 37154 30100 37156
rect 30044 37102 30046 37154
rect 30046 37102 30098 37154
rect 30098 37102 30100 37154
rect 30044 37100 30100 37102
rect 30044 36594 30100 36596
rect 30044 36542 30046 36594
rect 30046 36542 30098 36594
rect 30098 36542 30100 36594
rect 30044 36540 30100 36542
rect 30268 35922 30324 35924
rect 30268 35870 30270 35922
rect 30270 35870 30322 35922
rect 30322 35870 30324 35922
rect 30268 35868 30324 35870
rect 31948 38668 32004 38724
rect 30716 37938 30772 37940
rect 30716 37886 30718 37938
rect 30718 37886 30770 37938
rect 30770 37886 30772 37938
rect 30716 37884 30772 37886
rect 33292 38220 33348 38276
rect 33404 39228 33460 39284
rect 30940 37154 30996 37156
rect 30940 37102 30942 37154
rect 30942 37102 30994 37154
rect 30994 37102 30996 37154
rect 30940 37100 30996 37102
rect 30828 35980 30884 36036
rect 30492 35810 30548 35812
rect 30492 35758 30494 35810
rect 30494 35758 30546 35810
rect 30546 35758 30548 35810
rect 30492 35756 30548 35758
rect 29148 34914 29204 34916
rect 29148 34862 29150 34914
rect 29150 34862 29202 34914
rect 29202 34862 29204 34914
rect 29148 34860 29204 34862
rect 29260 34972 29316 35028
rect 27468 34300 27524 34356
rect 29484 34860 29540 34916
rect 29372 34690 29428 34692
rect 29372 34638 29374 34690
rect 29374 34638 29426 34690
rect 29426 34638 29428 34690
rect 29372 34636 29428 34638
rect 27132 33852 27188 33908
rect 26684 31836 26740 31892
rect 26684 30828 26740 30884
rect 26572 30210 26628 30212
rect 26572 30158 26574 30210
rect 26574 30158 26626 30210
rect 26626 30158 26628 30210
rect 26572 30156 26628 30158
rect 26908 30268 26964 30324
rect 26460 28812 26516 28868
rect 26684 29708 26740 29764
rect 26236 27804 26292 27860
rect 30268 34914 30324 34916
rect 30268 34862 30270 34914
rect 30270 34862 30322 34914
rect 30322 34862 30324 34914
rect 30268 34860 30324 34862
rect 29596 34130 29652 34132
rect 29596 34078 29598 34130
rect 29598 34078 29650 34130
rect 29650 34078 29652 34130
rect 29596 34076 29652 34078
rect 30380 33458 30436 33460
rect 30380 33406 30382 33458
rect 30382 33406 30434 33458
rect 30434 33406 30436 33458
rect 30380 33404 30436 33406
rect 27244 32450 27300 32452
rect 27244 32398 27246 32450
rect 27246 32398 27298 32450
rect 27298 32398 27300 32450
rect 27244 32396 27300 32398
rect 30044 33180 30100 33236
rect 29708 32732 29764 32788
rect 29148 32396 29204 32452
rect 27356 31890 27412 31892
rect 27356 31838 27358 31890
rect 27358 31838 27410 31890
rect 27410 31838 27412 31890
rect 27356 31836 27412 31838
rect 28252 31724 28308 31780
rect 28028 31164 28084 31220
rect 27356 30882 27412 30884
rect 27356 30830 27358 30882
rect 27358 30830 27410 30882
rect 27410 30830 27412 30882
rect 27356 30828 27412 30830
rect 27132 30380 27188 30436
rect 27020 29708 27076 29764
rect 25340 26178 25396 26180
rect 25340 26126 25342 26178
rect 25342 26126 25394 26178
rect 25394 26126 25396 26178
rect 25340 26124 25396 26126
rect 25340 25340 25396 25396
rect 25116 25228 25172 25284
rect 25452 24780 25508 24836
rect 26124 26066 26180 26068
rect 26124 26014 26126 26066
rect 26126 26014 26178 26066
rect 26178 26014 26180 26066
rect 26124 26012 26180 26014
rect 25564 25452 25620 25508
rect 25676 25228 25732 25284
rect 25340 23996 25396 24052
rect 25228 23884 25284 23940
rect 25340 23324 25396 23380
rect 26124 25116 26180 25172
rect 25788 24444 25844 24500
rect 25676 23042 25732 23044
rect 25676 22990 25678 23042
rect 25678 22990 25730 23042
rect 25730 22990 25732 23042
rect 25676 22988 25732 22990
rect 25452 21586 25508 21588
rect 25452 21534 25454 21586
rect 25454 21534 25506 21586
rect 25506 21534 25508 21586
rect 25452 21532 25508 21534
rect 25116 21420 25172 21476
rect 25452 21308 25508 21364
rect 24556 20802 24612 20804
rect 24556 20750 24558 20802
rect 24558 20750 24610 20802
rect 24610 20750 24612 20802
rect 24556 20748 24612 20750
rect 24668 19906 24724 19908
rect 24668 19854 24670 19906
rect 24670 19854 24722 19906
rect 24722 19854 24724 19906
rect 24668 19852 24724 19854
rect 25004 19234 25060 19236
rect 25004 19182 25006 19234
rect 25006 19182 25058 19234
rect 25058 19182 25060 19234
rect 25004 19180 25060 19182
rect 26348 24946 26404 24948
rect 26348 24894 26350 24946
rect 26350 24894 26402 24946
rect 26402 24894 26404 24946
rect 26348 24892 26404 24894
rect 25788 21362 25844 21364
rect 25788 21310 25790 21362
rect 25790 21310 25842 21362
rect 25842 21310 25844 21362
rect 25788 21308 25844 21310
rect 25564 19852 25620 19908
rect 25676 20188 25732 20244
rect 25228 19068 25284 19124
rect 23436 16380 23492 16436
rect 23100 15148 23156 15204
rect 23324 15596 23380 15652
rect 22876 14588 22932 14644
rect 22316 13634 22372 13636
rect 22316 13582 22318 13634
rect 22318 13582 22370 13634
rect 22370 13582 22372 13634
rect 22316 13580 22372 13582
rect 22316 13132 22372 13188
rect 22764 12962 22820 12964
rect 22764 12910 22766 12962
rect 22766 12910 22818 12962
rect 22818 12910 22820 12962
rect 22764 12908 22820 12910
rect 23436 13804 23492 13860
rect 24668 18338 24724 18340
rect 24668 18286 24670 18338
rect 24670 18286 24722 18338
rect 24722 18286 24724 18338
rect 24668 18284 24724 18286
rect 23884 17836 23940 17892
rect 24668 17276 24724 17332
rect 23772 17164 23828 17220
rect 24332 17164 24388 17220
rect 23884 16994 23940 16996
rect 23884 16942 23886 16994
rect 23886 16942 23938 16994
rect 23938 16942 23940 16994
rect 23884 16940 23940 16942
rect 23660 16716 23716 16772
rect 24220 16604 24276 16660
rect 23660 15538 23716 15540
rect 23660 15486 23662 15538
rect 23662 15486 23714 15538
rect 23714 15486 23716 15538
rect 23660 15484 23716 15486
rect 23772 16044 23828 16100
rect 25228 18396 25284 18452
rect 24892 18172 24948 18228
rect 25452 19346 25508 19348
rect 25452 19294 25454 19346
rect 25454 19294 25506 19346
rect 25506 19294 25508 19346
rect 25452 19292 25508 19294
rect 25676 19122 25732 19124
rect 25676 19070 25678 19122
rect 25678 19070 25730 19122
rect 25730 19070 25732 19122
rect 25676 19068 25732 19070
rect 25676 18844 25732 18900
rect 25452 18172 25508 18228
rect 25564 17836 25620 17892
rect 24668 16940 24724 16996
rect 24556 16828 24612 16884
rect 24220 15932 24276 15988
rect 23548 13244 23604 13300
rect 22988 12796 23044 12852
rect 23436 12402 23492 12404
rect 23436 12350 23438 12402
rect 23438 12350 23490 12402
rect 23490 12350 23492 12402
rect 23436 12348 23492 12350
rect 22092 11676 22148 11732
rect 23436 11506 23492 11508
rect 23436 11454 23438 11506
rect 23438 11454 23490 11506
rect 23490 11454 23492 11506
rect 23436 11452 23492 11454
rect 22876 11228 22932 11284
rect 23324 9996 23380 10052
rect 22316 9826 22372 9828
rect 22316 9774 22318 9826
rect 22318 9774 22370 9826
rect 22370 9774 22372 9826
rect 22316 9772 22372 9774
rect 21980 8764 22036 8820
rect 21868 7644 21924 7700
rect 18956 6690 19012 6692
rect 18956 6638 18958 6690
rect 18958 6638 19010 6690
rect 19010 6638 19012 6690
rect 18956 6636 19012 6638
rect 19628 6636 19684 6692
rect 18508 6018 18564 6020
rect 18508 5966 18510 6018
rect 18510 5966 18562 6018
rect 18562 5966 18564 6018
rect 18508 5964 18564 5966
rect 19404 5964 19460 6020
rect 21868 6748 21924 6804
rect 20300 6636 20356 6692
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 22316 8876 22372 8932
rect 22876 8146 22932 8148
rect 22876 8094 22878 8146
rect 22878 8094 22930 8146
rect 22930 8094 22932 8146
rect 22876 8092 22932 8094
rect 22316 7756 22372 7812
rect 25004 16380 25060 16436
rect 25116 17388 25172 17444
rect 25228 17164 25284 17220
rect 25228 16882 25284 16884
rect 25228 16830 25230 16882
rect 25230 16830 25282 16882
rect 25282 16830 25284 16882
rect 25228 16828 25284 16830
rect 26460 22988 26516 23044
rect 26460 22316 26516 22372
rect 26684 25564 26740 25620
rect 26684 24834 26740 24836
rect 26684 24782 26686 24834
rect 26686 24782 26738 24834
rect 26738 24782 26740 24834
rect 26684 24780 26740 24782
rect 26796 23996 26852 24052
rect 26684 21868 26740 21924
rect 26572 21756 26628 21812
rect 26572 21420 26628 21476
rect 28140 30156 28196 30212
rect 29596 31948 29652 32004
rect 29260 30940 29316 30996
rect 29484 30716 29540 30772
rect 28476 30098 28532 30100
rect 28476 30046 28478 30098
rect 28478 30046 28530 30098
rect 28530 30046 28532 30098
rect 28476 30044 28532 30046
rect 27580 29148 27636 29204
rect 28252 29596 28308 29652
rect 27804 28812 27860 28868
rect 27356 28642 27412 28644
rect 27356 28590 27358 28642
rect 27358 28590 27410 28642
rect 27410 28590 27412 28642
rect 27356 28588 27412 28590
rect 31164 37884 31220 37940
rect 31500 37490 31556 37492
rect 31500 37438 31502 37490
rect 31502 37438 31554 37490
rect 31554 37438 31556 37490
rect 31500 37436 31556 37438
rect 31724 37212 31780 37268
rect 32060 37154 32116 37156
rect 32060 37102 32062 37154
rect 32062 37102 32114 37154
rect 32114 37102 32116 37154
rect 32060 37100 32116 37102
rect 31836 36258 31892 36260
rect 31836 36206 31838 36258
rect 31838 36206 31890 36258
rect 31890 36206 31892 36258
rect 31836 36204 31892 36206
rect 31276 35084 31332 35140
rect 33068 37266 33124 37268
rect 33068 37214 33070 37266
rect 33070 37214 33122 37266
rect 33122 37214 33124 37266
rect 33068 37212 33124 37214
rect 33404 36876 33460 36932
rect 32508 36428 32564 36484
rect 33516 36428 33572 36484
rect 32396 36204 32452 36260
rect 32172 35980 32228 36036
rect 33180 34802 33236 34804
rect 33180 34750 33182 34802
rect 33182 34750 33234 34802
rect 33234 34750 33236 34802
rect 33180 34748 33236 34750
rect 32508 33852 32564 33908
rect 32732 33458 32788 33460
rect 32732 33406 32734 33458
rect 32734 33406 32786 33458
rect 32786 33406 32788 33458
rect 32732 33404 32788 33406
rect 33516 34076 33572 34132
rect 33964 46674 34020 46676
rect 33964 46622 33966 46674
rect 33966 46622 34018 46674
rect 34018 46622 34020 46674
rect 33964 46620 34020 46622
rect 33740 44828 33796 44884
rect 33740 44380 33796 44436
rect 34412 46956 34468 47012
rect 35420 48802 35476 48804
rect 35420 48750 35422 48802
rect 35422 48750 35474 48802
rect 35474 48750 35476 48802
rect 35420 48748 35476 48750
rect 35980 51602 36036 51604
rect 35980 51550 35982 51602
rect 35982 51550 36034 51602
rect 36034 51550 36036 51602
rect 35980 51548 36036 51550
rect 35980 51324 36036 51380
rect 35868 51154 35924 51156
rect 35868 51102 35870 51154
rect 35870 51102 35922 51154
rect 35922 51102 35924 51154
rect 35868 51100 35924 51102
rect 37660 52220 37716 52276
rect 36428 50316 36484 50372
rect 36204 49810 36260 49812
rect 36204 49758 36206 49810
rect 36206 49758 36258 49810
rect 36258 49758 36260 49810
rect 36204 49756 36260 49758
rect 37100 51436 37156 51492
rect 36988 50988 37044 51044
rect 36988 50594 37044 50596
rect 36988 50542 36990 50594
rect 36990 50542 37042 50594
rect 37042 50542 37044 50594
rect 36988 50540 37044 50542
rect 37212 50764 37268 50820
rect 36652 50316 36708 50372
rect 36876 50204 36932 50260
rect 36652 49532 36708 49588
rect 36764 50092 36820 50148
rect 36204 49026 36260 49028
rect 36204 48974 36206 49026
rect 36206 48974 36258 49026
rect 36258 48974 36260 49026
rect 36204 48972 36260 48974
rect 38108 53506 38164 53508
rect 38108 53454 38110 53506
rect 38110 53454 38162 53506
rect 38162 53454 38164 53506
rect 38108 53452 38164 53454
rect 38108 53004 38164 53060
rect 37996 52386 38052 52388
rect 37996 52334 37998 52386
rect 37998 52334 38050 52386
rect 38050 52334 38052 52386
rect 37996 52332 38052 52334
rect 38220 52780 38276 52836
rect 37884 51548 37940 51604
rect 37996 51938 38052 51940
rect 37996 51886 37998 51938
rect 37998 51886 38050 51938
rect 38050 51886 38052 51938
rect 37996 51884 38052 51886
rect 37772 51324 37828 51380
rect 37324 50204 37380 50260
rect 37100 49868 37156 49924
rect 36428 48860 36484 48916
rect 36876 49196 36932 49252
rect 36092 48802 36148 48804
rect 36092 48750 36094 48802
rect 36094 48750 36146 48802
rect 36146 48750 36148 48802
rect 36092 48748 36148 48750
rect 36204 48242 36260 48244
rect 36204 48190 36206 48242
rect 36206 48190 36258 48242
rect 36258 48190 36260 48242
rect 36204 48188 36260 48190
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 34748 46956 34804 47012
rect 34412 46620 34468 46676
rect 33964 45106 34020 45108
rect 33964 45054 33966 45106
rect 33966 45054 34018 45106
rect 34018 45054 34020 45106
rect 33964 45052 34020 45054
rect 35756 46956 35812 47012
rect 36316 46956 36372 47012
rect 35980 46450 36036 46452
rect 35980 46398 35982 46450
rect 35982 46398 36034 46450
rect 36034 46398 36036 46450
rect 35980 46396 36036 46398
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 34188 44994 34244 44996
rect 34188 44942 34190 44994
rect 34190 44942 34242 44994
rect 34242 44942 34244 44994
rect 34188 44940 34244 44942
rect 33964 44210 34020 44212
rect 33964 44158 33966 44210
rect 33966 44158 34018 44210
rect 34018 44158 34020 44210
rect 33964 44156 34020 44158
rect 34076 44098 34132 44100
rect 34076 44046 34078 44098
rect 34078 44046 34130 44098
rect 34130 44046 34132 44098
rect 34076 44044 34132 44046
rect 34188 42252 34244 42308
rect 34188 40124 34244 40180
rect 33740 39340 33796 39396
rect 33964 37660 34020 37716
rect 34636 44098 34692 44100
rect 34636 44046 34638 44098
rect 34638 44046 34690 44098
rect 34690 44046 34692 44098
rect 34636 44044 34692 44046
rect 34524 43932 34580 43988
rect 34524 43260 34580 43316
rect 35420 44994 35476 44996
rect 35420 44942 35422 44994
rect 35422 44942 35474 44994
rect 35474 44942 35476 44994
rect 35420 44940 35476 44942
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34748 43426 34804 43428
rect 34748 43374 34750 43426
rect 34750 43374 34802 43426
rect 34802 43374 34804 43426
rect 34748 43372 34804 43374
rect 35868 43426 35924 43428
rect 35868 43374 35870 43426
rect 35870 43374 35922 43426
rect 35922 43374 35924 43426
rect 35868 43372 35924 43374
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34748 42754 34804 42756
rect 34748 42702 34750 42754
rect 34750 42702 34802 42754
rect 34802 42702 34804 42754
rect 34748 42700 34804 42702
rect 34972 42530 35028 42532
rect 34972 42478 34974 42530
rect 34974 42478 35026 42530
rect 35026 42478 35028 42530
rect 34972 42476 35028 42478
rect 34748 42028 34804 42084
rect 34860 41356 34916 41412
rect 34636 41132 34692 41188
rect 35644 42252 35700 42308
rect 35196 42140 35252 42196
rect 35532 42082 35588 42084
rect 35532 42030 35534 42082
rect 35534 42030 35586 42082
rect 35586 42030 35588 42082
rect 35532 42028 35588 42030
rect 35084 41916 35140 41972
rect 35868 41970 35924 41972
rect 35868 41918 35870 41970
rect 35870 41918 35922 41970
rect 35922 41918 35924 41970
rect 35868 41916 35924 41918
rect 35308 41692 35364 41748
rect 35756 41804 35812 41860
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 34972 41020 35028 41076
rect 35084 41244 35140 41300
rect 35420 40124 35476 40180
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 37100 49026 37156 49028
rect 37100 48974 37102 49026
rect 37102 48974 37154 49026
rect 37154 48974 37156 49026
rect 37100 48972 37156 48974
rect 37548 49756 37604 49812
rect 38108 51660 38164 51716
rect 38220 51996 38276 52052
rect 38220 51436 38276 51492
rect 38668 53730 38724 53732
rect 38668 53678 38670 53730
rect 38670 53678 38722 53730
rect 38722 53678 38724 53730
rect 38668 53676 38724 53678
rect 38444 53340 38500 53396
rect 38444 52668 38500 52724
rect 38892 53676 38948 53732
rect 38668 53228 38724 53284
rect 39116 53730 39172 53732
rect 39116 53678 39118 53730
rect 39118 53678 39170 53730
rect 39170 53678 39172 53730
rect 39116 53676 39172 53678
rect 41020 57036 41076 57092
rect 40460 56700 40516 56756
rect 42140 56924 42196 56980
rect 42924 57036 42980 57092
rect 41692 56252 41748 56308
rect 42028 56812 42084 56868
rect 41804 55186 41860 55188
rect 41804 55134 41806 55186
rect 41806 55134 41858 55186
rect 41858 55134 41860 55186
rect 41804 55132 41860 55134
rect 39452 54236 39508 54292
rect 39564 53842 39620 53844
rect 39564 53790 39566 53842
rect 39566 53790 39618 53842
rect 39618 53790 39620 53842
rect 39564 53788 39620 53790
rect 39340 53676 39396 53732
rect 39452 53618 39508 53620
rect 39452 53566 39454 53618
rect 39454 53566 39506 53618
rect 39506 53566 39508 53618
rect 39452 53564 39508 53566
rect 41804 53676 41860 53732
rect 38444 52274 38500 52276
rect 38444 52222 38446 52274
rect 38446 52222 38498 52274
rect 38498 52222 38500 52274
rect 38444 52220 38500 52222
rect 38892 52780 38948 52836
rect 38892 52332 38948 52388
rect 38780 52050 38836 52052
rect 38780 51998 38782 52050
rect 38782 51998 38834 52050
rect 38834 51998 38836 52050
rect 38780 51996 38836 51998
rect 38780 51772 38836 51828
rect 38556 51602 38612 51604
rect 38556 51550 38558 51602
rect 38558 51550 38610 51602
rect 38610 51550 38612 51602
rect 38556 51548 38612 51550
rect 38444 51490 38500 51492
rect 38444 51438 38446 51490
rect 38446 51438 38498 51490
rect 38498 51438 38500 51490
rect 38444 51436 38500 51438
rect 38332 50764 38388 50820
rect 38220 50652 38276 50708
rect 38220 50428 38276 50484
rect 38444 50428 38500 50484
rect 38668 50428 38724 50484
rect 37996 50092 38052 50148
rect 38668 49980 38724 50036
rect 37436 49026 37492 49028
rect 37436 48974 37438 49026
rect 37438 48974 37490 49026
rect 37490 48974 37492 49026
rect 37436 48972 37492 48974
rect 37660 48914 37716 48916
rect 37660 48862 37662 48914
rect 37662 48862 37714 48914
rect 37714 48862 37716 48914
rect 37660 48860 37716 48862
rect 39004 51212 39060 51268
rect 38892 51100 38948 51156
rect 39228 53116 39284 53172
rect 39340 53452 39396 53508
rect 39228 52668 39284 52724
rect 39564 53452 39620 53508
rect 39900 53452 39956 53508
rect 39788 53340 39844 53396
rect 40908 53228 40964 53284
rect 40236 53116 40292 53172
rect 39788 52892 39844 52948
rect 39676 52834 39732 52836
rect 39676 52782 39678 52834
rect 39678 52782 39730 52834
rect 39730 52782 39732 52834
rect 39676 52780 39732 52782
rect 39452 52162 39508 52164
rect 39452 52110 39454 52162
rect 39454 52110 39506 52162
rect 39506 52110 39508 52162
rect 39452 52108 39508 52110
rect 40012 52108 40068 52164
rect 41132 52946 41188 52948
rect 41132 52894 41134 52946
rect 41134 52894 41186 52946
rect 41186 52894 41188 52946
rect 41132 52892 41188 52894
rect 41020 52722 41076 52724
rect 41020 52670 41022 52722
rect 41022 52670 41074 52722
rect 41074 52670 41076 52722
rect 41020 52668 41076 52670
rect 42252 53730 42308 53732
rect 42252 53678 42254 53730
rect 42254 53678 42306 53730
rect 42306 53678 42308 53730
rect 42252 53676 42308 53678
rect 42924 55186 42980 55188
rect 42924 55134 42926 55186
rect 42926 55134 42978 55186
rect 42978 55134 42980 55186
rect 42924 55132 42980 55134
rect 44044 56924 44100 56980
rect 43596 56306 43652 56308
rect 43596 56254 43598 56306
rect 43598 56254 43650 56306
rect 43650 56254 43652 56306
rect 43596 56252 43652 56254
rect 43484 55916 43540 55972
rect 44492 55970 44548 55972
rect 44492 55918 44494 55970
rect 44494 55918 44546 55970
rect 44546 55918 44548 55970
rect 44492 55916 44548 55918
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 44828 55804 44884 55860
rect 45388 55858 45444 55860
rect 45388 55806 45390 55858
rect 45390 55806 45442 55858
rect 45442 55806 45444 55858
rect 45388 55804 45444 55806
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 43036 54236 43092 54292
rect 43708 54236 43764 54292
rect 42588 53676 42644 53732
rect 42140 53170 42196 53172
rect 42140 53118 42142 53170
rect 42142 53118 42194 53170
rect 42194 53118 42196 53170
rect 42140 53116 42196 53118
rect 42588 53170 42644 53172
rect 42588 53118 42590 53170
rect 42590 53118 42642 53170
rect 42642 53118 42644 53170
rect 42588 53116 42644 53118
rect 40796 52386 40852 52388
rect 40796 52334 40798 52386
rect 40798 52334 40850 52386
rect 40850 52334 40852 52386
rect 40796 52332 40852 52334
rect 39452 51884 39508 51940
rect 40124 51772 40180 51828
rect 39676 51266 39732 51268
rect 39676 51214 39678 51266
rect 39678 51214 39730 51266
rect 39730 51214 39732 51266
rect 39676 51212 39732 51214
rect 39004 50764 39060 50820
rect 39228 50706 39284 50708
rect 39228 50654 39230 50706
rect 39230 50654 39282 50706
rect 39282 50654 39284 50706
rect 39228 50652 39284 50654
rect 39452 50652 39508 50708
rect 39116 50594 39172 50596
rect 39116 50542 39118 50594
rect 39118 50542 39170 50594
rect 39170 50542 39172 50594
rect 39116 50540 39172 50542
rect 39228 50428 39284 50484
rect 41916 52892 41972 52948
rect 41804 52274 41860 52276
rect 41804 52222 41806 52274
rect 41806 52222 41858 52274
rect 41858 52222 41860 52274
rect 41804 52220 41860 52222
rect 41580 52050 41636 52052
rect 41580 51998 41582 52050
rect 41582 51998 41634 52050
rect 41634 51998 41636 52050
rect 41580 51996 41636 51998
rect 41916 51660 41972 51716
rect 41244 51100 41300 51156
rect 41692 50876 41748 50932
rect 41580 50652 41636 50708
rect 40908 50540 40964 50596
rect 40236 50428 40292 50484
rect 39116 50092 39172 50148
rect 39116 49756 39172 49812
rect 40012 50370 40068 50372
rect 40012 50318 40014 50370
rect 40014 50318 40066 50370
rect 40066 50318 40068 50370
rect 40012 50316 40068 50318
rect 40012 49980 40068 50036
rect 39900 49756 39956 49812
rect 39788 49196 39844 49252
rect 39116 49026 39172 49028
rect 39116 48974 39118 49026
rect 39118 48974 39170 49026
rect 39170 48974 39172 49026
rect 39116 48972 39172 48974
rect 39788 49026 39844 49028
rect 39788 48974 39790 49026
rect 39790 48974 39842 49026
rect 39842 48974 39844 49026
rect 39788 48972 39844 48974
rect 38332 48860 38388 48916
rect 39452 48914 39508 48916
rect 39452 48862 39454 48914
rect 39454 48862 39506 48914
rect 39506 48862 39508 48914
rect 39452 48860 39508 48862
rect 41356 49980 41412 50036
rect 40684 49644 40740 49700
rect 41244 49644 41300 49700
rect 41356 49532 41412 49588
rect 39900 48860 39956 48916
rect 42028 52162 42084 52164
rect 42028 52110 42030 52162
rect 42030 52110 42082 52162
rect 42082 52110 42084 52162
rect 42028 52108 42084 52110
rect 42140 51772 42196 51828
rect 42252 51100 42308 51156
rect 42364 50876 42420 50932
rect 41916 50540 41972 50596
rect 42140 50540 42196 50596
rect 42028 49756 42084 49812
rect 42700 52050 42756 52052
rect 42700 51998 42702 52050
rect 42702 51998 42754 52050
rect 42754 51998 42756 52050
rect 42700 51996 42756 51998
rect 44828 54236 44884 54292
rect 45052 53676 45108 53732
rect 42812 51772 42868 51828
rect 43932 52946 43988 52948
rect 43932 52894 43934 52946
rect 43934 52894 43986 52946
rect 43986 52894 43988 52946
rect 43932 52892 43988 52894
rect 43484 51772 43540 51828
rect 43820 51884 43876 51940
rect 42700 50540 42756 50596
rect 42924 50652 42980 50708
rect 43708 51324 43764 51380
rect 42924 50482 42980 50484
rect 42924 50430 42926 50482
rect 42926 50430 42978 50482
rect 42978 50430 42980 50482
rect 42924 50428 42980 50430
rect 42364 50316 42420 50372
rect 41804 49196 41860 49252
rect 43372 51100 43428 51156
rect 43596 50764 43652 50820
rect 43036 50092 43092 50148
rect 45500 53676 45556 53732
rect 46956 53676 47012 53732
rect 46284 53618 46340 53620
rect 46284 53566 46286 53618
rect 46286 53566 46338 53618
rect 46338 53566 46340 53618
rect 46284 53564 46340 53566
rect 45948 52892 46004 52948
rect 45052 51324 45108 51380
rect 45612 51266 45668 51268
rect 45612 51214 45614 51266
rect 45614 51214 45666 51266
rect 45666 51214 45668 51266
rect 45612 51212 45668 51214
rect 45836 51154 45892 51156
rect 45836 51102 45838 51154
rect 45838 51102 45890 51154
rect 45890 51102 45892 51154
rect 45836 51100 45892 51102
rect 46732 51938 46788 51940
rect 46732 51886 46734 51938
rect 46734 51886 46786 51938
rect 46786 51886 46788 51938
rect 46732 51884 46788 51886
rect 46396 51436 46452 51492
rect 46732 51100 46788 51156
rect 46620 50764 46676 50820
rect 46172 50482 46228 50484
rect 46172 50430 46174 50482
rect 46174 50430 46226 50482
rect 46226 50430 46228 50482
rect 46172 50428 46228 50430
rect 43596 50316 43652 50372
rect 43036 49756 43092 49812
rect 43932 49810 43988 49812
rect 43932 49758 43934 49810
rect 43934 49758 43986 49810
rect 43986 49758 43988 49810
rect 43932 49756 43988 49758
rect 42924 49698 42980 49700
rect 42924 49646 42926 49698
rect 42926 49646 42978 49698
rect 42978 49646 42980 49698
rect 42924 49644 42980 49646
rect 43036 49250 43092 49252
rect 43036 49198 43038 49250
rect 43038 49198 43090 49250
rect 43090 49198 43092 49250
rect 43036 49196 43092 49198
rect 37996 48802 38052 48804
rect 37996 48750 37998 48802
rect 37998 48750 38050 48802
rect 38050 48750 38052 48802
rect 37996 48748 38052 48750
rect 44492 49698 44548 49700
rect 44492 49646 44494 49698
rect 44494 49646 44546 49698
rect 44546 49646 44548 49698
rect 44492 49644 44548 49646
rect 44940 49698 44996 49700
rect 44940 49646 44942 49698
rect 44942 49646 44994 49698
rect 44994 49646 44996 49698
rect 44940 49644 44996 49646
rect 45388 49644 45444 49700
rect 43372 48412 43428 48468
rect 43820 48636 43876 48692
rect 39228 47068 39284 47124
rect 37100 46956 37156 47012
rect 37772 46956 37828 47012
rect 37100 46396 37156 46452
rect 37548 45836 37604 45892
rect 36876 44604 36932 44660
rect 39676 46674 39732 46676
rect 39676 46622 39678 46674
rect 39678 46622 39730 46674
rect 39730 46622 39732 46674
rect 39676 46620 39732 46622
rect 42140 47346 42196 47348
rect 42140 47294 42142 47346
rect 42142 47294 42194 47346
rect 42194 47294 42196 47346
rect 42140 47292 42196 47294
rect 43372 48242 43428 48244
rect 43372 48190 43374 48242
rect 43374 48190 43426 48242
rect 43426 48190 43428 48242
rect 43372 48188 43428 48190
rect 44044 48354 44100 48356
rect 44044 48302 44046 48354
rect 44046 48302 44098 48354
rect 44098 48302 44100 48354
rect 44044 48300 44100 48302
rect 44828 48636 44884 48692
rect 44156 48188 44212 48244
rect 43260 48018 43316 48020
rect 43260 47966 43262 48018
rect 43262 47966 43314 48018
rect 43314 47966 43316 48018
rect 43260 47964 43316 47966
rect 44268 47570 44324 47572
rect 44268 47518 44270 47570
rect 44270 47518 44322 47570
rect 44322 47518 44324 47570
rect 44268 47516 44324 47518
rect 43260 47068 43316 47124
rect 44492 47068 44548 47124
rect 40236 46562 40292 46564
rect 40236 46510 40238 46562
rect 40238 46510 40290 46562
rect 40290 46510 40292 46562
rect 40236 46508 40292 46510
rect 38332 45836 38388 45892
rect 39228 45890 39284 45892
rect 39228 45838 39230 45890
rect 39230 45838 39282 45890
rect 39282 45838 39284 45890
rect 39228 45836 39284 45838
rect 39564 45388 39620 45444
rect 39900 45890 39956 45892
rect 39900 45838 39902 45890
rect 39902 45838 39954 45890
rect 39954 45838 39956 45890
rect 39900 45836 39956 45838
rect 40460 45890 40516 45892
rect 40460 45838 40462 45890
rect 40462 45838 40514 45890
rect 40514 45838 40516 45890
rect 40460 45836 40516 45838
rect 48748 53730 48804 53732
rect 48748 53678 48750 53730
rect 48750 53678 48802 53730
rect 48802 53678 48804 53730
rect 48748 53676 48804 53678
rect 48860 53564 48916 53620
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 49980 52946 50036 52948
rect 49980 52894 49982 52946
rect 49982 52894 50034 52946
rect 50034 52894 50036 52946
rect 49980 52892 50036 52894
rect 48860 52332 48916 52388
rect 47068 51938 47124 51940
rect 47068 51886 47070 51938
rect 47070 51886 47122 51938
rect 47122 51886 47124 51938
rect 47068 51884 47124 51886
rect 46956 51324 47012 51380
rect 47516 51100 47572 51156
rect 47068 50988 47124 51044
rect 47068 50706 47124 50708
rect 47068 50654 47070 50706
rect 47070 50654 47122 50706
rect 47122 50654 47124 50706
rect 47068 50652 47124 50654
rect 47516 50594 47572 50596
rect 47516 50542 47518 50594
rect 47518 50542 47570 50594
rect 47570 50542 47572 50594
rect 47516 50540 47572 50542
rect 47292 50482 47348 50484
rect 47292 50430 47294 50482
rect 47294 50430 47346 50482
rect 47346 50430 47348 50482
rect 47292 50428 47348 50430
rect 48076 51436 48132 51492
rect 47740 50876 47796 50932
rect 47964 51100 48020 51156
rect 47628 49868 47684 49924
rect 47740 50428 47796 50484
rect 46844 49196 46900 49252
rect 45388 48076 45444 48132
rect 46060 48300 46116 48356
rect 44716 47516 44772 47572
rect 45388 47516 45444 47572
rect 44828 47346 44884 47348
rect 44828 47294 44830 47346
rect 44830 47294 44882 47346
rect 44882 47294 44884 47346
rect 44828 47292 44884 47294
rect 45836 47516 45892 47572
rect 44940 46620 44996 46676
rect 41692 46562 41748 46564
rect 41692 46510 41694 46562
rect 41694 46510 41746 46562
rect 41746 46510 41748 46562
rect 41692 46508 41748 46510
rect 45052 46172 45108 46228
rect 40348 45276 40404 45332
rect 36092 44268 36148 44324
rect 36988 43596 37044 43652
rect 36204 42140 36260 42196
rect 37772 43596 37828 43652
rect 37996 44268 38052 44324
rect 38444 44210 38500 44212
rect 38444 44158 38446 44210
rect 38446 44158 38498 44210
rect 38498 44158 38500 44210
rect 38444 44156 38500 44158
rect 39564 45218 39620 45220
rect 39564 45166 39566 45218
rect 39566 45166 39618 45218
rect 39618 45166 39620 45218
rect 39564 45164 39620 45166
rect 39676 44882 39732 44884
rect 39676 44830 39678 44882
rect 39678 44830 39730 44882
rect 39730 44830 39732 44882
rect 39676 44828 39732 44830
rect 38780 44322 38836 44324
rect 38780 44270 38782 44322
rect 38782 44270 38834 44322
rect 38834 44270 38836 44322
rect 38780 44268 38836 44270
rect 39788 44322 39844 44324
rect 39788 44270 39790 44322
rect 39790 44270 39842 44322
rect 39842 44270 39844 44322
rect 39788 44268 39844 44270
rect 39116 44156 39172 44212
rect 38668 43820 38724 43876
rect 38444 43538 38500 43540
rect 38444 43486 38446 43538
rect 38446 43486 38498 43538
rect 38498 43486 38500 43538
rect 38444 43484 38500 43486
rect 38556 43260 38612 43316
rect 36204 41298 36260 41300
rect 36204 41246 36206 41298
rect 36206 41246 36258 41298
rect 36258 41246 36260 41298
rect 36204 41244 36260 41246
rect 36092 41132 36148 41188
rect 36988 42028 37044 42084
rect 37772 42140 37828 42196
rect 38892 43538 38948 43540
rect 38892 43486 38894 43538
rect 38894 43486 38946 43538
rect 38946 43486 38948 43538
rect 38892 43484 38948 43486
rect 38780 42700 38836 42756
rect 39228 44044 39284 44100
rect 40124 44044 40180 44100
rect 39900 43820 39956 43876
rect 39564 43708 39620 43764
rect 39900 43426 39956 43428
rect 39900 43374 39902 43426
rect 39902 43374 39954 43426
rect 39954 43374 39956 43426
rect 39900 43372 39956 43374
rect 40348 43650 40404 43652
rect 40348 43598 40350 43650
rect 40350 43598 40402 43650
rect 40402 43598 40404 43650
rect 40348 43596 40404 43598
rect 40236 43260 40292 43316
rect 39004 42812 39060 42868
rect 40348 42754 40404 42756
rect 40348 42702 40350 42754
rect 40350 42702 40402 42754
rect 40402 42702 40404 42754
rect 40348 42700 40404 42702
rect 39900 42588 39956 42644
rect 40124 42476 40180 42532
rect 40124 42028 40180 42084
rect 38332 41858 38388 41860
rect 38332 41806 38334 41858
rect 38334 41806 38386 41858
rect 38386 41806 38388 41858
rect 38332 41804 38388 41806
rect 39900 41804 39956 41860
rect 38332 41356 38388 41412
rect 37100 41244 37156 41300
rect 36652 41020 36708 41076
rect 37212 41074 37268 41076
rect 37212 41022 37214 41074
rect 37214 41022 37266 41074
rect 37266 41022 37268 41074
rect 37212 41020 37268 41022
rect 37100 40684 37156 40740
rect 37324 40348 37380 40404
rect 35980 39228 36036 39284
rect 36428 39730 36484 39732
rect 36428 39678 36430 39730
rect 36430 39678 36482 39730
rect 36482 39678 36484 39730
rect 36428 39676 36484 39678
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34636 38220 34692 38276
rect 34300 36540 34356 36596
rect 33964 36428 34020 36484
rect 33740 35810 33796 35812
rect 33740 35758 33742 35810
rect 33742 35758 33794 35810
rect 33794 35758 33796 35810
rect 33740 35756 33796 35758
rect 33852 35308 33908 35364
rect 33628 33964 33684 34020
rect 33180 33404 33236 33460
rect 30044 31948 30100 32004
rect 32396 32620 32452 32676
rect 31052 31836 31108 31892
rect 29708 31218 29764 31220
rect 29708 31166 29710 31218
rect 29710 31166 29762 31218
rect 29762 31166 29764 31218
rect 29708 31164 29764 31166
rect 31052 31164 31108 31220
rect 29708 30940 29764 30996
rect 30156 30770 30212 30772
rect 30156 30718 30158 30770
rect 30158 30718 30210 30770
rect 30210 30718 30212 30770
rect 30156 30716 30212 30718
rect 29372 30044 29428 30100
rect 28252 28866 28308 28868
rect 28252 28814 28254 28866
rect 28254 28814 28306 28866
rect 28306 28814 28308 28866
rect 28252 28812 28308 28814
rect 29148 28866 29204 28868
rect 29148 28814 29150 28866
rect 29150 28814 29202 28866
rect 29202 28814 29204 28866
rect 29148 28812 29204 28814
rect 28364 27692 28420 27748
rect 28476 26236 28532 26292
rect 30604 30044 30660 30100
rect 32508 31724 32564 31780
rect 33292 32620 33348 32676
rect 34076 34690 34132 34692
rect 34076 34638 34078 34690
rect 34078 34638 34130 34690
rect 34130 34638 34132 34690
rect 34076 34636 34132 34638
rect 33964 34076 34020 34132
rect 34300 35420 34356 35476
rect 34412 37548 34468 37604
rect 35084 37826 35140 37828
rect 35084 37774 35086 37826
rect 35086 37774 35138 37826
rect 35138 37774 35140 37826
rect 35084 37772 35140 37774
rect 39116 41020 39172 41076
rect 39340 41580 39396 41636
rect 38108 40962 38164 40964
rect 38108 40910 38110 40962
rect 38110 40910 38162 40962
rect 38162 40910 38164 40962
rect 38108 40908 38164 40910
rect 37100 39676 37156 39732
rect 38892 40962 38948 40964
rect 38892 40910 38894 40962
rect 38894 40910 38946 40962
rect 38946 40910 38948 40962
rect 38892 40908 38948 40910
rect 37884 40684 37940 40740
rect 38444 40626 38500 40628
rect 38444 40574 38446 40626
rect 38446 40574 38498 40626
rect 38498 40574 38500 40626
rect 38444 40572 38500 40574
rect 39004 40402 39060 40404
rect 39004 40350 39006 40402
rect 39006 40350 39058 40402
rect 39058 40350 39060 40402
rect 39004 40348 39060 40350
rect 39788 41020 39844 41076
rect 39340 40908 39396 40964
rect 39788 40514 39844 40516
rect 39788 40462 39790 40514
rect 39790 40462 39842 40514
rect 39842 40462 39844 40514
rect 39788 40460 39844 40462
rect 39228 40348 39284 40404
rect 37884 40290 37940 40292
rect 37884 40238 37886 40290
rect 37886 40238 37938 40290
rect 37938 40238 37940 40290
rect 37884 40236 37940 40238
rect 39900 39900 39956 39956
rect 38892 39788 38948 39844
rect 37548 39116 37604 39172
rect 36764 38332 36820 38388
rect 36204 37826 36260 37828
rect 36204 37774 36206 37826
rect 36206 37774 36258 37826
rect 36258 37774 36260 37826
rect 36204 37772 36260 37774
rect 36540 37884 36596 37940
rect 35084 37212 35140 37268
rect 35868 37548 35924 37604
rect 34636 36988 34692 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 36428 37548 36484 37604
rect 36204 37378 36260 37380
rect 36204 37326 36206 37378
rect 36206 37326 36258 37378
rect 36258 37326 36260 37378
rect 36204 37324 36260 37326
rect 36540 36652 36596 36708
rect 37212 38050 37268 38052
rect 37212 37998 37214 38050
rect 37214 37998 37266 38050
rect 37266 37998 37268 38050
rect 37212 37996 37268 37998
rect 38220 38834 38276 38836
rect 38220 38782 38222 38834
rect 38222 38782 38274 38834
rect 38274 38782 38276 38834
rect 38220 38780 38276 38782
rect 37884 38332 37940 38388
rect 38108 38332 38164 38388
rect 37324 37938 37380 37940
rect 37324 37886 37326 37938
rect 37326 37886 37378 37938
rect 37378 37886 37380 37938
rect 37324 37884 37380 37886
rect 37100 37660 37156 37716
rect 36876 37324 36932 37380
rect 36092 36482 36148 36484
rect 36092 36430 36094 36482
rect 36094 36430 36146 36482
rect 36146 36430 36148 36482
rect 36092 36428 36148 36430
rect 35756 36092 35812 36148
rect 34972 35308 35028 35364
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34860 35026 34916 35028
rect 34860 34974 34862 35026
rect 34862 34974 34914 35026
rect 34914 34974 34916 35026
rect 34860 34972 34916 34974
rect 37212 37378 37268 37380
rect 37212 37326 37214 37378
rect 37214 37326 37266 37378
rect 37266 37326 37268 37378
rect 37212 37324 37268 37326
rect 37660 37378 37716 37380
rect 37660 37326 37662 37378
rect 37662 37326 37714 37378
rect 37714 37326 37716 37378
rect 37660 37324 37716 37326
rect 37324 36764 37380 36820
rect 37212 36706 37268 36708
rect 37212 36654 37214 36706
rect 37214 36654 37266 36706
rect 37266 36654 37268 36706
rect 37212 36652 37268 36654
rect 36988 36482 37044 36484
rect 36988 36430 36990 36482
rect 36990 36430 37042 36482
rect 37042 36430 37044 36482
rect 36988 36428 37044 36430
rect 36652 35810 36708 35812
rect 36652 35758 36654 35810
rect 36654 35758 36706 35810
rect 36706 35758 36708 35810
rect 36652 35756 36708 35758
rect 37548 35698 37604 35700
rect 37548 35646 37550 35698
rect 37550 35646 37602 35698
rect 37602 35646 37604 35698
rect 37548 35644 37604 35646
rect 38220 38220 38276 38276
rect 38108 38108 38164 38164
rect 38220 38050 38276 38052
rect 38220 37998 38222 38050
rect 38222 37998 38274 38050
rect 38274 37998 38276 38050
rect 38220 37996 38276 37998
rect 38220 37548 38276 37604
rect 37996 37378 38052 37380
rect 37996 37326 37998 37378
rect 37998 37326 38050 37378
rect 38050 37326 38052 37378
rect 37996 37324 38052 37326
rect 38668 38834 38724 38836
rect 38668 38782 38670 38834
rect 38670 38782 38722 38834
rect 38722 38782 38724 38834
rect 38668 38780 38724 38782
rect 38444 38332 38500 38388
rect 38668 37100 38724 37156
rect 35756 34748 35812 34804
rect 34188 34076 34244 34132
rect 34300 34636 34356 34692
rect 34300 33628 34356 33684
rect 34412 33964 34468 34020
rect 33516 32284 33572 32340
rect 33068 31836 33124 31892
rect 32172 30716 32228 30772
rect 32172 30492 32228 30548
rect 32284 29426 32340 29428
rect 32284 29374 32286 29426
rect 32286 29374 32338 29426
rect 32338 29374 32340 29426
rect 32284 29372 32340 29374
rect 33068 29426 33124 29428
rect 33068 29374 33070 29426
rect 33070 29374 33122 29426
rect 33122 29374 33124 29426
rect 33068 29372 33124 29374
rect 32508 29314 32564 29316
rect 32508 29262 32510 29314
rect 32510 29262 32562 29314
rect 32562 29262 32564 29314
rect 32508 29260 32564 29262
rect 33068 28924 33124 28980
rect 33404 30492 33460 30548
rect 33740 31500 33796 31556
rect 28812 27692 28868 27748
rect 31836 27916 31892 27972
rect 28700 26290 28756 26292
rect 28700 26238 28702 26290
rect 28702 26238 28754 26290
rect 28754 26238 28756 26290
rect 28700 26236 28756 26238
rect 28588 25340 28644 25396
rect 27020 22258 27076 22260
rect 27020 22206 27022 22258
rect 27022 22206 27074 22258
rect 27074 22206 27076 22258
rect 27020 22204 27076 22206
rect 26908 22092 26964 22148
rect 27692 22370 27748 22372
rect 27692 22318 27694 22370
rect 27694 22318 27746 22370
rect 27746 22318 27748 22370
rect 27692 22316 27748 22318
rect 27580 22092 27636 22148
rect 27468 21644 27524 21700
rect 26236 20188 26292 20244
rect 26124 20076 26180 20132
rect 27132 20300 27188 20356
rect 27020 20076 27076 20132
rect 25900 18060 25956 18116
rect 26348 18956 26404 19012
rect 26460 18844 26516 18900
rect 26012 17836 26068 17892
rect 26460 18396 26516 18452
rect 26012 16994 26068 16996
rect 26012 16942 26014 16994
rect 26014 16942 26066 16994
rect 26066 16942 26068 16994
rect 26012 16940 26068 16942
rect 27020 19010 27076 19012
rect 27020 18958 27022 19010
rect 27022 18958 27074 19010
rect 27074 18958 27076 19010
rect 27020 18956 27076 18958
rect 28588 22988 28644 23044
rect 28924 25004 28980 25060
rect 28476 22204 28532 22260
rect 28588 21196 28644 21252
rect 28588 20914 28644 20916
rect 28588 20862 28590 20914
rect 28590 20862 28642 20914
rect 28642 20862 28644 20914
rect 28588 20860 28644 20862
rect 28700 21308 28756 21364
rect 28252 20300 28308 20356
rect 27580 19292 27636 19348
rect 28476 19740 28532 19796
rect 27804 18732 27860 18788
rect 27692 18620 27748 18676
rect 27692 18396 27748 18452
rect 27244 18172 27300 18228
rect 26796 18060 26852 18116
rect 26572 17666 26628 17668
rect 26572 17614 26574 17666
rect 26574 17614 26626 17666
rect 26626 17614 26628 17666
rect 26572 17612 26628 17614
rect 27132 17276 27188 17332
rect 26460 17106 26516 17108
rect 26460 17054 26462 17106
rect 26462 17054 26514 17106
rect 26514 17054 26516 17106
rect 26460 17052 26516 17054
rect 27244 17164 27300 17220
rect 25676 16828 25732 16884
rect 25676 16380 25732 16436
rect 25004 16044 25060 16100
rect 25452 16044 25508 16100
rect 24556 15986 24612 15988
rect 24556 15934 24558 15986
rect 24558 15934 24610 15986
rect 24610 15934 24612 15986
rect 24556 15932 24612 15934
rect 25340 15932 25396 15988
rect 24780 15820 24836 15876
rect 24892 15708 24948 15764
rect 24556 15314 24612 15316
rect 24556 15262 24558 15314
rect 24558 15262 24610 15314
rect 24610 15262 24612 15314
rect 24556 15260 24612 15262
rect 24220 14476 24276 14532
rect 24108 13804 24164 13860
rect 24220 14140 24276 14196
rect 24108 13468 24164 13524
rect 23772 12572 23828 12628
rect 23884 12348 23940 12404
rect 24444 13634 24500 13636
rect 24444 13582 24446 13634
rect 24446 13582 24498 13634
rect 24498 13582 24500 13634
rect 24444 13580 24500 13582
rect 24444 13356 24500 13412
rect 24444 13020 24500 13076
rect 24332 12962 24388 12964
rect 24332 12910 24334 12962
rect 24334 12910 24386 12962
rect 24386 12910 24388 12962
rect 24332 12908 24388 12910
rect 24668 14700 24724 14756
rect 23996 11676 24052 11732
rect 24332 11564 24388 11620
rect 24332 9772 24388 9828
rect 23772 8428 23828 8484
rect 23660 8316 23716 8372
rect 23100 6860 23156 6916
rect 23548 6914 23604 6916
rect 23548 6862 23550 6914
rect 23550 6862 23602 6914
rect 23602 6862 23604 6914
rect 23548 6860 23604 6862
rect 22764 6802 22820 6804
rect 22764 6750 22766 6802
rect 22766 6750 22818 6802
rect 22818 6750 22820 6802
rect 22764 6748 22820 6750
rect 19852 5234 19908 5236
rect 19852 5182 19854 5234
rect 19854 5182 19906 5234
rect 19906 5182 19908 5234
rect 19852 5180 19908 5182
rect 21532 5292 21588 5348
rect 20860 5180 20916 5236
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 22652 6188 22708 6244
rect 22652 5964 22708 6020
rect 24332 8764 24388 8820
rect 25004 15484 25060 15540
rect 25676 16098 25732 16100
rect 25676 16046 25678 16098
rect 25678 16046 25730 16098
rect 25730 16046 25732 16098
rect 25676 16044 25732 16046
rect 25676 15708 25732 15764
rect 26124 16716 26180 16772
rect 26124 16156 26180 16212
rect 27356 17388 27412 17444
rect 26908 16882 26964 16884
rect 26908 16830 26910 16882
rect 26910 16830 26962 16882
rect 26962 16830 26964 16882
rect 26908 16828 26964 16830
rect 26684 16268 26740 16324
rect 26796 16604 26852 16660
rect 26684 16098 26740 16100
rect 26684 16046 26686 16098
rect 26686 16046 26738 16098
rect 26738 16046 26740 16098
rect 26684 16044 26740 16046
rect 25788 15596 25844 15652
rect 25228 15314 25284 15316
rect 25228 15262 25230 15314
rect 25230 15262 25282 15314
rect 25282 15262 25284 15314
rect 25228 15260 25284 15262
rect 25452 15148 25508 15204
rect 25116 14140 25172 14196
rect 25228 15036 25284 15092
rect 25116 12962 25172 12964
rect 25116 12910 25118 12962
rect 25118 12910 25170 12962
rect 25170 12910 25172 12962
rect 25116 12908 25172 12910
rect 25004 12850 25060 12852
rect 25004 12798 25006 12850
rect 25006 12798 25058 12850
rect 25058 12798 25060 12850
rect 25004 12796 25060 12798
rect 24780 12124 24836 12180
rect 24556 11506 24612 11508
rect 24556 11454 24558 11506
rect 24558 11454 24610 11506
rect 24610 11454 24612 11506
rect 24556 11452 24612 11454
rect 24668 10780 24724 10836
rect 24556 9996 24612 10052
rect 24668 9884 24724 9940
rect 24556 9042 24612 9044
rect 24556 8990 24558 9042
rect 24558 8990 24610 9042
rect 24610 8990 24612 9042
rect 24556 8988 24612 8990
rect 23996 8258 24052 8260
rect 23996 8206 23998 8258
rect 23998 8206 24050 8258
rect 24050 8206 24052 8258
rect 23996 8204 24052 8206
rect 23884 8092 23940 8148
rect 24220 7756 24276 7812
rect 23996 7644 24052 7700
rect 23996 6690 24052 6692
rect 23996 6638 23998 6690
rect 23998 6638 24050 6690
rect 24050 6638 24052 6690
rect 23996 6636 24052 6638
rect 24220 6748 24276 6804
rect 24668 8258 24724 8260
rect 24668 8206 24670 8258
rect 24670 8206 24722 8258
rect 24722 8206 24724 8258
rect 24668 8204 24724 8206
rect 24444 8146 24500 8148
rect 24444 8094 24446 8146
rect 24446 8094 24498 8146
rect 24498 8094 24500 8146
rect 24444 8092 24500 8094
rect 25340 13970 25396 13972
rect 25340 13918 25342 13970
rect 25342 13918 25394 13970
rect 25394 13918 25396 13970
rect 25340 13916 25396 13918
rect 26124 15596 26180 15652
rect 25900 15372 25956 15428
rect 26460 15372 26516 15428
rect 26348 15314 26404 15316
rect 26348 15262 26350 15314
rect 26350 15262 26402 15314
rect 26402 15262 26404 15314
rect 26348 15260 26404 15262
rect 25564 14028 25620 14084
rect 25564 13468 25620 13524
rect 25564 13020 25620 13076
rect 25676 12962 25732 12964
rect 25676 12910 25678 12962
rect 25678 12910 25730 12962
rect 25730 12910 25732 12962
rect 25676 12908 25732 12910
rect 25340 12796 25396 12852
rect 26348 14700 26404 14756
rect 26124 14588 26180 14644
rect 26012 13356 26068 13412
rect 26684 15874 26740 15876
rect 26684 15822 26686 15874
rect 26686 15822 26738 15874
rect 26738 15822 26740 15874
rect 26684 15820 26740 15822
rect 26684 15596 26740 15652
rect 27916 17500 27972 17556
rect 27804 17442 27860 17444
rect 27804 17390 27806 17442
rect 27806 17390 27858 17442
rect 27858 17390 27860 17442
rect 27804 17388 27860 17390
rect 27580 17052 27636 17108
rect 27580 16882 27636 16884
rect 27580 16830 27582 16882
rect 27582 16830 27634 16882
rect 27634 16830 27636 16882
rect 27580 16828 27636 16830
rect 26796 15260 26852 15316
rect 26684 15148 26740 15204
rect 27020 16098 27076 16100
rect 27020 16046 27022 16098
rect 27022 16046 27074 16098
rect 27074 16046 27076 16098
rect 27020 16044 27076 16046
rect 27804 16044 27860 16100
rect 28252 17276 28308 17332
rect 28140 16322 28196 16324
rect 28140 16270 28142 16322
rect 28142 16270 28194 16322
rect 28194 16270 28196 16322
rect 28140 16268 28196 16270
rect 27356 15932 27412 15988
rect 27468 15596 27524 15652
rect 28028 15932 28084 15988
rect 27132 15372 27188 15428
rect 27468 15426 27524 15428
rect 27468 15374 27470 15426
rect 27470 15374 27522 15426
rect 27522 15374 27524 15426
rect 27468 15372 27524 15374
rect 26796 14754 26852 14756
rect 26796 14702 26798 14754
rect 26798 14702 26850 14754
rect 26850 14702 26852 14754
rect 26796 14700 26852 14702
rect 27132 13970 27188 13972
rect 27132 13918 27134 13970
rect 27134 13918 27186 13970
rect 27186 13918 27188 13970
rect 27132 13916 27188 13918
rect 26796 13746 26852 13748
rect 26796 13694 26798 13746
rect 26798 13694 26850 13746
rect 26850 13694 26852 13746
rect 26796 13692 26852 13694
rect 27132 13746 27188 13748
rect 27132 13694 27134 13746
rect 27134 13694 27186 13746
rect 27186 13694 27188 13746
rect 27132 13692 27188 13694
rect 26348 13522 26404 13524
rect 26348 13470 26350 13522
rect 26350 13470 26402 13522
rect 26402 13470 26404 13522
rect 26348 13468 26404 13470
rect 26908 13468 26964 13524
rect 26236 13074 26292 13076
rect 26236 13022 26238 13074
rect 26238 13022 26290 13074
rect 26290 13022 26292 13074
rect 26236 13020 26292 13022
rect 26124 12684 26180 12740
rect 27692 14530 27748 14532
rect 27692 14478 27694 14530
rect 27694 14478 27746 14530
rect 27746 14478 27748 14530
rect 27692 14476 27748 14478
rect 33292 28812 33348 28868
rect 32284 27916 32340 27972
rect 32396 28364 32452 28420
rect 31612 27074 31668 27076
rect 31612 27022 31614 27074
rect 31614 27022 31666 27074
rect 31666 27022 31668 27074
rect 31612 27020 31668 27022
rect 32284 27074 32340 27076
rect 32284 27022 32286 27074
rect 32286 27022 32338 27074
rect 32338 27022 32340 27074
rect 32284 27020 32340 27022
rect 29596 26796 29652 26852
rect 32508 27858 32564 27860
rect 32508 27806 32510 27858
rect 32510 27806 32562 27858
rect 32562 27806 32564 27858
rect 32508 27804 32564 27806
rect 33740 29596 33796 29652
rect 33516 29260 33572 29316
rect 33516 28588 33572 28644
rect 32956 28530 33012 28532
rect 32956 28478 32958 28530
rect 32958 28478 33010 28530
rect 33010 28478 33012 28530
rect 32956 28476 33012 28478
rect 34076 29596 34132 29652
rect 34300 31612 34356 31668
rect 33964 29426 34020 29428
rect 33964 29374 33966 29426
rect 33966 29374 34018 29426
rect 34018 29374 34020 29426
rect 33964 29372 34020 29374
rect 34748 33852 34804 33908
rect 35084 33852 35140 33908
rect 34972 33628 35028 33684
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35420 33234 35476 33236
rect 35420 33182 35422 33234
rect 35422 33182 35474 33234
rect 35474 33182 35476 33234
rect 35420 33180 35476 33182
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 36428 34972 36484 35028
rect 35980 33740 36036 33796
rect 35532 31948 35588 32004
rect 37884 34972 37940 35028
rect 36540 34242 36596 34244
rect 36540 34190 36542 34242
rect 36542 34190 36594 34242
rect 36594 34190 36596 34242
rect 36540 34188 36596 34190
rect 36428 33906 36484 33908
rect 36428 33854 36430 33906
rect 36430 33854 36482 33906
rect 36482 33854 36484 33906
rect 36428 33852 36484 33854
rect 36204 33234 36260 33236
rect 36204 33182 36206 33234
rect 36206 33182 36258 33234
rect 36258 33182 36260 33234
rect 36204 33180 36260 33182
rect 36428 33122 36484 33124
rect 36428 33070 36430 33122
rect 36430 33070 36482 33122
rect 36482 33070 36484 33122
rect 36428 33068 36484 33070
rect 36428 32732 36484 32788
rect 36204 31890 36260 31892
rect 36204 31838 36206 31890
rect 36206 31838 36258 31890
rect 36258 31838 36260 31890
rect 36204 31836 36260 31838
rect 35644 31724 35700 31780
rect 34524 31554 34580 31556
rect 34524 31502 34526 31554
rect 34526 31502 34578 31554
rect 34578 31502 34580 31554
rect 34524 31500 34580 31502
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 30156 35252 30212
rect 34636 30044 34692 30100
rect 34524 29260 34580 29316
rect 35196 29650 35252 29652
rect 35196 29598 35198 29650
rect 35198 29598 35250 29650
rect 35250 29598 35252 29650
rect 35196 29596 35252 29598
rect 35308 29426 35364 29428
rect 35308 29374 35310 29426
rect 35310 29374 35362 29426
rect 35362 29374 35364 29426
rect 35308 29372 35364 29374
rect 33852 28700 33908 28756
rect 34076 28642 34132 28644
rect 34076 28590 34078 28642
rect 34078 28590 34130 28642
rect 34130 28590 34132 28642
rect 34076 28588 34132 28590
rect 33740 28476 33796 28532
rect 33628 27468 33684 27524
rect 33740 27298 33796 27300
rect 33740 27246 33742 27298
rect 33742 27246 33794 27298
rect 33794 27246 33796 27298
rect 33740 27244 33796 27246
rect 33292 27074 33348 27076
rect 33292 27022 33294 27074
rect 33294 27022 33346 27074
rect 33346 27022 33348 27074
rect 33292 27020 33348 27022
rect 29372 25394 29428 25396
rect 29372 25342 29374 25394
rect 29374 25342 29426 25394
rect 29426 25342 29428 25394
rect 29372 25340 29428 25342
rect 29596 25340 29652 25396
rect 29148 24668 29204 24724
rect 29148 24220 29204 24276
rect 29372 23772 29428 23828
rect 31612 26290 31668 26292
rect 31612 26238 31614 26290
rect 31614 26238 31666 26290
rect 31666 26238 31668 26290
rect 31612 26236 31668 26238
rect 32060 26290 32116 26292
rect 32060 26238 32062 26290
rect 32062 26238 32114 26290
rect 32114 26238 32116 26290
rect 32060 26236 32116 26238
rect 30492 26124 30548 26180
rect 32508 26066 32564 26068
rect 32508 26014 32510 26066
rect 32510 26014 32562 26066
rect 32562 26014 32564 26066
rect 32508 26012 32564 26014
rect 32620 25340 32676 25396
rect 32060 25228 32116 25284
rect 32508 24946 32564 24948
rect 32508 24894 32510 24946
rect 32510 24894 32562 24946
rect 32562 24894 32564 24946
rect 32508 24892 32564 24894
rect 32284 24556 32340 24612
rect 30156 24220 30212 24276
rect 29820 22258 29876 22260
rect 29820 22206 29822 22258
rect 29822 22206 29874 22258
rect 29874 22206 29876 22258
rect 29820 22204 29876 22206
rect 29708 21810 29764 21812
rect 29708 21758 29710 21810
rect 29710 21758 29762 21810
rect 29762 21758 29764 21810
rect 29708 21756 29764 21758
rect 29036 21362 29092 21364
rect 29036 21310 29038 21362
rect 29038 21310 29090 21362
rect 29090 21310 29092 21362
rect 29036 21308 29092 21310
rect 29708 20972 29764 21028
rect 30044 21698 30100 21700
rect 30044 21646 30046 21698
rect 30046 21646 30098 21698
rect 30098 21646 30100 21698
rect 30044 21644 30100 21646
rect 29148 20860 29204 20916
rect 28924 20130 28980 20132
rect 28924 20078 28926 20130
rect 28926 20078 28978 20130
rect 28978 20078 28980 20130
rect 28924 20076 28980 20078
rect 28924 18620 28980 18676
rect 28364 15484 28420 15540
rect 28364 15314 28420 15316
rect 28364 15262 28366 15314
rect 28366 15262 28418 15314
rect 28418 15262 28420 15314
rect 28364 15260 28420 15262
rect 28364 14028 28420 14084
rect 27916 13746 27972 13748
rect 27916 13694 27918 13746
rect 27918 13694 27970 13746
rect 27970 13694 27972 13746
rect 27916 13692 27972 13694
rect 27468 13634 27524 13636
rect 27468 13582 27470 13634
rect 27470 13582 27522 13634
rect 27522 13582 27524 13634
rect 27468 13580 27524 13582
rect 28476 13468 28532 13524
rect 27356 13356 27412 13412
rect 27244 13132 27300 13188
rect 25340 11900 25396 11956
rect 25452 11394 25508 11396
rect 25452 11342 25454 11394
rect 25454 11342 25506 11394
rect 25506 11342 25508 11394
rect 25452 11340 25508 11342
rect 26348 12066 26404 12068
rect 26348 12014 26350 12066
rect 26350 12014 26402 12066
rect 26402 12014 26404 12066
rect 26348 12012 26404 12014
rect 27580 12908 27636 12964
rect 26460 11900 26516 11956
rect 26348 11788 26404 11844
rect 25228 10220 25284 10276
rect 25004 9938 25060 9940
rect 25004 9886 25006 9938
rect 25006 9886 25058 9938
rect 25058 9886 25060 9938
rect 25004 9884 25060 9886
rect 25228 9548 25284 9604
rect 24668 7698 24724 7700
rect 24668 7646 24670 7698
rect 24670 7646 24722 7698
rect 24722 7646 24724 7698
rect 24668 7644 24724 7646
rect 26012 9996 26068 10052
rect 25564 9602 25620 9604
rect 25564 9550 25566 9602
rect 25566 9550 25618 9602
rect 25618 9550 25620 9602
rect 25564 9548 25620 9550
rect 25228 8988 25284 9044
rect 25900 9100 25956 9156
rect 26012 9212 26068 9268
rect 25564 8652 25620 8708
rect 25340 8428 25396 8484
rect 23884 6188 23940 6244
rect 23212 5292 23268 5348
rect 22092 5180 22148 5236
rect 21756 5068 21812 5124
rect 22876 5122 22932 5124
rect 22876 5070 22878 5122
rect 22878 5070 22930 5122
rect 22930 5070 22932 5122
rect 22876 5068 22932 5070
rect 24332 6188 24388 6244
rect 24220 5964 24276 6020
rect 24892 6802 24948 6804
rect 24892 6750 24894 6802
rect 24894 6750 24946 6802
rect 24946 6750 24948 6802
rect 24892 6748 24948 6750
rect 26124 6636 26180 6692
rect 26236 9436 26292 9492
rect 27020 12572 27076 12628
rect 27020 12178 27076 12180
rect 27020 12126 27022 12178
rect 27022 12126 27074 12178
rect 27074 12126 27076 12178
rect 27020 12124 27076 12126
rect 26908 12066 26964 12068
rect 26908 12014 26910 12066
rect 26910 12014 26962 12066
rect 26962 12014 26964 12066
rect 26908 12012 26964 12014
rect 26684 11394 26740 11396
rect 26684 11342 26686 11394
rect 26686 11342 26738 11394
rect 26738 11342 26740 11394
rect 26684 11340 26740 11342
rect 28028 12908 28084 12964
rect 27916 12178 27972 12180
rect 27916 12126 27918 12178
rect 27918 12126 27970 12178
rect 27970 12126 27972 12178
rect 27916 12124 27972 12126
rect 27468 11340 27524 11396
rect 26796 9996 26852 10052
rect 26572 9436 26628 9492
rect 26460 8988 26516 9044
rect 26908 8876 26964 8932
rect 26460 8652 26516 8708
rect 26684 8652 26740 8708
rect 26572 8428 26628 8484
rect 24220 4956 24276 5012
rect 26236 5794 26292 5796
rect 26236 5742 26238 5794
rect 26238 5742 26290 5794
rect 26290 5742 26292 5794
rect 26236 5740 26292 5742
rect 25340 4956 25396 5012
rect 25676 4562 25732 4564
rect 25676 4510 25678 4562
rect 25678 4510 25730 4562
rect 25730 4510 25732 4562
rect 25676 4508 25732 4510
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 27132 8316 27188 8372
rect 28252 10668 28308 10724
rect 27692 10444 27748 10500
rect 28588 10498 28644 10500
rect 28588 10446 28590 10498
rect 28590 10446 28642 10498
rect 28642 10446 28644 10498
rect 28588 10444 28644 10446
rect 29484 20300 29540 20356
rect 29820 20300 29876 20356
rect 29484 19964 29540 20020
rect 29260 19794 29316 19796
rect 29260 19742 29262 19794
rect 29262 19742 29314 19794
rect 29314 19742 29316 19794
rect 29260 19740 29316 19742
rect 30044 20188 30100 20244
rect 33180 26850 33236 26852
rect 33180 26798 33182 26850
rect 33182 26798 33234 26850
rect 33234 26798 33236 26850
rect 33180 26796 33236 26798
rect 33628 26908 33684 26964
rect 33516 26796 33572 26852
rect 33516 26290 33572 26292
rect 33516 26238 33518 26290
rect 33518 26238 33570 26290
rect 33570 26238 33572 26290
rect 33516 26236 33572 26238
rect 33628 26460 33684 26516
rect 33180 26178 33236 26180
rect 33180 26126 33182 26178
rect 33182 26126 33234 26178
rect 33234 26126 33236 26178
rect 33180 26124 33236 26126
rect 33068 26012 33124 26068
rect 33068 25228 33124 25284
rect 31276 23826 31332 23828
rect 31276 23774 31278 23826
rect 31278 23774 31330 23826
rect 31330 23774 31332 23826
rect 31276 23772 31332 23774
rect 30716 22988 30772 23044
rect 30492 21810 30548 21812
rect 30492 21758 30494 21810
rect 30494 21758 30546 21810
rect 30546 21758 30548 21810
rect 30492 21756 30548 21758
rect 30380 21644 30436 21700
rect 33628 25340 33684 25396
rect 33964 27468 34020 27524
rect 34748 28700 34804 28756
rect 34188 27244 34244 27300
rect 34076 26796 34132 26852
rect 34524 26962 34580 26964
rect 34524 26910 34526 26962
rect 34526 26910 34578 26962
rect 34578 26910 34580 26962
rect 34524 26908 34580 26910
rect 34412 26460 34468 26516
rect 33292 24668 33348 24724
rect 33852 25116 33908 25172
rect 34076 24722 34132 24724
rect 34076 24670 34078 24722
rect 34078 24670 34130 24722
rect 34130 24670 34132 24722
rect 34076 24668 34132 24670
rect 33516 24556 33572 24612
rect 34300 25004 34356 25060
rect 34524 26066 34580 26068
rect 34524 26014 34526 26066
rect 34526 26014 34578 26066
rect 34578 26014 34580 26066
rect 34524 26012 34580 26014
rect 34636 24892 34692 24948
rect 34412 24780 34468 24836
rect 33852 23548 33908 23604
rect 34300 23378 34356 23380
rect 34300 23326 34302 23378
rect 34302 23326 34354 23378
rect 34354 23326 34356 23378
rect 34300 23324 34356 23326
rect 34188 23266 34244 23268
rect 34188 23214 34190 23266
rect 34190 23214 34242 23266
rect 34242 23214 34244 23266
rect 34188 23212 34244 23214
rect 33516 23100 33572 23156
rect 34748 23660 34804 23716
rect 34748 23100 34804 23156
rect 34636 22988 34692 23044
rect 32732 22428 32788 22484
rect 34188 22482 34244 22484
rect 34188 22430 34190 22482
rect 34190 22430 34242 22482
rect 34242 22430 34244 22482
rect 34188 22428 34244 22430
rect 33292 21868 33348 21924
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35308 28418 35364 28420
rect 35308 28366 35310 28418
rect 35310 28366 35362 28418
rect 35362 28366 35364 28418
rect 35308 28364 35364 28366
rect 35084 27916 35140 27972
rect 35532 27804 35588 27860
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35756 30210 35812 30212
rect 35756 30158 35758 30210
rect 35758 30158 35810 30210
rect 35810 30158 35812 30210
rect 35756 30156 35812 30158
rect 36988 33292 37044 33348
rect 37100 33068 37156 33124
rect 37100 32732 37156 32788
rect 37212 33180 37268 33236
rect 36652 32284 36708 32340
rect 36428 28364 36484 28420
rect 36092 27804 36148 27860
rect 36540 27970 36596 27972
rect 36540 27918 36542 27970
rect 36542 27918 36594 27970
rect 36594 27918 36596 27970
rect 36540 27916 36596 27918
rect 36428 27074 36484 27076
rect 36428 27022 36430 27074
rect 36430 27022 36482 27074
rect 36482 27022 36484 27074
rect 36428 27020 36484 27022
rect 36204 26962 36260 26964
rect 36204 26910 36206 26962
rect 36206 26910 36258 26962
rect 36258 26910 36260 26962
rect 36204 26908 36260 26910
rect 35644 26850 35700 26852
rect 35644 26798 35646 26850
rect 35646 26798 35698 26850
rect 35698 26798 35700 26850
rect 35644 26796 35700 26798
rect 35308 26290 35364 26292
rect 35308 26238 35310 26290
rect 35310 26238 35362 26290
rect 35362 26238 35364 26290
rect 35308 26236 35364 26238
rect 35980 26290 36036 26292
rect 35980 26238 35982 26290
rect 35982 26238 36034 26290
rect 36034 26238 36036 26290
rect 35980 26236 36036 26238
rect 35532 26012 35588 26068
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34972 25116 35028 25172
rect 35420 24834 35476 24836
rect 35420 24782 35422 24834
rect 35422 24782 35474 24834
rect 35474 24782 35476 24834
rect 35420 24780 35476 24782
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35420 24162 35476 24164
rect 35420 24110 35422 24162
rect 35422 24110 35474 24162
rect 35474 24110 35476 24162
rect 35420 24108 35476 24110
rect 35532 23996 35588 24052
rect 35644 23660 35700 23716
rect 35868 23826 35924 23828
rect 35868 23774 35870 23826
rect 35870 23774 35922 23826
rect 35922 23774 35924 23826
rect 35868 23772 35924 23774
rect 35756 23100 35812 23156
rect 35084 22988 35140 23044
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34972 22540 35028 22596
rect 35532 22428 35588 22484
rect 34972 21868 35028 21924
rect 32396 21308 32452 21364
rect 29820 17388 29876 17444
rect 29820 16828 29876 16884
rect 29596 16492 29652 16548
rect 29260 15372 29316 15428
rect 30156 18620 30212 18676
rect 31836 18284 31892 18340
rect 32284 18338 32340 18340
rect 32284 18286 32286 18338
rect 32286 18286 32338 18338
rect 32338 18286 32340 18338
rect 32284 18284 32340 18286
rect 30044 16268 30100 16324
rect 30380 16156 30436 16212
rect 31276 16994 31332 16996
rect 31276 16942 31278 16994
rect 31278 16942 31330 16994
rect 31330 16942 31332 16994
rect 31276 16940 31332 16942
rect 36316 24108 36372 24164
rect 36204 23772 36260 23828
rect 38108 34188 38164 34244
rect 38332 35756 38388 35812
rect 40236 40012 40292 40068
rect 39900 39564 39956 39620
rect 38892 37436 38948 37492
rect 39452 36540 39508 36596
rect 38780 35644 38836 35700
rect 38780 35196 38836 35252
rect 39788 37548 39844 37604
rect 41468 45836 41524 45892
rect 44044 45890 44100 45892
rect 44044 45838 44046 45890
rect 44046 45838 44098 45890
rect 44098 45838 44100 45890
rect 44044 45836 44100 45838
rect 44380 45276 44436 45332
rect 41468 45218 41524 45220
rect 41468 45166 41470 45218
rect 41470 45166 41522 45218
rect 41522 45166 41524 45218
rect 41468 45164 41524 45166
rect 42364 45218 42420 45220
rect 42364 45166 42366 45218
rect 42366 45166 42418 45218
rect 42418 45166 42420 45218
rect 42364 45164 42420 45166
rect 41580 45106 41636 45108
rect 41580 45054 41582 45106
rect 41582 45054 41634 45106
rect 41634 45054 41636 45106
rect 41580 45052 41636 45054
rect 42476 45106 42532 45108
rect 42476 45054 42478 45106
rect 42478 45054 42530 45106
rect 42530 45054 42532 45106
rect 42476 45052 42532 45054
rect 44492 45836 44548 45892
rect 44940 45890 44996 45892
rect 44940 45838 44942 45890
rect 44942 45838 44994 45890
rect 44994 45838 44996 45890
rect 44940 45836 44996 45838
rect 46396 48076 46452 48132
rect 46508 47852 46564 47908
rect 46060 47458 46116 47460
rect 46060 47406 46062 47458
rect 46062 47406 46114 47458
rect 46114 47406 46116 47458
rect 46060 47404 46116 47406
rect 48860 51212 48916 51268
rect 48188 50988 48244 51044
rect 48076 50594 48132 50596
rect 48076 50542 48078 50594
rect 48078 50542 48130 50594
rect 48130 50542 48132 50594
rect 48076 50540 48132 50542
rect 48300 50594 48356 50596
rect 48300 50542 48302 50594
rect 48302 50542 48354 50594
rect 48354 50542 48356 50594
rect 48300 50540 48356 50542
rect 47964 50428 48020 50484
rect 49420 52274 49476 52276
rect 49420 52222 49422 52274
rect 49422 52222 49474 52274
rect 49474 52222 49476 52274
rect 49420 52220 49476 52222
rect 51436 52892 51492 52948
rect 49980 52220 50036 52276
rect 49756 52108 49812 52164
rect 49196 51996 49252 52052
rect 49420 51996 49476 52052
rect 49308 50594 49364 50596
rect 49308 50542 49310 50594
rect 49310 50542 49362 50594
rect 49362 50542 49364 50594
rect 49308 50540 49364 50542
rect 49420 50876 49476 50932
rect 48524 50204 48580 50260
rect 48748 49922 48804 49924
rect 48748 49870 48750 49922
rect 48750 49870 48802 49922
rect 48802 49870 48804 49922
rect 48748 49868 48804 49870
rect 49084 49756 49140 49812
rect 49084 49250 49140 49252
rect 49084 49198 49086 49250
rect 49086 49198 49138 49250
rect 49138 49198 49140 49250
rect 49084 49196 49140 49198
rect 47740 48636 47796 48692
rect 46956 48354 47012 48356
rect 46956 48302 46958 48354
rect 46958 48302 47010 48354
rect 47010 48302 47012 48354
rect 46956 48300 47012 48302
rect 46060 47068 46116 47124
rect 45836 46674 45892 46676
rect 45836 46622 45838 46674
rect 45838 46622 45890 46674
rect 45890 46622 45892 46674
rect 45836 46620 45892 46622
rect 46172 46562 46228 46564
rect 46172 46510 46174 46562
rect 46174 46510 46226 46562
rect 46226 46510 46228 46562
rect 46172 46508 46228 46510
rect 46620 46562 46676 46564
rect 46620 46510 46622 46562
rect 46622 46510 46674 46562
rect 46674 46510 46676 46562
rect 46620 46508 46676 46510
rect 45724 46450 45780 46452
rect 45724 46398 45726 46450
rect 45726 46398 45778 46450
rect 45778 46398 45780 46450
rect 45724 46396 45780 46398
rect 45836 46172 45892 46228
rect 47292 47964 47348 48020
rect 47180 47404 47236 47460
rect 47964 48188 48020 48244
rect 48636 48242 48692 48244
rect 48636 48190 48638 48242
rect 48638 48190 48690 48242
rect 48690 48190 48692 48242
rect 48636 48188 48692 48190
rect 48860 48130 48916 48132
rect 48860 48078 48862 48130
rect 48862 48078 48914 48130
rect 48914 48078 48916 48130
rect 48860 48076 48916 48078
rect 48188 47964 48244 48020
rect 47404 46732 47460 46788
rect 47068 46172 47124 46228
rect 47292 46396 47348 46452
rect 46620 45890 46676 45892
rect 46620 45838 46622 45890
rect 46622 45838 46674 45890
rect 46674 45838 46676 45890
rect 46620 45836 46676 45838
rect 49980 51996 50036 52052
rect 50204 51996 50260 52052
rect 49868 51436 49924 51492
rect 49868 51100 49924 51156
rect 50652 52332 50708 52388
rect 50764 52162 50820 52164
rect 50764 52110 50766 52162
rect 50766 52110 50818 52162
rect 50818 52110 50820 52162
rect 50764 52108 50820 52110
rect 50988 51938 51044 51940
rect 50988 51886 50990 51938
rect 50990 51886 51042 51938
rect 51042 51886 51044 51938
rect 50988 51884 51044 51886
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 51884 52220 51940 52276
rect 50876 51436 50932 51492
rect 50316 51100 50372 51156
rect 49980 50428 50036 50484
rect 50764 50652 50820 50708
rect 51660 51378 51716 51380
rect 51660 51326 51662 51378
rect 51662 51326 51714 51378
rect 51714 51326 51716 51378
rect 51660 51324 51716 51326
rect 52444 51884 52500 51940
rect 51772 51212 51828 51268
rect 52668 51324 52724 51380
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 49532 49084 49588 49140
rect 49756 49196 49812 49252
rect 50540 49250 50596 49252
rect 50540 49198 50542 49250
rect 50542 49198 50594 49250
rect 50594 49198 50596 49250
rect 50540 49196 50596 49198
rect 54572 51266 54628 51268
rect 54572 51214 54574 51266
rect 54574 51214 54626 51266
rect 54626 51214 54628 51266
rect 54572 51212 54628 51214
rect 55580 50706 55636 50708
rect 55580 50654 55582 50706
rect 55582 50654 55634 50706
rect 55634 50654 55636 50706
rect 55580 50652 55636 50654
rect 51324 50428 51380 50484
rect 53452 50482 53508 50484
rect 53452 50430 53454 50482
rect 53454 50430 53506 50482
rect 53506 50430 53508 50482
rect 53452 50428 53508 50430
rect 49868 49084 49924 49140
rect 49084 47852 49140 47908
rect 48524 47516 48580 47572
rect 48300 47458 48356 47460
rect 48300 47406 48302 47458
rect 48302 47406 48354 47458
rect 48354 47406 48356 47458
rect 48300 47404 48356 47406
rect 48748 47292 48804 47348
rect 48636 47068 48692 47124
rect 49084 46732 49140 46788
rect 48860 46562 48916 46564
rect 48860 46510 48862 46562
rect 48862 46510 48914 46562
rect 48914 46510 48916 46562
rect 48860 46508 48916 46510
rect 49644 48412 49700 48468
rect 49756 47964 49812 48020
rect 50092 47852 50148 47908
rect 49644 47628 49700 47684
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50652 48412 50708 48468
rect 50540 48300 50596 48356
rect 49868 47458 49924 47460
rect 49868 47406 49870 47458
rect 49870 47406 49922 47458
rect 49922 47406 49924 47458
rect 49868 47404 49924 47406
rect 50316 47404 50372 47460
rect 51324 48412 51380 48468
rect 51436 48300 51492 48356
rect 50652 47964 50708 48020
rect 51548 48076 51604 48132
rect 51548 47628 51604 47684
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50988 46956 51044 47012
rect 51212 47458 51268 47460
rect 51212 47406 51214 47458
rect 51214 47406 51266 47458
rect 51266 47406 51268 47458
rect 51212 47404 51268 47406
rect 53340 48130 53396 48132
rect 53340 48078 53342 48130
rect 53342 48078 53394 48130
rect 53394 48078 53396 48130
rect 53340 48076 53396 48078
rect 51660 46956 51716 47012
rect 50540 46674 50596 46676
rect 50540 46622 50542 46674
rect 50542 46622 50594 46674
rect 50594 46622 50596 46674
rect 50540 46620 50596 46622
rect 49308 46060 49364 46116
rect 42364 44828 42420 44884
rect 41804 44044 41860 44100
rect 44156 44098 44212 44100
rect 44156 44046 44158 44098
rect 44158 44046 44210 44098
rect 44210 44046 44212 44098
rect 44156 44044 44212 44046
rect 41244 43538 41300 43540
rect 41244 43486 41246 43538
rect 41246 43486 41298 43538
rect 41298 43486 41300 43538
rect 41244 43484 41300 43486
rect 41468 43372 41524 43428
rect 40796 43260 40852 43316
rect 41132 42812 41188 42868
rect 42140 43538 42196 43540
rect 42140 43486 42142 43538
rect 42142 43486 42194 43538
rect 42194 43486 42196 43538
rect 42140 43484 42196 43486
rect 43260 43484 43316 43540
rect 41804 42252 41860 42308
rect 42028 41186 42084 41188
rect 42028 41134 42030 41186
rect 42030 41134 42082 41186
rect 42082 41134 42084 41186
rect 42028 41132 42084 41134
rect 41580 41074 41636 41076
rect 41580 41022 41582 41074
rect 41582 41022 41634 41074
rect 41634 41022 41636 41074
rect 41580 41020 41636 41022
rect 41692 40962 41748 40964
rect 41692 40910 41694 40962
rect 41694 40910 41746 40962
rect 41746 40910 41748 40962
rect 41692 40908 41748 40910
rect 41916 40572 41972 40628
rect 41356 40402 41412 40404
rect 41356 40350 41358 40402
rect 41358 40350 41410 40402
rect 41410 40350 41412 40402
rect 41356 40348 41412 40350
rect 42476 40908 42532 40964
rect 41580 40124 41636 40180
rect 41468 39900 41524 39956
rect 41244 39618 41300 39620
rect 41244 39566 41246 39618
rect 41246 39566 41298 39618
rect 41298 39566 41300 39618
rect 41244 39564 41300 39566
rect 40684 39452 40740 39508
rect 40348 36594 40404 36596
rect 40348 36542 40350 36594
rect 40350 36542 40402 36594
rect 40402 36542 40404 36594
rect 40348 36540 40404 36542
rect 39676 36428 39732 36484
rect 41916 39730 41972 39732
rect 41916 39678 41918 39730
rect 41918 39678 41970 39730
rect 41970 39678 41972 39730
rect 41916 39676 41972 39678
rect 41580 38834 41636 38836
rect 41580 38782 41582 38834
rect 41582 38782 41634 38834
rect 41634 38782 41636 38834
rect 41580 38780 41636 38782
rect 40908 37154 40964 37156
rect 40908 37102 40910 37154
rect 40910 37102 40962 37154
rect 40962 37102 40964 37154
rect 40908 37100 40964 37102
rect 40684 36092 40740 36148
rect 40236 35420 40292 35476
rect 38780 34130 38836 34132
rect 38780 34078 38782 34130
rect 38782 34078 38834 34130
rect 38834 34078 38836 34130
rect 38780 34076 38836 34078
rect 39900 34076 39956 34132
rect 39676 33068 39732 33124
rect 37324 31836 37380 31892
rect 36988 31666 37044 31668
rect 36988 31614 36990 31666
rect 36990 31614 37042 31666
rect 37042 31614 37044 31666
rect 36988 31612 37044 31614
rect 37548 31778 37604 31780
rect 37548 31726 37550 31778
rect 37550 31726 37602 31778
rect 37602 31726 37604 31778
rect 37548 31724 37604 31726
rect 38220 31666 38276 31668
rect 38220 31614 38222 31666
rect 38222 31614 38274 31666
rect 38274 31614 38276 31666
rect 38220 31612 38276 31614
rect 38220 30210 38276 30212
rect 38220 30158 38222 30210
rect 38222 30158 38274 30210
rect 38274 30158 38276 30210
rect 38220 30156 38276 30158
rect 36988 29036 37044 29092
rect 37660 29036 37716 29092
rect 37212 28642 37268 28644
rect 37212 28590 37214 28642
rect 37214 28590 37266 28642
rect 37266 28590 37268 28642
rect 37212 28588 37268 28590
rect 36988 27020 37044 27076
rect 37324 27804 37380 27860
rect 38108 29820 38164 29876
rect 38108 28588 38164 28644
rect 37772 27244 37828 27300
rect 38668 31836 38724 31892
rect 39900 31836 39956 31892
rect 39228 31612 39284 31668
rect 38556 28028 38612 28084
rect 38556 27858 38612 27860
rect 38556 27806 38558 27858
rect 38558 27806 38610 27858
rect 38610 27806 38612 27858
rect 38556 27804 38612 27806
rect 39004 30434 39060 30436
rect 39004 30382 39006 30434
rect 39006 30382 39058 30434
rect 39058 30382 39060 30434
rect 39004 30380 39060 30382
rect 39228 29820 39284 29876
rect 39676 31500 39732 31556
rect 40124 31724 40180 31780
rect 39900 31106 39956 31108
rect 39900 31054 39902 31106
rect 39902 31054 39954 31106
rect 39954 31054 39956 31106
rect 39900 31052 39956 31054
rect 41020 35196 41076 35252
rect 40908 34130 40964 34132
rect 40908 34078 40910 34130
rect 40910 34078 40962 34130
rect 40962 34078 40964 34130
rect 40908 34076 40964 34078
rect 42028 38780 42084 38836
rect 42140 38892 42196 38948
rect 43036 41916 43092 41972
rect 44380 42364 44436 42420
rect 44044 41970 44100 41972
rect 44044 41918 44046 41970
rect 44046 41918 44098 41970
rect 44098 41918 44100 41970
rect 44044 41916 44100 41918
rect 43372 41132 43428 41188
rect 42812 40236 42868 40292
rect 42700 40124 42756 40180
rect 43260 40012 43316 40068
rect 43708 40962 43764 40964
rect 43708 40910 43710 40962
rect 43710 40910 43762 40962
rect 43762 40910 43764 40962
rect 43708 40908 43764 40910
rect 42588 39676 42644 39732
rect 42700 38780 42756 38836
rect 43372 38668 43428 38724
rect 44268 41074 44324 41076
rect 44268 41022 44270 41074
rect 44270 41022 44322 41074
rect 44322 41022 44324 41074
rect 44268 41020 44324 41022
rect 44156 40962 44212 40964
rect 44156 40910 44158 40962
rect 44158 40910 44210 40962
rect 44210 40910 44212 40962
rect 44156 40908 44212 40910
rect 44380 40684 44436 40740
rect 43820 40460 43876 40516
rect 44044 40236 44100 40292
rect 43708 39394 43764 39396
rect 43708 39342 43710 39394
rect 43710 39342 43762 39394
rect 43762 39342 43764 39394
rect 43708 39340 43764 39342
rect 43932 38668 43988 38724
rect 41692 37100 41748 37156
rect 42140 35196 42196 35252
rect 42028 34130 42084 34132
rect 42028 34078 42030 34130
rect 42030 34078 42082 34130
rect 42082 34078 42084 34130
rect 42028 34076 42084 34078
rect 41692 33628 41748 33684
rect 44268 39506 44324 39508
rect 44268 39454 44270 39506
rect 44270 39454 44322 39506
rect 44322 39454 44324 39506
rect 44268 39452 44324 39454
rect 44156 38556 44212 38612
rect 42812 37938 42868 37940
rect 42812 37886 42814 37938
rect 42814 37886 42866 37938
rect 42866 37886 42868 37938
rect 42812 37884 42868 37886
rect 43708 37884 43764 37940
rect 43484 37436 43540 37492
rect 43820 37436 43876 37492
rect 43932 37324 43988 37380
rect 42476 37100 42532 37156
rect 42476 36652 42532 36708
rect 43484 36988 43540 37044
rect 42812 36092 42868 36148
rect 42588 34076 42644 34132
rect 43372 36876 43428 36932
rect 43932 36876 43988 36932
rect 43484 36428 43540 36484
rect 40348 33122 40404 33124
rect 40348 33070 40350 33122
rect 40350 33070 40402 33122
rect 40402 33070 40404 33122
rect 40348 33068 40404 33070
rect 41468 32172 41524 32228
rect 40348 31836 40404 31892
rect 40236 30716 40292 30772
rect 40348 31554 40404 31556
rect 40348 31502 40350 31554
rect 40350 31502 40402 31554
rect 40402 31502 40404 31554
rect 40348 31500 40404 31502
rect 39900 29538 39956 29540
rect 39900 29486 39902 29538
rect 39902 29486 39954 29538
rect 39954 29486 39956 29538
rect 39900 29484 39956 29486
rect 40908 31500 40964 31556
rect 41468 31836 41524 31892
rect 41804 31724 41860 31780
rect 41916 31836 41972 31892
rect 41804 31500 41860 31556
rect 41580 31052 41636 31108
rect 41020 30716 41076 30772
rect 40572 30604 40628 30660
rect 39340 28588 39396 28644
rect 40572 28588 40628 28644
rect 40348 28028 40404 28084
rect 38892 27356 38948 27412
rect 38332 27132 38388 27188
rect 39564 27244 39620 27300
rect 37212 26908 37268 26964
rect 37436 26908 37492 26964
rect 37100 26236 37156 26292
rect 37212 26178 37268 26180
rect 37212 26126 37214 26178
rect 37214 26126 37266 26178
rect 37266 26126 37268 26178
rect 37212 26124 37268 26126
rect 36988 25116 37044 25172
rect 36652 24108 36708 24164
rect 36428 23548 36484 23604
rect 36540 23212 36596 23268
rect 36652 23100 36708 23156
rect 38668 26850 38724 26852
rect 38668 26798 38670 26850
rect 38670 26798 38722 26850
rect 38722 26798 38724 26850
rect 38668 26796 38724 26798
rect 38892 26850 38948 26852
rect 38892 26798 38894 26850
rect 38894 26798 38946 26850
rect 38946 26798 38948 26850
rect 38892 26796 38948 26798
rect 37324 24050 37380 24052
rect 37324 23998 37326 24050
rect 37326 23998 37378 24050
rect 37378 23998 37380 24050
rect 37324 23996 37380 23998
rect 37100 23772 37156 23828
rect 36204 22540 36260 22596
rect 36428 22540 36484 22596
rect 37212 23938 37268 23940
rect 37212 23886 37214 23938
rect 37214 23886 37266 23938
rect 37266 23886 37268 23938
rect 37212 23884 37268 23886
rect 37212 23212 37268 23268
rect 37884 25116 37940 25172
rect 38220 24780 38276 24836
rect 38556 24780 38612 24836
rect 37996 24668 38052 24724
rect 38332 23938 38388 23940
rect 38332 23886 38334 23938
rect 38334 23886 38386 23938
rect 38386 23886 38388 23938
rect 38332 23884 38388 23886
rect 37772 23324 37828 23380
rect 38444 23660 38500 23716
rect 38892 24834 38948 24836
rect 38892 24782 38894 24834
rect 38894 24782 38946 24834
rect 38946 24782 38948 24834
rect 38892 24780 38948 24782
rect 38556 23378 38612 23380
rect 38556 23326 38558 23378
rect 38558 23326 38610 23378
rect 38610 23326 38612 23378
rect 38556 23324 38612 23326
rect 38668 24556 38724 24612
rect 38668 23436 38724 23492
rect 38220 23100 38276 23156
rect 37436 22540 37492 22596
rect 37324 22482 37380 22484
rect 37324 22430 37326 22482
rect 37326 22430 37378 22482
rect 37378 22430 37380 22482
rect 37324 22428 37380 22430
rect 33740 21532 33796 21588
rect 33516 21362 33572 21364
rect 33516 21310 33518 21362
rect 33518 21310 33570 21362
rect 33570 21310 33572 21362
rect 33516 21308 33572 21310
rect 34076 20188 34132 20244
rect 33292 18508 33348 18564
rect 33516 19292 33572 19348
rect 32732 18172 32788 18228
rect 31948 16828 32004 16884
rect 31612 16658 31668 16660
rect 31612 16606 31614 16658
rect 31614 16606 31666 16658
rect 31666 16606 31668 16658
rect 31612 16604 31668 16606
rect 30828 16380 30884 16436
rect 30828 16210 30884 16212
rect 30828 16158 30830 16210
rect 30830 16158 30882 16210
rect 30882 16158 30884 16210
rect 30828 16156 30884 16158
rect 31836 16156 31892 16212
rect 31276 15260 31332 15316
rect 27580 9154 27636 9156
rect 27580 9102 27582 9154
rect 27582 9102 27634 9154
rect 27634 9102 27636 9154
rect 27580 9100 27636 9102
rect 27804 9042 27860 9044
rect 27804 8990 27806 9042
rect 27806 8990 27858 9042
rect 27858 8990 27860 9042
rect 27804 8988 27860 8990
rect 27916 8316 27972 8372
rect 28588 8370 28644 8372
rect 28588 8318 28590 8370
rect 28590 8318 28642 8370
rect 28642 8318 28644 8370
rect 28588 8316 28644 8318
rect 29596 13468 29652 13524
rect 29372 12962 29428 12964
rect 29372 12910 29374 12962
rect 29374 12910 29426 12962
rect 29426 12910 29428 12962
rect 29372 12908 29428 12910
rect 29708 12962 29764 12964
rect 29708 12910 29710 12962
rect 29710 12910 29762 12962
rect 29762 12910 29764 12962
rect 29708 12908 29764 12910
rect 29596 11900 29652 11956
rect 29148 9212 29204 9268
rect 29260 11282 29316 11284
rect 29260 11230 29262 11282
rect 29262 11230 29314 11282
rect 29314 11230 29316 11282
rect 29260 11228 29316 11230
rect 33740 18956 33796 19012
rect 35644 21532 35700 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 32956 16380 33012 16436
rect 32732 16044 32788 16100
rect 32508 15484 32564 15540
rect 31500 14700 31556 14756
rect 29932 13580 29988 13636
rect 30604 14306 30660 14308
rect 30604 14254 30606 14306
rect 30606 14254 30658 14306
rect 30658 14254 30660 14306
rect 30604 14252 30660 14254
rect 31276 13468 31332 13524
rect 29932 12402 29988 12404
rect 29932 12350 29934 12402
rect 29934 12350 29986 12402
rect 29986 12350 29988 12402
rect 29932 12348 29988 12350
rect 31612 14252 31668 14308
rect 33404 15538 33460 15540
rect 33404 15486 33406 15538
rect 33406 15486 33458 15538
rect 33458 15486 33460 15538
rect 33404 15484 33460 15486
rect 33180 13746 33236 13748
rect 33180 13694 33182 13746
rect 33182 13694 33234 13746
rect 33234 13694 33236 13746
rect 33180 13692 33236 13694
rect 33628 18284 33684 18340
rect 36988 21868 37044 21924
rect 35420 19852 35476 19908
rect 35532 20300 35588 20356
rect 34636 19346 34692 19348
rect 34636 19294 34638 19346
rect 34638 19294 34690 19346
rect 34690 19294 34692 19346
rect 34636 19292 34692 19294
rect 34300 18284 34356 18340
rect 34860 18338 34916 18340
rect 34860 18286 34862 18338
rect 34862 18286 34914 18338
rect 34914 18286 34916 18338
rect 34860 18284 34916 18286
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 39116 24332 39172 24388
rect 39004 23548 39060 23604
rect 38556 22594 38612 22596
rect 38556 22542 38558 22594
rect 38558 22542 38610 22594
rect 38610 22542 38612 22594
rect 38556 22540 38612 22542
rect 40012 27356 40068 27412
rect 40012 27020 40068 27076
rect 40460 27186 40516 27188
rect 40460 27134 40462 27186
rect 40462 27134 40514 27186
rect 40514 27134 40516 27186
rect 40460 27132 40516 27134
rect 40348 27020 40404 27076
rect 40124 26290 40180 26292
rect 40124 26238 40126 26290
rect 40126 26238 40178 26290
rect 40178 26238 40180 26290
rect 40124 26236 40180 26238
rect 39900 26124 39956 26180
rect 40124 25618 40180 25620
rect 40124 25566 40126 25618
rect 40126 25566 40178 25618
rect 40178 25566 40180 25618
rect 40124 25564 40180 25566
rect 39900 25506 39956 25508
rect 39900 25454 39902 25506
rect 39902 25454 39954 25506
rect 39954 25454 39956 25506
rect 39900 25452 39956 25454
rect 40012 24722 40068 24724
rect 40012 24670 40014 24722
rect 40014 24670 40066 24722
rect 40066 24670 40068 24722
rect 40012 24668 40068 24670
rect 39564 23548 39620 23604
rect 39564 23324 39620 23380
rect 39116 22540 39172 22596
rect 38892 22428 38948 22484
rect 37772 21868 37828 21924
rect 39788 23324 39844 23380
rect 39676 23266 39732 23268
rect 39676 23214 39678 23266
rect 39678 23214 39730 23266
rect 39730 23214 39732 23266
rect 39676 23212 39732 23214
rect 39900 22428 39956 22484
rect 40012 23436 40068 23492
rect 40236 23548 40292 23604
rect 40124 22482 40180 22484
rect 40124 22430 40126 22482
rect 40126 22430 40178 22482
rect 40178 22430 40180 22482
rect 40124 22428 40180 22430
rect 40012 22316 40068 22372
rect 41132 28924 41188 28980
rect 41692 30716 41748 30772
rect 41692 29260 41748 29316
rect 41468 28700 41524 28756
rect 42924 32508 42980 32564
rect 42812 32396 42868 32452
rect 41916 28754 41972 28756
rect 41916 28702 41918 28754
rect 41918 28702 41970 28754
rect 41970 28702 41972 28754
rect 41916 28700 41972 28702
rect 42028 30210 42084 30212
rect 42028 30158 42030 30210
rect 42030 30158 42082 30210
rect 42082 30158 42084 30210
rect 42028 30156 42084 30158
rect 41244 27634 41300 27636
rect 41244 27582 41246 27634
rect 41246 27582 41298 27634
rect 41298 27582 41300 27634
rect 41244 27580 41300 27582
rect 41804 27580 41860 27636
rect 42028 27468 42084 27524
rect 42588 30716 42644 30772
rect 43372 32786 43428 32788
rect 43372 32734 43374 32786
rect 43374 32734 43426 32786
rect 43426 32734 43428 32786
rect 43372 32732 43428 32734
rect 43596 33740 43652 33796
rect 43708 35196 43764 35252
rect 44156 36652 44212 36708
rect 44828 44604 44884 44660
rect 44828 43596 44884 43652
rect 46844 43650 46900 43652
rect 46844 43598 46846 43650
rect 46846 43598 46898 43650
rect 46898 43598 46900 43650
rect 46844 43596 46900 43598
rect 45388 43426 45444 43428
rect 45388 43374 45390 43426
rect 45390 43374 45442 43426
rect 45442 43374 45444 43426
rect 45388 43372 45444 43374
rect 46172 43426 46228 43428
rect 46172 43374 46174 43426
rect 46174 43374 46226 43426
rect 46226 43374 46228 43426
rect 46172 43372 46228 43374
rect 45276 42978 45332 42980
rect 45276 42926 45278 42978
rect 45278 42926 45330 42978
rect 45330 42926 45332 42978
rect 45276 42924 45332 42926
rect 46060 43314 46116 43316
rect 46060 43262 46062 43314
rect 46062 43262 46114 43314
rect 46114 43262 46116 43314
rect 46060 43260 46116 43262
rect 44828 40796 44884 40852
rect 45052 40572 45108 40628
rect 45052 40236 45108 40292
rect 44828 39452 44884 39508
rect 44604 39340 44660 39396
rect 45388 40124 45444 40180
rect 45612 42252 45668 42308
rect 47292 43260 47348 43316
rect 51548 46114 51604 46116
rect 51548 46062 51550 46114
rect 51550 46062 51602 46114
rect 51602 46062 51604 46114
rect 51548 46060 51604 46062
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 51660 44940 51716 44996
rect 48188 44098 48244 44100
rect 48188 44046 48190 44098
rect 48190 44046 48242 44098
rect 48242 44046 48244 44098
rect 48188 44044 48244 44046
rect 46620 42812 46676 42868
rect 46284 42754 46340 42756
rect 46284 42702 46286 42754
rect 46286 42702 46338 42754
rect 46338 42702 46340 42754
rect 46284 42700 46340 42702
rect 46844 42588 46900 42644
rect 46620 42028 46676 42084
rect 46060 41746 46116 41748
rect 46060 41694 46062 41746
rect 46062 41694 46114 41746
rect 46114 41694 46116 41746
rect 46060 41692 46116 41694
rect 45948 40684 46004 40740
rect 45612 40236 45668 40292
rect 45052 39340 45108 39396
rect 44604 38834 44660 38836
rect 44604 38782 44606 38834
rect 44606 38782 44658 38834
rect 44658 38782 44660 38834
rect 44604 38780 44660 38782
rect 44828 38556 44884 38612
rect 45388 39618 45444 39620
rect 45388 39566 45390 39618
rect 45390 39566 45442 39618
rect 45442 39566 45444 39618
rect 45388 39564 45444 39566
rect 45612 39452 45668 39508
rect 45276 39394 45332 39396
rect 45276 39342 45278 39394
rect 45278 39342 45330 39394
rect 45330 39342 45332 39394
rect 45276 39340 45332 39342
rect 45500 39394 45556 39396
rect 45500 39342 45502 39394
rect 45502 39342 45554 39394
rect 45554 39342 45556 39394
rect 45500 39340 45556 39342
rect 45836 39506 45892 39508
rect 45836 39454 45838 39506
rect 45838 39454 45890 39506
rect 45890 39454 45892 39506
rect 45836 39452 45892 39454
rect 46844 40684 46900 40740
rect 46284 39900 46340 39956
rect 46956 40236 47012 40292
rect 46284 39618 46340 39620
rect 46284 39566 46286 39618
rect 46286 39566 46338 39618
rect 46338 39566 46340 39618
rect 46284 39564 46340 39566
rect 46172 39506 46228 39508
rect 46172 39454 46174 39506
rect 46174 39454 46226 39506
rect 46226 39454 46228 39506
rect 46172 39452 46228 39454
rect 45948 38946 46004 38948
rect 45948 38894 45950 38946
rect 45950 38894 46002 38946
rect 46002 38894 46004 38946
rect 45948 38892 46004 38894
rect 45724 38668 45780 38724
rect 45052 38108 45108 38164
rect 44492 37772 44548 37828
rect 44828 37772 44884 37828
rect 44380 37324 44436 37380
rect 45164 37938 45220 37940
rect 45164 37886 45166 37938
rect 45166 37886 45218 37938
rect 45218 37886 45220 37938
rect 45164 37884 45220 37886
rect 45388 37938 45444 37940
rect 45388 37886 45390 37938
rect 45390 37886 45442 37938
rect 45442 37886 45444 37938
rect 45388 37884 45444 37886
rect 46396 38722 46452 38724
rect 46396 38670 46398 38722
rect 46398 38670 46450 38722
rect 46450 38670 46452 38722
rect 46396 38668 46452 38670
rect 45836 38108 45892 38164
rect 45612 37884 45668 37940
rect 45276 37154 45332 37156
rect 45276 37102 45278 37154
rect 45278 37102 45330 37154
rect 45330 37102 45332 37154
rect 45276 37100 45332 37102
rect 45836 37938 45892 37940
rect 45836 37886 45838 37938
rect 45838 37886 45890 37938
rect 45890 37886 45892 37938
rect 45836 37884 45892 37886
rect 46396 37938 46452 37940
rect 46396 37886 46398 37938
rect 46398 37886 46450 37938
rect 46450 37886 46452 37938
rect 46396 37884 46452 37886
rect 45500 36988 45556 37044
rect 45724 37436 45780 37492
rect 45276 36482 45332 36484
rect 45276 36430 45278 36482
rect 45278 36430 45330 36482
rect 45330 36430 45332 36482
rect 45276 36428 45332 36430
rect 44940 36204 44996 36260
rect 44268 35644 44324 35700
rect 44716 35698 44772 35700
rect 44716 35646 44718 35698
rect 44718 35646 44770 35698
rect 44770 35646 44772 35698
rect 44716 35644 44772 35646
rect 45164 36092 45220 36148
rect 45500 36204 45556 36260
rect 45836 37266 45892 37268
rect 45836 37214 45838 37266
rect 45838 37214 45890 37266
rect 45890 37214 45892 37266
rect 45836 37212 45892 37214
rect 46060 36988 46116 37044
rect 46172 36876 46228 36932
rect 45164 35868 45220 35924
rect 45724 35698 45780 35700
rect 45724 35646 45726 35698
rect 45726 35646 45778 35698
rect 45778 35646 45780 35698
rect 45724 35644 45780 35646
rect 44380 35196 44436 35252
rect 43932 34690 43988 34692
rect 43932 34638 43934 34690
rect 43934 34638 43986 34690
rect 43986 34638 43988 34690
rect 43932 34636 43988 34638
rect 43820 34242 43876 34244
rect 43820 34190 43822 34242
rect 43822 34190 43874 34242
rect 43874 34190 43876 34242
rect 43820 34188 43876 34190
rect 43932 33516 43988 33572
rect 45948 35922 46004 35924
rect 45948 35870 45950 35922
rect 45950 35870 46002 35922
rect 46002 35870 46004 35922
rect 45948 35868 46004 35870
rect 45276 35196 45332 35252
rect 47404 42754 47460 42756
rect 47404 42702 47406 42754
rect 47406 42702 47458 42754
rect 47458 42702 47460 42754
rect 47404 42700 47460 42702
rect 52332 44994 52388 44996
rect 52332 44942 52334 44994
rect 52334 44942 52386 44994
rect 52386 44942 52388 44994
rect 52332 44940 52388 44942
rect 49084 44044 49140 44100
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 48188 42700 48244 42756
rect 48748 43372 48804 43428
rect 49084 42588 49140 42644
rect 49756 42588 49812 42644
rect 48748 41804 48804 41860
rect 48188 40572 48244 40628
rect 47740 40290 47796 40292
rect 47740 40238 47742 40290
rect 47742 40238 47794 40290
rect 47794 40238 47796 40290
rect 47740 40236 47796 40238
rect 47292 39788 47348 39844
rect 47852 39788 47908 39844
rect 47852 39228 47908 39284
rect 47964 39618 48020 39620
rect 47964 39566 47966 39618
rect 47966 39566 48018 39618
rect 48018 39566 48020 39618
rect 47964 39564 48020 39566
rect 46956 38892 47012 38948
rect 47740 39004 47796 39060
rect 47852 38946 47908 38948
rect 47852 38894 47854 38946
rect 47854 38894 47906 38946
rect 47906 38894 47908 38946
rect 47852 38892 47908 38894
rect 46620 38834 46676 38836
rect 46620 38782 46622 38834
rect 46622 38782 46674 38834
rect 46674 38782 46676 38834
rect 46620 38780 46676 38782
rect 46396 36764 46452 36820
rect 46620 37212 46676 37268
rect 46284 36652 46340 36708
rect 45164 34188 45220 34244
rect 44716 33740 44772 33796
rect 45724 34802 45780 34804
rect 45724 34750 45726 34802
rect 45726 34750 45778 34802
rect 45778 34750 45780 34802
rect 45724 34748 45780 34750
rect 47404 37100 47460 37156
rect 46844 36988 46900 37044
rect 47180 36428 47236 36484
rect 45500 33740 45556 33796
rect 47068 36316 47124 36372
rect 47068 35868 47124 35924
rect 46396 34802 46452 34804
rect 46396 34750 46398 34802
rect 46398 34750 46450 34802
rect 46450 34750 46452 34802
rect 46396 34748 46452 34750
rect 47068 35308 47124 35364
rect 47292 35420 47348 35476
rect 43260 31276 43316 31332
rect 42364 30156 42420 30212
rect 43484 31276 43540 31332
rect 43372 30044 43428 30100
rect 42252 29372 42308 29428
rect 43260 29986 43316 29988
rect 43260 29934 43262 29986
rect 43262 29934 43314 29986
rect 43314 29934 43316 29986
rect 43260 29932 43316 29934
rect 42588 28588 42644 28644
rect 41244 26850 41300 26852
rect 41244 26798 41246 26850
rect 41246 26798 41298 26850
rect 41298 26798 41300 26850
rect 41244 26796 41300 26798
rect 41132 26572 41188 26628
rect 40796 25506 40852 25508
rect 40796 25454 40798 25506
rect 40798 25454 40850 25506
rect 40850 25454 40852 25506
rect 40796 25452 40852 25454
rect 40908 25116 40964 25172
rect 42140 27244 42196 27300
rect 41916 27074 41972 27076
rect 41916 27022 41918 27074
rect 41918 27022 41970 27074
rect 41970 27022 41972 27074
rect 41916 27020 41972 27022
rect 41356 26236 41412 26292
rect 41244 25340 41300 25396
rect 41356 25228 41412 25284
rect 41132 25004 41188 25060
rect 41244 24780 41300 24836
rect 40684 23660 40740 23716
rect 40796 24668 40852 24724
rect 41020 24722 41076 24724
rect 41020 24670 41022 24722
rect 41022 24670 41074 24722
rect 41074 24670 41076 24722
rect 41020 24668 41076 24670
rect 40796 23324 40852 23380
rect 40908 23772 40964 23828
rect 40684 22370 40740 22372
rect 40684 22318 40686 22370
rect 40686 22318 40738 22370
rect 40738 22318 40740 22370
rect 40684 22316 40740 22318
rect 41132 22652 41188 22708
rect 41916 26290 41972 26292
rect 41916 26238 41918 26290
rect 41918 26238 41970 26290
rect 41970 26238 41972 26290
rect 41916 26236 41972 26238
rect 41692 25452 41748 25508
rect 42476 28418 42532 28420
rect 42476 28366 42478 28418
rect 42478 28366 42530 28418
rect 42530 28366 42532 28418
rect 42476 28364 42532 28366
rect 43820 32732 43876 32788
rect 43708 32562 43764 32564
rect 43708 32510 43710 32562
rect 43710 32510 43762 32562
rect 43762 32510 43764 32562
rect 43708 32508 43764 32510
rect 43820 32450 43876 32452
rect 43820 32398 43822 32450
rect 43822 32398 43874 32450
rect 43874 32398 43876 32450
rect 43820 32396 43876 32398
rect 43932 31612 43988 31668
rect 44044 31724 44100 31780
rect 44268 31724 44324 31780
rect 44156 31106 44212 31108
rect 44156 31054 44158 31106
rect 44158 31054 44210 31106
rect 44210 31054 44212 31106
rect 44156 31052 44212 31054
rect 43484 29372 43540 29428
rect 43372 28754 43428 28756
rect 43372 28702 43374 28754
rect 43374 28702 43426 28754
rect 43426 28702 43428 28754
rect 43372 28700 43428 28702
rect 43596 28924 43652 28980
rect 44492 29314 44548 29316
rect 44492 29262 44494 29314
rect 44494 29262 44546 29314
rect 44546 29262 44548 29314
rect 44492 29260 44548 29262
rect 43820 28812 43876 28868
rect 45388 32956 45444 33012
rect 44828 32284 44884 32340
rect 44716 30940 44772 30996
rect 44940 31890 44996 31892
rect 44940 31838 44942 31890
rect 44942 31838 44994 31890
rect 44994 31838 44996 31890
rect 44940 31836 44996 31838
rect 45388 31276 45444 31332
rect 44940 31164 44996 31220
rect 45276 30994 45332 30996
rect 45276 30942 45278 30994
rect 45278 30942 45330 30994
rect 45330 30942 45332 30994
rect 45276 30940 45332 30942
rect 45500 31218 45556 31220
rect 45500 31166 45502 31218
rect 45502 31166 45554 31218
rect 45554 31166 45556 31218
rect 45500 31164 45556 31166
rect 45836 33516 45892 33572
rect 46508 33292 46564 33348
rect 46396 32786 46452 32788
rect 46396 32734 46398 32786
rect 46398 32734 46450 32786
rect 46450 32734 46452 32786
rect 46396 32732 46452 32734
rect 47068 33628 47124 33684
rect 47180 33292 47236 33348
rect 47180 33122 47236 33124
rect 47180 33070 47182 33122
rect 47182 33070 47234 33122
rect 47234 33070 47236 33122
rect 47180 33068 47236 33070
rect 46844 32956 46900 33012
rect 47628 36594 47684 36596
rect 47628 36542 47630 36594
rect 47630 36542 47682 36594
rect 47682 36542 47684 36594
rect 47628 36540 47684 36542
rect 47516 36370 47572 36372
rect 47516 36318 47518 36370
rect 47518 36318 47570 36370
rect 47570 36318 47572 36370
rect 47516 36316 47572 36318
rect 47740 36204 47796 36260
rect 48860 41020 48916 41076
rect 51100 43426 51156 43428
rect 51100 43374 51102 43426
rect 51102 43374 51154 43426
rect 51154 43374 51156 43426
rect 51100 43372 51156 43374
rect 51324 43148 51380 43204
rect 51660 43314 51716 43316
rect 51660 43262 51662 43314
rect 51662 43262 51714 43314
rect 51714 43262 51716 43314
rect 51660 43260 51716 43262
rect 50316 42476 50372 42532
rect 49420 41692 49476 41748
rect 49980 41410 50036 41412
rect 49980 41358 49982 41410
rect 49982 41358 50034 41410
rect 50034 41358 50036 41410
rect 49980 41356 50036 41358
rect 49980 41074 50036 41076
rect 49980 41022 49982 41074
rect 49982 41022 50034 41074
rect 50034 41022 50036 41074
rect 49980 41020 50036 41022
rect 50428 42700 50484 42756
rect 50764 42476 50820 42532
rect 50988 42476 51044 42532
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 48748 38892 48804 38948
rect 49196 40626 49252 40628
rect 49196 40574 49198 40626
rect 49198 40574 49250 40626
rect 49250 40574 49252 40626
rect 49196 40572 49252 40574
rect 49420 40460 49476 40516
rect 48972 39564 49028 39620
rect 48300 38780 48356 38836
rect 48300 38556 48356 38612
rect 49084 40236 49140 40292
rect 49084 39506 49140 39508
rect 49084 39454 49086 39506
rect 49086 39454 49138 39506
rect 49138 39454 49140 39506
rect 49084 39452 49140 39454
rect 48188 37884 48244 37940
rect 48076 36092 48132 36148
rect 47516 35308 47572 35364
rect 47628 34748 47684 34804
rect 47516 32732 47572 32788
rect 46284 32338 46340 32340
rect 46284 32286 46286 32338
rect 46286 32286 46338 32338
rect 46338 32286 46340 32338
rect 46284 32284 46340 32286
rect 46284 31836 46340 31892
rect 45052 30770 45108 30772
rect 45052 30718 45054 30770
rect 45054 30718 45106 30770
rect 45106 30718 45108 30770
rect 45052 30716 45108 30718
rect 44716 29372 44772 29428
rect 44268 29036 44324 29092
rect 44044 28700 44100 28756
rect 43036 27468 43092 27524
rect 42924 27244 42980 27300
rect 42252 27020 42308 27076
rect 42812 27074 42868 27076
rect 42812 27022 42814 27074
rect 42814 27022 42866 27074
rect 42866 27022 42868 27074
rect 42812 27020 42868 27022
rect 42476 25788 42532 25844
rect 42588 26572 42644 26628
rect 42252 25506 42308 25508
rect 42252 25454 42254 25506
rect 42254 25454 42306 25506
rect 42306 25454 42308 25506
rect 42252 25452 42308 25454
rect 42028 25228 42084 25284
rect 42476 25228 42532 25284
rect 42140 25116 42196 25172
rect 41804 24108 41860 24164
rect 41356 23772 41412 23828
rect 41692 23548 41748 23604
rect 42028 23772 42084 23828
rect 41804 23660 41860 23716
rect 41244 23212 41300 23268
rect 42252 23212 42308 23268
rect 42140 23042 42196 23044
rect 42140 22990 42142 23042
rect 42142 22990 42194 23042
rect 42194 22990 42196 23042
rect 42140 22988 42196 22990
rect 42028 22652 42084 22708
rect 41244 22540 41300 22596
rect 42028 22482 42084 22484
rect 42028 22430 42030 22482
rect 42030 22430 42082 22482
rect 42082 22430 42084 22482
rect 42028 22428 42084 22430
rect 40236 22204 40292 22260
rect 41020 22092 41076 22148
rect 40124 21980 40180 22036
rect 39900 21644 39956 21700
rect 40236 21474 40292 21476
rect 40236 21422 40238 21474
rect 40238 21422 40290 21474
rect 40290 21422 40292 21474
rect 40236 21420 40292 21422
rect 37100 19906 37156 19908
rect 37100 19854 37102 19906
rect 37102 19854 37154 19906
rect 37154 19854 37156 19906
rect 37100 19852 37156 19854
rect 39116 20524 39172 20580
rect 41244 21532 41300 21588
rect 41804 21420 41860 21476
rect 42252 22092 42308 22148
rect 43260 28252 43316 28308
rect 43596 27468 43652 27524
rect 44268 28476 44324 28532
rect 44828 28700 44884 28756
rect 45164 29426 45220 29428
rect 45164 29374 45166 29426
rect 45166 29374 45218 29426
rect 45218 29374 45220 29426
rect 45164 29372 45220 29374
rect 45164 29148 45220 29204
rect 44940 28028 44996 28084
rect 44044 27020 44100 27076
rect 43260 26908 43316 26964
rect 43484 26908 43540 26964
rect 43932 26796 43988 26852
rect 43484 25788 43540 25844
rect 42812 25506 42868 25508
rect 42812 25454 42814 25506
rect 42814 25454 42866 25506
rect 42866 25454 42868 25506
rect 42812 25452 42868 25454
rect 42700 24668 42756 24724
rect 42812 23324 42868 23380
rect 42476 22876 42532 22932
rect 42588 22428 42644 22484
rect 42812 22092 42868 22148
rect 42476 21980 42532 22036
rect 43036 23100 43092 23156
rect 43596 25564 43652 25620
rect 43148 22316 43204 22372
rect 43484 23548 43540 23604
rect 43372 22258 43428 22260
rect 43372 22206 43374 22258
rect 43374 22206 43426 22258
rect 43426 22206 43428 22258
rect 43372 22204 43428 22206
rect 43036 21586 43092 21588
rect 43036 21534 43038 21586
rect 43038 21534 43090 21586
rect 43090 21534 43092 21586
rect 43036 21532 43092 21534
rect 43708 25452 43764 25508
rect 45612 30716 45668 30772
rect 45612 30044 45668 30100
rect 45724 29820 45780 29876
rect 45836 29708 45892 29764
rect 46060 29596 46116 29652
rect 45836 29484 45892 29540
rect 45724 29372 45780 29428
rect 45388 28700 45444 28756
rect 45500 28812 45556 28868
rect 45052 27298 45108 27300
rect 45052 27246 45054 27298
rect 45054 27246 45106 27298
rect 45106 27246 45108 27298
rect 45052 27244 45108 27246
rect 45276 27132 45332 27188
rect 45276 26460 45332 26516
rect 44044 25340 44100 25396
rect 44156 25228 44212 25284
rect 44268 24556 44324 24612
rect 45388 26236 45444 26292
rect 45388 25788 45444 25844
rect 44940 25506 44996 25508
rect 44940 25454 44942 25506
rect 44942 25454 44994 25506
rect 44994 25454 44996 25506
rect 44940 25452 44996 25454
rect 44940 24556 44996 24612
rect 43820 23154 43876 23156
rect 43820 23102 43822 23154
rect 43822 23102 43874 23154
rect 43874 23102 43876 23154
rect 43820 23100 43876 23102
rect 45164 23938 45220 23940
rect 45164 23886 45166 23938
rect 45166 23886 45218 23938
rect 45218 23886 45220 23938
rect 45164 23884 45220 23886
rect 46172 28588 46228 28644
rect 46508 30994 46564 30996
rect 46508 30942 46510 30994
rect 46510 30942 46562 30994
rect 46562 30942 46564 30994
rect 46508 30940 46564 30942
rect 46508 30380 46564 30436
rect 46396 30210 46452 30212
rect 46396 30158 46398 30210
rect 46398 30158 46450 30210
rect 46450 30158 46452 30210
rect 46396 30156 46452 30158
rect 46956 32674 47012 32676
rect 46956 32622 46958 32674
rect 46958 32622 47010 32674
rect 47010 32622 47012 32674
rect 46956 32620 47012 32622
rect 47740 32508 47796 32564
rect 47852 35644 47908 35700
rect 46732 32060 46788 32116
rect 46844 31388 46900 31444
rect 47628 31554 47684 31556
rect 47628 31502 47630 31554
rect 47630 31502 47682 31554
rect 47682 31502 47684 31554
rect 47628 31500 47684 31502
rect 47180 30940 47236 30996
rect 46732 30882 46788 30884
rect 46732 30830 46734 30882
rect 46734 30830 46786 30882
rect 46786 30830 46788 30882
rect 46732 30828 46788 30830
rect 46844 30268 46900 30324
rect 47740 30322 47796 30324
rect 47740 30270 47742 30322
rect 47742 30270 47794 30322
rect 47794 30270 47796 30322
rect 47740 30268 47796 30270
rect 46956 30156 47012 30212
rect 46956 29650 47012 29652
rect 46956 29598 46958 29650
rect 46958 29598 47010 29650
rect 47010 29598 47012 29650
rect 46956 29596 47012 29598
rect 48188 34242 48244 34244
rect 48188 34190 48190 34242
rect 48190 34190 48242 34242
rect 48242 34190 48244 34242
rect 48188 34188 48244 34190
rect 47964 32844 48020 32900
rect 48860 36876 48916 36932
rect 48972 36540 49028 36596
rect 48748 36428 48804 36484
rect 49420 39788 49476 39844
rect 49756 40402 49812 40404
rect 49756 40350 49758 40402
rect 49758 40350 49810 40402
rect 49810 40350 49812 40402
rect 49756 40348 49812 40350
rect 49644 40290 49700 40292
rect 49644 40238 49646 40290
rect 49646 40238 49698 40290
rect 49698 40238 49700 40290
rect 49644 40236 49700 40238
rect 50764 40962 50820 40964
rect 50764 40910 50766 40962
rect 50766 40910 50818 40962
rect 50818 40910 50820 40962
rect 50764 40908 50820 40910
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 53788 43260 53844 43316
rect 51660 42642 51716 42644
rect 51660 42590 51662 42642
rect 51662 42590 51714 42642
rect 51714 42590 51716 42642
rect 51660 42588 51716 42590
rect 51884 42028 51940 42084
rect 51324 41356 51380 41412
rect 50204 40348 50260 40404
rect 50092 40236 50148 40292
rect 50316 39900 50372 39956
rect 50204 39788 50260 39844
rect 49532 39676 49588 39732
rect 49308 39618 49364 39620
rect 49308 39566 49310 39618
rect 49310 39566 49362 39618
rect 49362 39566 49364 39618
rect 49308 39564 49364 39566
rect 49756 39618 49812 39620
rect 49756 39566 49758 39618
rect 49758 39566 49810 39618
rect 49810 39566 49812 39618
rect 49756 39564 49812 39566
rect 49644 39506 49700 39508
rect 49644 39454 49646 39506
rect 49646 39454 49698 39506
rect 49698 39454 49700 39506
rect 49644 39452 49700 39454
rect 49644 39004 49700 39060
rect 49756 38946 49812 38948
rect 49756 38894 49758 38946
rect 49758 38894 49810 38946
rect 49810 38894 49812 38946
rect 49756 38892 49812 38894
rect 48748 35474 48804 35476
rect 48748 35422 48750 35474
rect 48750 35422 48802 35474
rect 48802 35422 48804 35474
rect 48748 35420 48804 35422
rect 48748 34748 48804 34804
rect 48524 34300 48580 34356
rect 48748 34130 48804 34132
rect 48748 34078 48750 34130
rect 48750 34078 48802 34130
rect 48802 34078 48804 34130
rect 48748 34076 48804 34078
rect 50428 40124 50484 40180
rect 50988 40514 51044 40516
rect 50988 40462 50990 40514
rect 50990 40462 51042 40514
rect 51042 40462 51044 40514
rect 50988 40460 51044 40462
rect 53004 42082 53060 42084
rect 53004 42030 53006 42082
rect 53006 42030 53058 42082
rect 53058 42030 53060 42082
rect 53004 42028 53060 42030
rect 51996 41692 52052 41748
rect 52220 41916 52276 41972
rect 51884 40908 51940 40964
rect 53676 41970 53732 41972
rect 53676 41918 53678 41970
rect 53678 41918 53730 41970
rect 53730 41918 53732 41970
rect 53676 41916 53732 41918
rect 52780 41692 52836 41748
rect 52556 40626 52612 40628
rect 52556 40574 52558 40626
rect 52558 40574 52610 40626
rect 52610 40574 52612 40626
rect 52556 40572 52612 40574
rect 51324 40514 51380 40516
rect 51324 40462 51326 40514
rect 51326 40462 51378 40514
rect 51378 40462 51380 40514
rect 51324 40460 51380 40462
rect 51884 40514 51940 40516
rect 51884 40462 51886 40514
rect 51886 40462 51938 40514
rect 51938 40462 51940 40514
rect 51884 40460 51940 40462
rect 50764 40402 50820 40404
rect 50764 40350 50766 40402
rect 50766 40350 50818 40402
rect 50818 40350 50820 40402
rect 50764 40348 50820 40350
rect 51660 40348 51716 40404
rect 50876 40290 50932 40292
rect 50876 40238 50878 40290
rect 50878 40238 50930 40290
rect 50930 40238 50932 40290
rect 50876 40236 50932 40238
rect 50652 40124 50708 40180
rect 50988 40012 51044 40068
rect 50652 39788 50708 39844
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50428 39004 50484 39060
rect 50316 38780 50372 38836
rect 51660 38668 51716 38724
rect 53340 38722 53396 38724
rect 53340 38670 53342 38722
rect 53342 38670 53394 38722
rect 53394 38670 53396 38722
rect 53340 38668 53396 38670
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50428 36876 50484 36932
rect 49868 36652 49924 36708
rect 50204 36540 50260 36596
rect 50204 36092 50260 36148
rect 49420 35644 49476 35700
rect 48972 35196 49028 35252
rect 48972 34636 49028 34692
rect 49308 34914 49364 34916
rect 49308 34862 49310 34914
rect 49310 34862 49362 34914
rect 49362 34862 49364 34914
rect 49308 34860 49364 34862
rect 49084 34524 49140 34580
rect 49420 34748 49476 34804
rect 48188 31666 48244 31668
rect 48188 31614 48190 31666
rect 48190 31614 48242 31666
rect 48242 31614 48244 31666
rect 48188 31612 48244 31614
rect 48412 31666 48468 31668
rect 48412 31614 48414 31666
rect 48414 31614 48466 31666
rect 48466 31614 48468 31666
rect 48412 31612 48468 31614
rect 48188 31052 48244 31108
rect 47964 30268 48020 30324
rect 47292 29820 47348 29876
rect 46620 29426 46676 29428
rect 46620 29374 46622 29426
rect 46622 29374 46674 29426
rect 46674 29374 46676 29426
rect 46620 29372 46676 29374
rect 47068 29426 47124 29428
rect 47068 29374 47070 29426
rect 47070 29374 47122 29426
rect 47122 29374 47124 29426
rect 47068 29372 47124 29374
rect 46396 29148 46452 29204
rect 47180 29148 47236 29204
rect 46620 28812 46676 28868
rect 46396 28700 46452 28756
rect 45836 27244 45892 27300
rect 45724 27074 45780 27076
rect 45724 27022 45726 27074
rect 45726 27022 45778 27074
rect 45778 27022 45780 27074
rect 45724 27020 45780 27022
rect 46060 26348 46116 26404
rect 45836 25564 45892 25620
rect 45948 26124 46004 26180
rect 46172 25788 46228 25844
rect 45724 25340 45780 25396
rect 45948 24556 46004 24612
rect 45612 24108 45668 24164
rect 47404 29650 47460 29652
rect 47404 29598 47406 29650
rect 47406 29598 47458 29650
rect 47458 29598 47460 29650
rect 47404 29596 47460 29598
rect 47404 29260 47460 29316
rect 46732 27916 46788 27972
rect 46620 27020 46676 27076
rect 46732 26348 46788 26404
rect 46956 28418 47012 28420
rect 46956 28366 46958 28418
rect 46958 28366 47010 28418
rect 47010 28366 47012 28418
rect 46956 28364 47012 28366
rect 46844 26236 46900 26292
rect 46956 25618 47012 25620
rect 46956 25566 46958 25618
rect 46958 25566 47010 25618
rect 47010 25566 47012 25618
rect 46956 25564 47012 25566
rect 47292 28530 47348 28532
rect 47292 28478 47294 28530
rect 47294 28478 47346 28530
rect 47346 28478 47348 28530
rect 47292 28476 47348 28478
rect 48076 29986 48132 29988
rect 48076 29934 48078 29986
rect 48078 29934 48130 29986
rect 48130 29934 48132 29986
rect 48076 29932 48132 29934
rect 48860 31276 48916 31332
rect 48748 30156 48804 30212
rect 49084 32844 49140 32900
rect 49420 33964 49476 34020
rect 49196 33068 49252 33124
rect 49980 35644 50036 35700
rect 49644 34188 49700 34244
rect 49756 34524 49812 34580
rect 50092 34748 50148 34804
rect 50204 34242 50260 34244
rect 50204 34190 50206 34242
rect 50206 34190 50258 34242
rect 50258 34190 50260 34242
rect 50204 34188 50260 34190
rect 50204 33852 50260 33908
rect 49196 32732 49252 32788
rect 49532 32508 49588 32564
rect 49084 31500 49140 31556
rect 49420 31218 49476 31220
rect 49420 31166 49422 31218
rect 49422 31166 49474 31218
rect 49474 31166 49476 31218
rect 49420 31164 49476 31166
rect 49420 30828 49476 30884
rect 49196 30380 49252 30436
rect 49756 32562 49812 32564
rect 49756 32510 49758 32562
rect 49758 32510 49810 32562
rect 49810 32510 49812 32562
rect 49756 32508 49812 32510
rect 49756 32284 49812 32340
rect 49756 31276 49812 31332
rect 50204 32508 50260 32564
rect 50988 37884 51044 37940
rect 51100 37826 51156 37828
rect 51100 37774 51102 37826
rect 51102 37774 51154 37826
rect 51154 37774 51156 37826
rect 51100 37772 51156 37774
rect 51100 37212 51156 37268
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50428 34860 50484 34916
rect 50764 35868 50820 35924
rect 50764 35698 50820 35700
rect 50764 35646 50766 35698
rect 50766 35646 50818 35698
rect 50818 35646 50820 35698
rect 50764 35644 50820 35646
rect 51772 38050 51828 38052
rect 51772 37998 51774 38050
rect 51774 37998 51826 38050
rect 51826 37998 51828 38050
rect 51772 37996 51828 37998
rect 52780 37996 52836 38052
rect 52556 37884 52612 37940
rect 52556 36876 52612 36932
rect 51660 36764 51716 36820
rect 52332 36764 52388 36820
rect 52108 36258 52164 36260
rect 52108 36206 52110 36258
rect 52110 36206 52162 36258
rect 52162 36206 52164 36258
rect 52108 36204 52164 36206
rect 51212 35868 51268 35924
rect 51548 35308 51604 35364
rect 51100 34748 51156 34804
rect 51772 34860 51828 34916
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 51660 34300 51716 34356
rect 50652 34242 50708 34244
rect 50652 34190 50654 34242
rect 50654 34190 50706 34242
rect 50706 34190 50708 34242
rect 50652 34188 50708 34190
rect 50428 34076 50484 34132
rect 51100 34076 51156 34132
rect 50988 33740 51044 33796
rect 50876 33346 50932 33348
rect 50876 33294 50878 33346
rect 50878 33294 50930 33346
rect 50930 33294 50932 33346
rect 50876 33292 50932 33294
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50764 32562 50820 32564
rect 50764 32510 50766 32562
rect 50766 32510 50818 32562
rect 50818 32510 50820 32562
rect 50764 32508 50820 32510
rect 50316 32284 50372 32340
rect 52668 36316 52724 36372
rect 52332 34860 52388 34916
rect 52668 35084 52724 35140
rect 53564 37996 53620 38052
rect 54572 38050 54628 38052
rect 54572 37998 54574 38050
rect 54574 37998 54626 38050
rect 54626 37998 54628 38050
rect 54572 37996 54628 37998
rect 52892 36652 52948 36708
rect 52892 35868 52948 35924
rect 52892 35196 52948 35252
rect 51660 33964 51716 34020
rect 51212 33906 51268 33908
rect 51212 33854 51214 33906
rect 51214 33854 51266 33906
rect 51266 33854 51268 33906
rect 51212 33852 51268 33854
rect 51212 33628 51268 33684
rect 52108 33234 52164 33236
rect 52108 33182 52110 33234
rect 52110 33182 52162 33234
rect 52162 33182 52164 33234
rect 52108 33180 52164 33182
rect 53340 35196 53396 35252
rect 54124 37266 54180 37268
rect 54124 37214 54126 37266
rect 54126 37214 54178 37266
rect 54178 37214 54180 37266
rect 54124 37212 54180 37214
rect 53564 36988 53620 37044
rect 53228 34802 53284 34804
rect 53228 34750 53230 34802
rect 53230 34750 53282 34802
rect 53282 34750 53284 34802
rect 53228 34748 53284 34750
rect 53452 34802 53508 34804
rect 53452 34750 53454 34802
rect 53454 34750 53506 34802
rect 53506 34750 53508 34802
rect 53452 34748 53508 34750
rect 54796 37042 54852 37044
rect 54796 36990 54798 37042
rect 54798 36990 54850 37042
rect 54850 36990 54852 37042
rect 54796 36988 54852 36990
rect 54572 36652 54628 36708
rect 54684 36876 54740 36932
rect 54012 36428 54068 36484
rect 54572 36428 54628 36484
rect 54124 36316 54180 36372
rect 54460 36316 54516 36372
rect 54236 36204 54292 36260
rect 53676 35196 53732 35252
rect 53676 34300 53732 34356
rect 53564 33180 53620 33236
rect 52220 32786 52276 32788
rect 52220 32734 52222 32786
rect 52222 32734 52274 32786
rect 52274 32734 52276 32786
rect 52220 32732 52276 32734
rect 51660 32674 51716 32676
rect 51660 32622 51662 32674
rect 51662 32622 51714 32674
rect 51714 32622 51716 32674
rect 51660 32620 51716 32622
rect 51772 32562 51828 32564
rect 51772 32510 51774 32562
rect 51774 32510 51826 32562
rect 51826 32510 51828 32562
rect 51772 32508 51828 32510
rect 50988 32172 51044 32228
rect 51324 31948 51380 32004
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50204 30828 50260 30884
rect 51996 31948 52052 32004
rect 51436 31554 51492 31556
rect 51436 31502 51438 31554
rect 51438 31502 51490 31554
rect 51490 31502 51492 31554
rect 51436 31500 51492 31502
rect 48524 29986 48580 29988
rect 48524 29934 48526 29986
rect 48526 29934 48578 29986
rect 48578 29934 48580 29986
rect 48524 29932 48580 29934
rect 48300 29260 48356 29316
rect 49420 29986 49476 29988
rect 49420 29934 49422 29986
rect 49422 29934 49474 29986
rect 49474 29934 49476 29986
rect 49420 29932 49476 29934
rect 49644 29986 49700 29988
rect 49644 29934 49646 29986
rect 49646 29934 49698 29986
rect 49698 29934 49700 29986
rect 49644 29932 49700 29934
rect 47404 27186 47460 27188
rect 47404 27134 47406 27186
rect 47406 27134 47458 27186
rect 47458 27134 47460 27186
rect 47404 27132 47460 27134
rect 49868 29596 49924 29652
rect 47852 27858 47908 27860
rect 47852 27806 47854 27858
rect 47854 27806 47906 27858
rect 47906 27806 47908 27858
rect 47852 27804 47908 27806
rect 48860 28252 48916 28308
rect 48188 27132 48244 27188
rect 48748 27074 48804 27076
rect 48748 27022 48750 27074
rect 48750 27022 48802 27074
rect 48802 27022 48804 27074
rect 48748 27020 48804 27022
rect 49196 27580 49252 27636
rect 48524 26850 48580 26852
rect 48524 26798 48526 26850
rect 48526 26798 48578 26850
rect 48578 26798 48580 26850
rect 48524 26796 48580 26798
rect 47628 26402 47684 26404
rect 47628 26350 47630 26402
rect 47630 26350 47682 26402
rect 47682 26350 47684 26402
rect 47628 26348 47684 26350
rect 47516 25788 47572 25844
rect 47516 25564 47572 25620
rect 47292 25452 47348 25508
rect 46508 24722 46564 24724
rect 46508 24670 46510 24722
rect 46510 24670 46562 24722
rect 46562 24670 46564 24722
rect 46508 24668 46564 24670
rect 45388 23660 45444 23716
rect 45388 23154 45444 23156
rect 45388 23102 45390 23154
rect 45390 23102 45442 23154
rect 45442 23102 45444 23154
rect 45388 23100 45444 23102
rect 44828 22652 44884 22708
rect 46396 23996 46452 24052
rect 46508 23826 46564 23828
rect 46508 23774 46510 23826
rect 46510 23774 46562 23826
rect 46562 23774 46564 23826
rect 46508 23772 46564 23774
rect 46060 23266 46116 23268
rect 46060 23214 46062 23266
rect 46062 23214 46114 23266
rect 46114 23214 46116 23266
rect 46060 23212 46116 23214
rect 46060 22540 46116 22596
rect 44268 22204 44324 22260
rect 45276 22258 45332 22260
rect 45276 22206 45278 22258
rect 45278 22206 45330 22258
rect 45330 22206 45332 22258
rect 45276 22204 45332 22206
rect 43932 21474 43988 21476
rect 43932 21422 43934 21474
rect 43934 21422 43986 21474
rect 43986 21422 43988 21474
rect 43932 21420 43988 21422
rect 44044 22092 44100 22148
rect 41580 20578 41636 20580
rect 41580 20526 41582 20578
rect 41582 20526 41634 20578
rect 41634 20526 41636 20578
rect 41580 20524 41636 20526
rect 45500 22258 45556 22260
rect 45500 22206 45502 22258
rect 45502 22206 45554 22258
rect 45554 22206 45556 22258
rect 45500 22204 45556 22206
rect 45388 22092 45444 22148
rect 44268 21308 44324 21364
rect 44940 20860 44996 20916
rect 46060 22370 46116 22372
rect 46060 22318 46062 22370
rect 46062 22318 46114 22370
rect 46114 22318 46116 22370
rect 46060 22316 46116 22318
rect 46060 22092 46116 22148
rect 46284 22876 46340 22932
rect 46172 21644 46228 21700
rect 46732 24220 46788 24276
rect 47180 25004 47236 25060
rect 47180 24220 47236 24276
rect 47068 23996 47124 24052
rect 47292 23996 47348 24052
rect 46508 22482 46564 22484
rect 46508 22430 46510 22482
rect 46510 22430 46562 22482
rect 46562 22430 46564 22482
rect 46508 22428 46564 22430
rect 47068 23436 47124 23492
rect 47628 24220 47684 24276
rect 47740 25228 47796 25284
rect 47964 24610 48020 24612
rect 47964 24558 47966 24610
rect 47966 24558 48018 24610
rect 48018 24558 48020 24610
rect 47964 24556 48020 24558
rect 48636 26460 48692 26516
rect 48860 26514 48916 26516
rect 48860 26462 48862 26514
rect 48862 26462 48914 26514
rect 48914 26462 48916 26514
rect 48860 26460 48916 26462
rect 48972 26236 49028 26292
rect 48636 24556 48692 24612
rect 48188 24444 48244 24500
rect 47852 24332 47908 24388
rect 47404 23884 47460 23940
rect 47628 23436 47684 23492
rect 47068 22428 47124 22484
rect 47292 21644 47348 21700
rect 47964 23436 48020 23492
rect 47516 21980 47572 22036
rect 47628 22316 47684 22372
rect 47852 22428 47908 22484
rect 49644 29260 49700 29316
rect 49532 28252 49588 28308
rect 49756 29148 49812 29204
rect 50204 29820 50260 29876
rect 49980 28476 50036 28532
rect 49980 27580 50036 27636
rect 49868 26684 49924 26740
rect 49196 25004 49252 25060
rect 49084 24668 49140 24724
rect 49420 25004 49476 25060
rect 49084 24444 49140 24500
rect 48972 23772 49028 23828
rect 48188 23548 48244 23604
rect 47964 22204 48020 22260
rect 47740 21532 47796 21588
rect 46844 20860 46900 20916
rect 47180 20860 47236 20916
rect 47852 21756 47908 21812
rect 48524 23436 48580 23492
rect 48972 23436 49028 23492
rect 49532 24946 49588 24948
rect 49532 24894 49534 24946
rect 49534 24894 49586 24946
rect 49586 24894 49588 24946
rect 49532 24892 49588 24894
rect 49532 24722 49588 24724
rect 49532 24670 49534 24722
rect 49534 24670 49586 24722
rect 49586 24670 49588 24722
rect 49532 24668 49588 24670
rect 49196 24220 49252 24276
rect 49420 23884 49476 23940
rect 49308 23772 49364 23828
rect 49644 23772 49700 23828
rect 49532 23548 49588 23604
rect 48636 23212 48692 23268
rect 49308 23154 49364 23156
rect 49308 23102 49310 23154
rect 49310 23102 49362 23154
rect 49362 23102 49364 23154
rect 49308 23100 49364 23102
rect 49084 22876 49140 22932
rect 48860 22428 48916 22484
rect 48412 22370 48468 22372
rect 48412 22318 48414 22370
rect 48414 22318 48466 22370
rect 48466 22318 48468 22370
rect 48412 22316 48468 22318
rect 49420 22258 49476 22260
rect 49420 22206 49422 22258
rect 49422 22206 49474 22258
rect 49474 22206 49476 22258
rect 49420 22204 49476 22206
rect 48636 22146 48692 22148
rect 48636 22094 48638 22146
rect 48638 22094 48690 22146
rect 48690 22094 48692 22146
rect 48636 22092 48692 22094
rect 48748 21980 48804 22036
rect 49644 23324 49700 23380
rect 50988 30604 51044 30660
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50428 28028 50484 28084
rect 50428 27580 50484 27636
rect 50652 28028 50708 28084
rect 50764 27356 50820 27412
rect 50316 26348 50372 26404
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 51660 31836 51716 31892
rect 51548 30044 51604 30100
rect 51212 28812 51268 28868
rect 51436 29932 51492 29988
rect 52668 31778 52724 31780
rect 52668 31726 52670 31778
rect 52670 31726 52722 31778
rect 52722 31726 52724 31778
rect 52668 31724 52724 31726
rect 51884 31666 51940 31668
rect 51884 31614 51886 31666
rect 51886 31614 51938 31666
rect 51938 31614 51940 31666
rect 51884 31612 51940 31614
rect 51884 31106 51940 31108
rect 51884 31054 51886 31106
rect 51886 31054 51938 31106
rect 51938 31054 51940 31106
rect 51884 31052 51940 31054
rect 52108 31106 52164 31108
rect 52108 31054 52110 31106
rect 52110 31054 52162 31106
rect 52162 31054 52164 31106
rect 52108 31052 52164 31054
rect 52556 31276 52612 31332
rect 52780 31164 52836 31220
rect 53452 31724 53508 31780
rect 51884 30210 51940 30212
rect 51884 30158 51886 30210
rect 51886 30158 51938 30210
rect 51938 30158 51940 30210
rect 51884 30156 51940 30158
rect 52780 30882 52836 30884
rect 52780 30830 52782 30882
rect 52782 30830 52834 30882
rect 52834 30830 52836 30882
rect 52780 30828 52836 30830
rect 54124 34076 54180 34132
rect 55468 36764 55524 36820
rect 56364 36764 56420 36820
rect 55020 36540 55076 36596
rect 55412 36540 55468 36596
rect 54684 35980 54740 36036
rect 55132 35868 55188 35924
rect 54796 35698 54852 35700
rect 54796 35646 54798 35698
rect 54798 35646 54850 35698
rect 54850 35646 54852 35698
rect 54796 35644 54852 35646
rect 55356 35698 55412 35700
rect 55356 35646 55358 35698
rect 55358 35646 55410 35698
rect 55410 35646 55412 35698
rect 55356 35644 55412 35646
rect 55132 35308 55188 35364
rect 55580 36316 55636 36372
rect 56028 36316 56084 36372
rect 55580 36092 55636 36148
rect 54460 34860 54516 34916
rect 54236 33740 54292 33796
rect 53900 33628 53956 33684
rect 54236 33292 54292 33348
rect 54012 32508 54068 32564
rect 53788 31276 53844 31332
rect 53788 31052 53844 31108
rect 53676 30322 53732 30324
rect 53676 30270 53678 30322
rect 53678 30270 53730 30322
rect 53730 30270 53732 30322
rect 53676 30268 53732 30270
rect 53116 30156 53172 30212
rect 53004 30098 53060 30100
rect 53004 30046 53006 30098
rect 53006 30046 53058 30098
rect 53058 30046 53060 30098
rect 53004 30044 53060 30046
rect 50988 27132 51044 27188
rect 51436 27580 51492 27636
rect 51212 27020 51268 27076
rect 52780 29986 52836 29988
rect 52780 29934 52782 29986
rect 52782 29934 52834 29986
rect 52834 29934 52836 29986
rect 52780 29932 52836 29934
rect 52892 29484 52948 29540
rect 53788 30044 53844 30100
rect 53564 29932 53620 29988
rect 53116 29372 53172 29428
rect 51772 28812 51828 28868
rect 51660 28476 51716 28532
rect 51660 28028 51716 28084
rect 51772 27970 51828 27972
rect 51772 27918 51774 27970
rect 51774 27918 51826 27970
rect 51826 27918 51828 27970
rect 51772 27916 51828 27918
rect 51660 27580 51716 27636
rect 51660 27356 51716 27412
rect 50988 26290 51044 26292
rect 50988 26238 50990 26290
rect 50990 26238 51042 26290
rect 51042 26238 51044 26290
rect 50988 26236 51044 26238
rect 50876 25788 50932 25844
rect 50876 25618 50932 25620
rect 50876 25566 50878 25618
rect 50878 25566 50930 25618
rect 50930 25566 50932 25618
rect 50876 25564 50932 25566
rect 50652 25506 50708 25508
rect 50652 25454 50654 25506
rect 50654 25454 50706 25506
rect 50706 25454 50708 25506
rect 50652 25452 50708 25454
rect 50204 25004 50260 25060
rect 49868 24220 49924 24276
rect 49868 23660 49924 23716
rect 49980 24780 50036 24836
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 51548 26460 51604 26516
rect 51324 26290 51380 26292
rect 51324 26238 51326 26290
rect 51326 26238 51378 26290
rect 51378 26238 51380 26290
rect 51324 26236 51380 26238
rect 51324 25564 51380 25620
rect 50988 24892 51044 24948
rect 51100 24834 51156 24836
rect 51100 24782 51102 24834
rect 51102 24782 51154 24834
rect 51154 24782 51156 24834
rect 51100 24780 51156 24782
rect 50316 24668 50372 24724
rect 50988 24668 51044 24724
rect 50092 24556 50148 24612
rect 50428 24498 50484 24500
rect 50428 24446 50430 24498
rect 50430 24446 50482 24498
rect 50482 24446 50484 24498
rect 50428 24444 50484 24446
rect 50204 24332 50260 24388
rect 50764 23996 50820 24052
rect 50876 23938 50932 23940
rect 50876 23886 50878 23938
rect 50878 23886 50930 23938
rect 50930 23886 50932 23938
rect 50876 23884 50932 23886
rect 49980 23492 50036 23548
rect 49756 22764 49812 22820
rect 49868 22988 49924 23044
rect 50092 22876 50148 22932
rect 49980 22258 50036 22260
rect 49980 22206 49982 22258
rect 49982 22206 50034 22258
rect 50034 22206 50036 22258
rect 49980 22204 50036 22206
rect 48972 21586 49028 21588
rect 48972 21534 48974 21586
rect 48974 21534 49026 21586
rect 49026 21534 49028 21586
rect 48972 21532 49028 21534
rect 49756 21980 49812 22036
rect 49644 21756 49700 21812
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50316 23324 50372 23380
rect 50764 23324 50820 23380
rect 50540 23154 50596 23156
rect 50540 23102 50542 23154
rect 50542 23102 50594 23154
rect 50594 23102 50596 23154
rect 50540 23100 50596 23102
rect 50764 22988 50820 23044
rect 50764 22540 50820 22596
rect 50428 22316 50484 22372
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 51436 25228 51492 25284
rect 51548 25452 51604 25508
rect 51436 23938 51492 23940
rect 51436 23886 51438 23938
rect 51438 23886 51490 23938
rect 51490 23886 51492 23938
rect 51436 23884 51492 23886
rect 51660 25340 51716 25396
rect 51660 23324 51716 23380
rect 52780 28476 52836 28532
rect 52332 27858 52388 27860
rect 52332 27806 52334 27858
rect 52334 27806 52386 27858
rect 52386 27806 52388 27858
rect 52332 27804 52388 27806
rect 51996 26850 52052 26852
rect 51996 26798 51998 26850
rect 51998 26798 52050 26850
rect 52050 26798 52052 26850
rect 51996 26796 52052 26798
rect 51884 26460 51940 26516
rect 52332 27020 52388 27076
rect 53564 28924 53620 28980
rect 52780 27186 52836 27188
rect 52780 27134 52782 27186
rect 52782 27134 52834 27186
rect 52834 27134 52836 27186
rect 52780 27132 52836 27134
rect 53228 27356 53284 27412
rect 53676 28812 53732 28868
rect 53340 27020 53396 27076
rect 52556 26236 52612 26292
rect 52556 25676 52612 25732
rect 52892 25618 52948 25620
rect 52892 25566 52894 25618
rect 52894 25566 52946 25618
rect 52946 25566 52948 25618
rect 52892 25564 52948 25566
rect 51996 25340 52052 25396
rect 52668 25228 52724 25284
rect 52556 24780 52612 24836
rect 51996 24722 52052 24724
rect 51996 24670 51998 24722
rect 51998 24670 52050 24722
rect 52050 24670 52052 24722
rect 51996 24668 52052 24670
rect 51436 23212 51492 23268
rect 51884 23212 51940 23268
rect 51100 22930 51156 22932
rect 51100 22878 51102 22930
rect 51102 22878 51154 22930
rect 51154 22878 51156 22930
rect 51100 22876 51156 22878
rect 51212 22482 51268 22484
rect 51212 22430 51214 22482
rect 51214 22430 51266 22482
rect 51266 22430 51268 22482
rect 51212 22428 51268 22430
rect 51772 22876 51828 22932
rect 52332 23378 52388 23380
rect 52332 23326 52334 23378
rect 52334 23326 52386 23378
rect 52386 23326 52388 23378
rect 52332 23324 52388 23326
rect 53900 29260 53956 29316
rect 53788 28700 53844 28756
rect 54012 28588 54068 28644
rect 53788 27916 53844 27972
rect 56140 36092 56196 36148
rect 55580 35084 55636 35140
rect 55804 35532 55860 35588
rect 55356 34860 55412 34916
rect 54684 34636 54740 34692
rect 55916 35420 55972 35476
rect 56700 35868 56756 35924
rect 57036 36092 57092 36148
rect 57260 36258 57316 36260
rect 57260 36206 57262 36258
rect 57262 36206 57314 36258
rect 57314 36206 57316 36258
rect 57260 36204 57316 36206
rect 57820 36258 57876 36260
rect 57820 36206 57822 36258
rect 57822 36206 57874 36258
rect 57874 36206 57876 36258
rect 57820 36204 57876 36206
rect 57372 35980 57428 36036
rect 56700 35586 56756 35588
rect 56700 35534 56702 35586
rect 56702 35534 56754 35586
rect 56754 35534 56756 35586
rect 56700 35532 56756 35534
rect 56812 34914 56868 34916
rect 56812 34862 56814 34914
rect 56814 34862 56866 34914
rect 56866 34862 56868 34914
rect 56812 34860 56868 34862
rect 56588 34802 56644 34804
rect 56588 34750 56590 34802
rect 56590 34750 56642 34802
rect 56642 34750 56644 34802
rect 56588 34748 56644 34750
rect 57148 35308 57204 35364
rect 57036 35084 57092 35140
rect 56812 34636 56868 34692
rect 56028 34242 56084 34244
rect 56028 34190 56030 34242
rect 56030 34190 56082 34242
rect 56082 34190 56084 34242
rect 56028 34188 56084 34190
rect 56476 33964 56532 34020
rect 54796 32674 54852 32676
rect 54796 32622 54798 32674
rect 54798 32622 54850 32674
rect 54850 32622 54852 32674
rect 54796 32620 54852 32622
rect 54348 31276 54404 31332
rect 54572 31052 54628 31108
rect 56812 34130 56868 34132
rect 56812 34078 56814 34130
rect 56814 34078 56866 34130
rect 56866 34078 56868 34130
rect 56812 34076 56868 34078
rect 55244 32620 55300 32676
rect 57148 34188 57204 34244
rect 57260 34860 57316 34916
rect 57708 35474 57764 35476
rect 57708 35422 57710 35474
rect 57710 35422 57762 35474
rect 57762 35422 57764 35474
rect 57708 35420 57764 35422
rect 57820 35308 57876 35364
rect 57708 34690 57764 34692
rect 57708 34638 57710 34690
rect 57710 34638 57762 34690
rect 57762 34638 57764 34690
rect 57708 34636 57764 34638
rect 57932 33292 57988 33348
rect 56700 31500 56756 31556
rect 54908 30994 54964 30996
rect 54908 30942 54910 30994
rect 54910 30942 54962 30994
rect 54962 30942 54964 30994
rect 54908 30940 54964 30942
rect 55356 30994 55412 30996
rect 55356 30942 55358 30994
rect 55358 30942 55410 30994
rect 55410 30942 55412 30994
rect 55356 30940 55412 30942
rect 54572 30322 54628 30324
rect 54572 30270 54574 30322
rect 54574 30270 54626 30322
rect 54626 30270 54628 30322
rect 54572 30268 54628 30270
rect 57372 30940 57428 30996
rect 58044 30940 58100 30996
rect 54796 29426 54852 29428
rect 54796 29374 54798 29426
rect 54798 29374 54850 29426
rect 54850 29374 54852 29426
rect 54796 29372 54852 29374
rect 54460 29260 54516 29316
rect 54236 28924 54292 28980
rect 54124 28028 54180 28084
rect 54908 28754 54964 28756
rect 54908 28702 54910 28754
rect 54910 28702 54962 28754
rect 54962 28702 54964 28754
rect 54908 28700 54964 28702
rect 55356 28812 55412 28868
rect 56252 28812 56308 28868
rect 55468 28364 55524 28420
rect 54460 27916 54516 27972
rect 55020 28140 55076 28196
rect 55020 27858 55076 27860
rect 55020 27806 55022 27858
rect 55022 27806 55074 27858
rect 55074 27806 55076 27858
rect 55020 27804 55076 27806
rect 54236 27746 54292 27748
rect 54236 27694 54238 27746
rect 54238 27694 54290 27746
rect 54290 27694 54292 27746
rect 54236 27692 54292 27694
rect 54348 27580 54404 27636
rect 53676 26796 53732 26852
rect 53340 24780 53396 24836
rect 53900 26402 53956 26404
rect 53900 26350 53902 26402
rect 53902 26350 53954 26402
rect 53954 26350 53956 26402
rect 53900 26348 53956 26350
rect 56476 28642 56532 28644
rect 56476 28590 56478 28642
rect 56478 28590 56530 28642
rect 56530 28590 56532 28642
rect 56476 28588 56532 28590
rect 55692 28140 55748 28196
rect 56812 28028 56868 28084
rect 56588 27970 56644 27972
rect 56588 27918 56590 27970
rect 56590 27918 56642 27970
rect 56642 27918 56644 27970
rect 56588 27916 56644 27918
rect 55580 27692 55636 27748
rect 57708 27692 57764 27748
rect 54460 26962 54516 26964
rect 54460 26910 54462 26962
rect 54462 26910 54514 26962
rect 54514 26910 54516 26962
rect 54460 26908 54516 26910
rect 54908 26908 54964 26964
rect 53900 25730 53956 25732
rect 53900 25678 53902 25730
rect 53902 25678 53954 25730
rect 53954 25678 53956 25730
rect 53900 25676 53956 25678
rect 54460 25394 54516 25396
rect 54460 25342 54462 25394
rect 54462 25342 54514 25394
rect 54514 25342 54516 25394
rect 54460 25340 54516 25342
rect 53676 24668 53732 24724
rect 53228 24220 53284 24276
rect 52780 23826 52836 23828
rect 52780 23774 52782 23826
rect 52782 23774 52834 23826
rect 52834 23774 52836 23826
rect 52780 23772 52836 23774
rect 52108 23100 52164 23156
rect 53004 23266 53060 23268
rect 53004 23214 53006 23266
rect 53006 23214 53058 23266
rect 53058 23214 53060 23266
rect 53004 23212 53060 23214
rect 51996 22316 52052 22372
rect 49644 21586 49700 21588
rect 49644 21534 49646 21586
rect 49646 21534 49698 21586
rect 49698 21534 49700 21586
rect 49644 21532 49700 21534
rect 49084 21420 49140 21476
rect 49532 21362 49588 21364
rect 49532 21310 49534 21362
rect 49534 21310 49586 21362
rect 49586 21310 49588 21362
rect 49532 21308 49588 21310
rect 48300 21196 48356 21252
rect 48636 20914 48692 20916
rect 48636 20862 48638 20914
rect 48638 20862 48690 20914
rect 48690 20862 48692 20914
rect 48636 20860 48692 20862
rect 53340 22988 53396 23044
rect 49868 20914 49924 20916
rect 49868 20862 49870 20914
rect 49870 20862 49922 20914
rect 49922 20862 49924 20914
rect 49868 20860 49924 20862
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 38556 19852 38612 19908
rect 35308 18956 35364 19012
rect 33628 15484 33684 15540
rect 33852 15596 33908 15652
rect 34748 16044 34804 16100
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35084 16604 35140 16660
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35532 16044 35588 16100
rect 34524 15260 34580 15316
rect 34188 15202 34244 15204
rect 34188 15150 34190 15202
rect 34190 15150 34242 15202
rect 34242 15150 34244 15202
rect 34188 15148 34244 15150
rect 30716 12348 30772 12404
rect 30380 11618 30436 11620
rect 30380 11566 30382 11618
rect 30382 11566 30434 11618
rect 30434 11566 30436 11618
rect 30380 11564 30436 11566
rect 30716 11564 30772 11620
rect 31500 11676 31556 11732
rect 30604 11452 30660 11508
rect 29596 10834 29652 10836
rect 29596 10782 29598 10834
rect 29598 10782 29650 10834
rect 29650 10782 29652 10834
rect 29596 10780 29652 10782
rect 30268 10834 30324 10836
rect 30268 10782 30270 10834
rect 30270 10782 30322 10834
rect 30322 10782 30324 10834
rect 30268 10780 30324 10782
rect 30940 11282 30996 11284
rect 30940 11230 30942 11282
rect 30942 11230 30994 11282
rect 30994 11230 30996 11282
rect 30940 11228 30996 11230
rect 31500 10780 31556 10836
rect 30828 10722 30884 10724
rect 30828 10670 30830 10722
rect 30830 10670 30882 10722
rect 30882 10670 30884 10722
rect 30828 10668 30884 10670
rect 30156 9602 30212 9604
rect 30156 9550 30158 9602
rect 30158 9550 30210 9602
rect 30210 9550 30212 9602
rect 30156 9548 30212 9550
rect 31388 9548 31444 9604
rect 33964 11900 34020 11956
rect 34300 12012 34356 12068
rect 33628 11676 33684 11732
rect 33852 11340 33908 11396
rect 35084 15148 35140 15204
rect 35420 15202 35476 15204
rect 35420 15150 35422 15202
rect 35422 15150 35474 15202
rect 35474 15150 35476 15202
rect 35420 15148 35476 15150
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34972 14028 35028 14084
rect 35084 13580 35140 13636
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 36988 18956 37044 19012
rect 37548 19010 37604 19012
rect 37548 18958 37550 19010
rect 37550 18958 37602 19010
rect 37602 18958 37604 19010
rect 37548 18956 37604 18958
rect 38220 18956 38276 19012
rect 39788 19906 39844 19908
rect 39788 19854 39790 19906
rect 39790 19854 39842 19906
rect 39842 19854 39844 19906
rect 39788 19852 39844 19854
rect 42140 19906 42196 19908
rect 42140 19854 42142 19906
rect 42142 19854 42194 19906
rect 42194 19854 42196 19906
rect 42140 19852 42196 19854
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 36988 18284 37044 18340
rect 36092 17554 36148 17556
rect 36092 17502 36094 17554
rect 36094 17502 36146 17554
rect 36146 17502 36148 17554
rect 36092 17500 36148 17502
rect 37436 17500 37492 17556
rect 36428 16604 36484 16660
rect 36092 15874 36148 15876
rect 36092 15822 36094 15874
rect 36094 15822 36146 15874
rect 36146 15822 36148 15874
rect 36092 15820 36148 15822
rect 37548 15820 37604 15876
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 35756 14028 35812 14084
rect 34524 11676 34580 11732
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35980 12066 36036 12068
rect 35980 12014 35982 12066
rect 35982 12014 36034 12066
rect 36034 12014 36036 12066
rect 35980 12012 36036 12014
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 35532 11618 35588 11620
rect 35532 11566 35534 11618
rect 35534 11566 35586 11618
rect 35586 11566 35588 11618
rect 35532 11564 35588 11566
rect 35980 11788 36036 11844
rect 35756 11340 35812 11396
rect 37100 12124 37156 12180
rect 39116 12178 39172 12180
rect 39116 12126 39118 12178
rect 39118 12126 39170 12178
rect 39170 12126 39172 12178
rect 39116 12124 39172 12126
rect 38444 11788 38500 11844
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 31276 8316 31332 8372
rect 32844 8370 32900 8372
rect 32844 8318 32846 8370
rect 32846 8318 32898 8370
rect 32898 8318 32900 8370
rect 32844 8316 32900 8318
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 27020 5740 27076 5796
rect 26684 4508 26740 4564
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 28252 5740 28308 5796
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 27916 4172 27972 4228
rect 29596 4226 29652 4228
rect 29596 4174 29598 4226
rect 29598 4174 29650 4226
rect 29650 4174 29652 4226
rect 29596 4172 29652 4174
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 15586 57036 15596 57092
rect 15652 57036 17500 57092
rect 17556 57036 17566 57092
rect 32274 57036 32284 57092
rect 32340 57036 34188 57092
rect 34244 57036 34254 57092
rect 34962 57036 34972 57092
rect 35028 57036 37996 57092
rect 38052 57036 38062 57092
rect 41010 57036 41020 57092
rect 41076 57036 42924 57092
rect 42980 57036 42990 57092
rect 33618 56924 33628 56980
rect 33684 56924 36428 56980
rect 36484 56924 36494 56980
rect 42130 56924 42140 56980
rect 42196 56924 44044 56980
rect 44100 56924 44110 56980
rect 38994 56812 39004 56868
rect 39060 56812 42028 56868
rect 42084 56812 42094 56868
rect 37650 56700 37660 56756
rect 37716 56700 40460 56756
rect 40516 56700 40526 56756
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4610 56252 4620 56308
rect 4676 56252 5516 56308
rect 5572 56252 5582 56308
rect 15698 56252 15708 56308
rect 15764 56252 15774 56308
rect 29586 56252 29596 56308
rect 29652 56252 30716 56308
rect 30772 56252 30782 56308
rect 30930 56252 30940 56308
rect 30996 56252 32620 56308
rect 32676 56252 32686 56308
rect 34066 56252 34076 56308
rect 34132 56252 35308 56308
rect 35364 56252 35374 56308
rect 36754 56252 36764 56308
rect 36820 56252 39116 56308
rect 39172 56252 39182 56308
rect 41682 56252 41692 56308
rect 41748 56252 43596 56308
rect 43652 56252 43662 56308
rect 5842 56140 5852 56196
rect 5908 56140 8428 56196
rect 8484 56140 8494 56196
rect 15708 56084 15764 56252
rect 14802 56028 14812 56084
rect 14868 56028 15764 56084
rect 33842 56028 33852 56084
rect 33908 56028 35980 56084
rect 36036 56028 36046 56084
rect 15138 55916 15148 55972
rect 15204 55916 17052 55972
rect 17108 55916 17118 55972
rect 27794 55916 27804 55972
rect 27860 55916 29932 55972
rect 29988 55916 29998 55972
rect 43474 55916 43484 55972
rect 43540 55916 44492 55972
rect 44548 55916 44558 55972
rect 44818 55804 44828 55860
rect 44884 55804 45388 55860
rect 45444 55804 45454 55860
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 17938 55468 17948 55524
rect 18004 55468 19180 55524
rect 19236 55468 19246 55524
rect 35298 55468 35308 55524
rect 35364 55468 37548 55524
rect 37604 55468 37614 55524
rect 16482 55356 16492 55412
rect 16548 55356 18508 55412
rect 18564 55356 19852 55412
rect 19908 55356 19918 55412
rect 36306 55356 36316 55412
rect 36372 55356 37436 55412
rect 37492 55356 37502 55412
rect 16594 55244 16604 55300
rect 16660 55244 17612 55300
rect 17668 55244 18284 55300
rect 18340 55244 18350 55300
rect 18946 55244 18956 55300
rect 19012 55244 20188 55300
rect 20244 55244 20254 55300
rect 16818 55132 16828 55188
rect 16884 55132 19628 55188
rect 19684 55132 19694 55188
rect 41794 55132 41804 55188
rect 41860 55132 42924 55188
rect 42980 55132 42990 55188
rect 17826 55020 17836 55076
rect 17892 55020 18844 55076
rect 18900 55020 18910 55076
rect 25106 54908 25116 54964
rect 25172 54908 26124 54964
rect 26180 54908 26190 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 17938 54684 17948 54740
rect 18004 54684 19180 54740
rect 19236 54684 19246 54740
rect 28242 54684 28252 54740
rect 28308 54684 29260 54740
rect 29316 54684 29326 54740
rect 9202 54460 9212 54516
rect 9268 54460 9996 54516
rect 10052 54460 12124 54516
rect 12180 54460 12190 54516
rect 17378 54460 17388 54516
rect 17444 54460 19516 54516
rect 19572 54460 19582 54516
rect 23090 54460 23100 54516
rect 23156 54460 24332 54516
rect 24388 54460 24398 54516
rect 23874 54348 23884 54404
rect 23940 54348 24668 54404
rect 24724 54348 25228 54404
rect 25284 54348 25788 54404
rect 25844 54348 29148 54404
rect 29204 54348 29708 54404
rect 29764 54348 30940 54404
rect 30996 54348 32060 54404
rect 32116 54348 32508 54404
rect 32564 54348 34188 54404
rect 34244 54348 34254 54404
rect 16258 54236 16268 54292
rect 16324 54236 17500 54292
rect 17556 54236 18284 54292
rect 18340 54236 18350 54292
rect 39106 54236 39116 54292
rect 39172 54236 39452 54292
rect 39508 54236 39518 54292
rect 43026 54236 43036 54292
rect 43092 54236 43708 54292
rect 43764 54236 44828 54292
rect 44884 54236 44894 54292
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 26450 54012 26460 54068
rect 26516 54012 33516 54068
rect 33572 54012 33582 54068
rect 12898 53900 12908 53956
rect 12964 53900 13468 53956
rect 13524 53900 13534 53956
rect 16482 53900 16492 53956
rect 16548 53900 17164 53956
rect 17220 53900 18620 53956
rect 18676 53900 18686 53956
rect 28242 53900 28252 53956
rect 28308 53900 39620 53956
rect 39564 53844 39620 53900
rect 4050 53788 4060 53844
rect 4116 53788 9324 53844
rect 9380 53788 9390 53844
rect 10658 53788 10668 53844
rect 10724 53788 13580 53844
rect 13636 53788 13646 53844
rect 35196 53788 38556 53844
rect 38612 53788 38622 53844
rect 39554 53788 39564 53844
rect 39620 53788 39630 53844
rect 21522 53676 21532 53732
rect 21588 53676 22204 53732
rect 22260 53676 22270 53732
rect 35196 53620 35252 53788
rect 37874 53676 37884 53732
rect 37940 53676 38332 53732
rect 38388 53676 38668 53732
rect 38724 53676 38734 53732
rect 38882 53676 38892 53732
rect 38948 53676 39116 53732
rect 39172 53676 39182 53732
rect 39330 53676 39340 53732
rect 39396 53676 41804 53732
rect 41860 53676 42252 53732
rect 42308 53676 42318 53732
rect 42578 53676 42588 53732
rect 42644 53676 45052 53732
rect 45108 53676 45500 53732
rect 45556 53676 46956 53732
rect 47012 53676 48748 53732
rect 48804 53676 48814 53732
rect 20962 53564 20972 53620
rect 21028 53564 23548 53620
rect 23604 53564 23614 53620
rect 30370 53564 30380 53620
rect 30436 53564 34748 53620
rect 34804 53564 34814 53620
rect 35186 53564 35196 53620
rect 35252 53564 35262 53620
rect 37986 53564 37996 53620
rect 38052 53564 39452 53620
rect 39508 53564 39518 53620
rect 46274 53564 46284 53620
rect 46340 53564 48860 53620
rect 48916 53564 48926 53620
rect 16818 53452 16828 53508
rect 16884 53452 17836 53508
rect 17892 53452 17902 53508
rect 38098 53452 38108 53508
rect 38164 53452 39340 53508
rect 39396 53452 39406 53508
rect 39554 53452 39564 53508
rect 39620 53452 39900 53508
rect 39956 53452 39966 53508
rect 34066 53340 34076 53396
rect 34132 53340 38444 53396
rect 38500 53340 38510 53396
rect 39218 53340 39228 53396
rect 39284 53340 39788 53396
rect 39844 53340 39854 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 34514 53228 34524 53284
rect 34580 53228 35868 53284
rect 35924 53228 35934 53284
rect 38658 53228 38668 53284
rect 38724 53228 40908 53284
rect 40964 53228 40974 53284
rect 23762 53116 23772 53172
rect 23828 53116 24220 53172
rect 24276 53116 24286 53172
rect 33170 53116 33180 53172
rect 33236 53116 33964 53172
rect 34020 53116 34030 53172
rect 39218 53116 39228 53172
rect 39284 53116 40236 53172
rect 40292 53116 42140 53172
rect 42196 53116 42588 53172
rect 42644 53116 42654 53172
rect 8082 53004 8092 53060
rect 8148 53004 8540 53060
rect 8596 53004 9548 53060
rect 9604 53004 9614 53060
rect 22418 53004 22428 53060
rect 22484 53004 24052 53060
rect 24546 53004 24556 53060
rect 24612 53004 25004 53060
rect 25060 53004 25340 53060
rect 25396 53004 25406 53060
rect 35298 53004 35308 53060
rect 35364 53004 38108 53060
rect 38164 53004 38174 53060
rect 23996 52948 24052 53004
rect 3826 52892 3836 52948
rect 3892 52892 4508 52948
rect 4564 52892 4574 52948
rect 4946 52892 4956 52948
rect 5012 52892 5022 52948
rect 11442 52892 11452 52948
rect 11508 52892 12796 52948
rect 12852 52892 12862 52948
rect 18732 52892 19180 52948
rect 19236 52892 19246 52948
rect 19842 52892 19852 52948
rect 19908 52892 20636 52948
rect 20692 52892 20702 52948
rect 22194 52892 22204 52948
rect 22260 52892 23548 52948
rect 23604 52892 23614 52948
rect 23986 52892 23996 52948
rect 24052 52892 24062 52948
rect 32274 52892 32284 52948
rect 32340 52892 37212 52948
rect 37268 52892 37278 52948
rect 37874 52892 37884 52948
rect 37940 52892 39788 52948
rect 39844 52892 39854 52948
rect 41122 52892 41132 52948
rect 41188 52892 41916 52948
rect 41972 52892 41982 52948
rect 43922 52892 43932 52948
rect 43988 52892 45948 52948
rect 46004 52892 46014 52948
rect 49970 52892 49980 52948
rect 50036 52892 51436 52948
rect 51492 52892 51502 52948
rect 4956 52836 5012 52892
rect 18732 52836 18788 52892
rect 3266 52780 3276 52836
rect 3332 52780 6188 52836
rect 6244 52780 6254 52836
rect 10882 52780 10892 52836
rect 10948 52780 12012 52836
rect 12068 52780 13468 52836
rect 13524 52780 13916 52836
rect 13972 52780 13982 52836
rect 17714 52780 17724 52836
rect 17780 52780 18732 52836
rect 18788 52780 18798 52836
rect 19282 52780 19292 52836
rect 19348 52780 20860 52836
rect 20916 52780 20926 52836
rect 35410 52780 35420 52836
rect 35476 52780 35644 52836
rect 35700 52780 35710 52836
rect 38210 52780 38220 52836
rect 38276 52780 38892 52836
rect 38948 52780 39676 52836
rect 39732 52780 39742 52836
rect 25554 52668 25564 52724
rect 25620 52668 27132 52724
rect 27188 52668 27198 52724
rect 35298 52668 35308 52724
rect 35364 52668 35700 52724
rect 36306 52668 36316 52724
rect 36372 52668 38444 52724
rect 38500 52668 38668 52724
rect 39218 52668 39228 52724
rect 39284 52668 41020 52724
rect 41076 52668 41086 52724
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 35644 52500 35700 52668
rect 13682 52444 13692 52500
rect 13748 52444 15932 52500
rect 15988 52444 15998 52500
rect 20738 52444 20748 52500
rect 20804 52444 25564 52500
rect 25620 52444 25630 52500
rect 35634 52444 35644 52500
rect 35700 52444 35710 52500
rect 4386 52332 4396 52388
rect 4452 52332 5012 52388
rect 6402 52332 6412 52388
rect 6468 52332 7532 52388
rect 7588 52332 7598 52388
rect 12562 52332 12572 52388
rect 12628 52332 14812 52388
rect 14868 52332 14878 52388
rect 36194 52332 36204 52388
rect 36260 52332 37996 52388
rect 38052 52332 38062 52388
rect 4956 52276 5012 52332
rect 38612 52276 38668 52668
rect 38882 52332 38892 52388
rect 38948 52332 40796 52388
rect 40852 52332 40862 52388
rect 48850 52332 48860 52388
rect 48916 52332 50652 52388
rect 50708 52332 50718 52388
rect 4946 52220 4956 52276
rect 5012 52220 6300 52276
rect 6356 52220 6748 52276
rect 6804 52220 6814 52276
rect 11554 52220 11564 52276
rect 11620 52220 12460 52276
rect 12516 52220 15708 52276
rect 15764 52220 15774 52276
rect 18946 52220 18956 52276
rect 19012 52220 20188 52276
rect 20244 52220 20748 52276
rect 20804 52220 20814 52276
rect 24546 52220 24556 52276
rect 24612 52220 25228 52276
rect 25284 52220 25294 52276
rect 35522 52220 35532 52276
rect 35588 52220 36316 52276
rect 36372 52220 36382 52276
rect 37650 52220 37660 52276
rect 37716 52220 38444 52276
rect 38500 52220 38510 52276
rect 38612 52220 41804 52276
rect 41860 52220 41870 52276
rect 49410 52220 49420 52276
rect 49476 52220 49980 52276
rect 50036 52220 50046 52276
rect 50204 52220 51884 52276
rect 51940 52220 51950 52276
rect 50204 52164 50260 52220
rect 6626 52108 6636 52164
rect 6692 52108 7196 52164
rect 7252 52108 7262 52164
rect 13122 52108 13132 52164
rect 13188 52108 13804 52164
rect 13860 52108 13870 52164
rect 15474 52108 15484 52164
rect 15540 52108 17948 52164
rect 18004 52108 18732 52164
rect 18788 52108 19740 52164
rect 19796 52108 20076 52164
rect 20132 52108 20972 52164
rect 21028 52108 21038 52164
rect 22978 52108 22988 52164
rect 23044 52108 23548 52164
rect 23604 52108 23614 52164
rect 39442 52108 39452 52164
rect 39508 52108 40012 52164
rect 40068 52108 42028 52164
rect 42084 52108 42094 52164
rect 49746 52108 49756 52164
rect 49812 52108 50260 52164
rect 50316 52108 50764 52164
rect 50820 52108 50830 52164
rect 50316 52052 50372 52108
rect 3602 51996 3612 52052
rect 3668 51996 4396 52052
rect 4452 51996 4462 52052
rect 9202 51996 9212 52052
rect 9268 51996 11676 52052
rect 11732 51996 11742 52052
rect 20626 51996 20636 52052
rect 20692 51996 22764 52052
rect 22820 51996 23100 52052
rect 23156 51996 23166 52052
rect 31154 51996 31164 52052
rect 31220 51996 34860 52052
rect 34916 51996 34926 52052
rect 35746 51996 35756 52052
rect 35812 51996 36316 52052
rect 36372 51996 38220 52052
rect 38276 51996 38286 52052
rect 38770 51996 38780 52052
rect 38836 51996 40404 52052
rect 41570 51996 41580 52052
rect 41636 51996 42700 52052
rect 42756 51996 42766 52052
rect 49186 51996 49196 52052
rect 49252 51996 49420 52052
rect 49476 51996 49980 52052
rect 50036 51996 50204 52052
rect 50260 51996 50372 52052
rect 40348 51940 40404 51996
rect 2482 51884 2492 51940
rect 2548 51884 4284 51940
rect 4340 51884 4350 51940
rect 35298 51884 35308 51940
rect 35364 51884 35644 51940
rect 35700 51884 35710 51940
rect 37986 51884 37996 51940
rect 38052 51884 39452 51940
rect 39508 51884 39518 51940
rect 40348 51884 43820 51940
rect 43876 51884 43886 51940
rect 46722 51884 46732 51940
rect 46788 51884 47068 51940
rect 47124 51884 47134 51940
rect 50978 51884 50988 51940
rect 51044 51884 52444 51940
rect 52500 51884 52510 51940
rect 38770 51772 38780 51828
rect 38836 51772 38874 51828
rect 40114 51772 40124 51828
rect 40180 51772 42140 51828
rect 42196 51772 42812 51828
rect 42868 51772 43484 51828
rect 43540 51772 43550 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 18274 51660 18284 51716
rect 18340 51660 19068 51716
rect 19124 51660 19134 51716
rect 22866 51660 22876 51716
rect 22932 51660 25228 51716
rect 25284 51660 25294 51716
rect 38098 51660 38108 51716
rect 38164 51660 41916 51716
rect 41972 51660 41982 51716
rect 22306 51548 22316 51604
rect 22372 51548 23660 51604
rect 23716 51548 23726 51604
rect 28578 51548 28588 51604
rect 28644 51548 30492 51604
rect 30548 51548 31836 51604
rect 31892 51548 31902 51604
rect 35522 51548 35532 51604
rect 35588 51548 35980 51604
rect 36036 51548 36046 51604
rect 37874 51548 37884 51604
rect 37940 51548 38556 51604
rect 38612 51548 38622 51604
rect 10322 51436 10332 51492
rect 10388 51436 11340 51492
rect 11396 51436 14476 51492
rect 14532 51436 14542 51492
rect 15362 51436 15372 51492
rect 15428 51436 17388 51492
rect 17444 51436 18284 51492
rect 18340 51436 18620 51492
rect 18676 51436 18686 51492
rect 23090 51436 23100 51492
rect 23156 51436 24332 51492
rect 24388 51436 24398 51492
rect 34178 51436 34188 51492
rect 34244 51436 35420 51492
rect 35476 51436 37100 51492
rect 37156 51436 37166 51492
rect 38210 51436 38220 51492
rect 38276 51436 38444 51492
rect 38500 51436 38510 51492
rect 46386 51436 46396 51492
rect 46452 51436 48076 51492
rect 48132 51436 48142 51492
rect 49858 51436 49868 51492
rect 49924 51436 50876 51492
rect 50932 51436 50942 51492
rect 14018 51324 14028 51380
rect 14084 51324 14364 51380
rect 14420 51324 15148 51380
rect 15586 51324 15596 51380
rect 15652 51324 16156 51380
rect 16212 51324 16222 51380
rect 34402 51324 34412 51380
rect 34468 51324 35644 51380
rect 35700 51324 35710 51380
rect 35970 51324 35980 51380
rect 36036 51324 37772 51380
rect 37828 51324 37838 51380
rect 42140 51324 43708 51380
rect 43764 51324 45052 51380
rect 45108 51324 45118 51380
rect 46946 51324 46956 51380
rect 47012 51324 51660 51380
rect 51716 51324 52668 51380
rect 52724 51324 52734 51380
rect 15092 51268 15148 51324
rect 42140 51268 42196 51324
rect 15092 51212 15260 51268
rect 15316 51212 16044 51268
rect 16100 51212 17612 51268
rect 17668 51212 17678 51268
rect 20066 51212 20076 51268
rect 20132 51212 22092 51268
rect 22148 51212 22158 51268
rect 24434 51212 24444 51268
rect 24500 51212 27356 51268
rect 27412 51212 27422 51268
rect 33954 51212 33964 51268
rect 34020 51212 34972 51268
rect 35028 51212 39004 51268
rect 39060 51212 39676 51268
rect 39732 51212 39742 51268
rect 42130 51212 42140 51268
rect 42196 51212 42206 51268
rect 45602 51212 45612 51268
rect 45668 51212 48860 51268
rect 48916 51212 51772 51268
rect 51828 51212 54572 51268
rect 54628 51212 54638 51268
rect 8754 51100 8764 51156
rect 8820 51100 10108 51156
rect 10164 51100 10174 51156
rect 11330 51100 11340 51156
rect 11396 51100 12012 51156
rect 12068 51100 12078 51156
rect 16818 51100 16828 51156
rect 16884 51100 18396 51156
rect 18452 51100 18956 51156
rect 19012 51100 19022 51156
rect 34738 51100 34748 51156
rect 34804 51100 35868 51156
rect 35924 51100 35934 51156
rect 38770 51100 38780 51156
rect 38836 51100 38892 51156
rect 38948 51100 38958 51156
rect 41234 51100 41244 51156
rect 41300 51100 42252 51156
rect 42308 51100 43372 51156
rect 43428 51100 43438 51156
rect 45826 51100 45836 51156
rect 45892 51100 46732 51156
rect 46788 51100 47516 51156
rect 47572 51100 47964 51156
rect 48020 51100 48030 51156
rect 49858 51100 49868 51156
rect 49924 51100 50316 51156
rect 50372 51100 50382 51156
rect 10210 50988 10220 51044
rect 10276 50988 13692 51044
rect 13748 50988 13758 51044
rect 19618 50988 19628 51044
rect 19684 50988 20188 51044
rect 20244 50988 20254 51044
rect 35634 50988 35644 51044
rect 35700 50988 36988 51044
rect 37044 50988 39284 51044
rect 47058 50988 47068 51044
rect 47124 50988 48188 51044
rect 48244 50988 48254 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 18946 50876 18956 50932
rect 19012 50876 19852 50932
rect 19908 50876 19918 50932
rect 39228 50820 39284 50988
rect 41682 50876 41692 50932
rect 41748 50876 42364 50932
rect 42420 50876 42430 50932
rect 47730 50876 47740 50932
rect 47796 50876 49420 50932
rect 49476 50876 49486 50932
rect 3826 50764 3836 50820
rect 3892 50764 4620 50820
rect 4676 50764 6748 50820
rect 6804 50764 6814 50820
rect 15138 50764 15148 50820
rect 15204 50764 16604 50820
rect 16660 50764 19404 50820
rect 19460 50764 19470 50820
rect 19964 50764 23436 50820
rect 23492 50764 23502 50820
rect 37202 50764 37212 50820
rect 37268 50764 38332 50820
rect 38388 50764 38398 50820
rect 38994 50764 39004 50820
rect 39060 50764 39070 50820
rect 39228 50764 42420 50820
rect 43586 50764 43596 50820
rect 43652 50764 46620 50820
rect 46676 50764 46686 50820
rect 4946 50652 4956 50708
rect 5012 50652 6636 50708
rect 6692 50652 6702 50708
rect 12898 50652 12908 50708
rect 12964 50652 13468 50708
rect 13524 50652 13534 50708
rect 4050 50540 4060 50596
rect 4116 50540 5964 50596
rect 6020 50540 6860 50596
rect 6916 50540 6926 50596
rect 12562 50540 12572 50596
rect 12628 50540 14364 50596
rect 14420 50540 15036 50596
rect 15092 50540 15102 50596
rect 19964 50484 20020 50764
rect 39004 50708 39060 50764
rect 34402 50652 34412 50708
rect 34468 50652 37044 50708
rect 38210 50652 38220 50708
rect 38276 50652 39060 50708
rect 39190 50652 39228 50708
rect 39284 50652 39294 50708
rect 39442 50652 39452 50708
rect 39508 50652 41580 50708
rect 41636 50652 41972 50708
rect 36988 50596 37044 50652
rect 41916 50596 41972 50652
rect 21970 50540 21980 50596
rect 22036 50540 23884 50596
rect 23940 50540 23950 50596
rect 34290 50540 34300 50596
rect 34356 50540 35420 50596
rect 35476 50540 35486 50596
rect 36978 50540 36988 50596
rect 37044 50540 39116 50596
rect 39172 50540 40908 50596
rect 40964 50540 40974 50596
rect 41906 50540 41916 50596
rect 41972 50540 41982 50596
rect 42102 50540 42140 50596
rect 42196 50540 42206 50596
rect 9986 50428 9996 50484
rect 10052 50428 10892 50484
rect 10948 50428 11788 50484
rect 11844 50428 12348 50484
rect 12404 50428 14924 50484
rect 14980 50428 14990 50484
rect 18274 50428 18284 50484
rect 18340 50428 19180 50484
rect 19236 50428 19246 50484
rect 19394 50428 19404 50484
rect 19460 50428 19740 50484
rect 19796 50428 19806 50484
rect 19954 50428 19964 50484
rect 20020 50428 20030 50484
rect 22642 50428 22652 50484
rect 22708 50428 22876 50484
rect 22932 50428 22942 50484
rect 24098 50428 24108 50484
rect 24164 50428 25452 50484
rect 25508 50428 26908 50484
rect 26964 50428 26974 50484
rect 35074 50428 35084 50484
rect 35140 50428 38220 50484
rect 38276 50428 38286 50484
rect 38434 50428 38444 50484
rect 38500 50428 38668 50484
rect 38724 50428 38734 50484
rect 39218 50428 39228 50484
rect 39284 50428 40236 50484
rect 40292 50428 40302 50484
rect 42364 50372 42420 50764
rect 49420 50708 49476 50876
rect 42914 50652 42924 50708
rect 42980 50652 47068 50708
rect 47124 50652 47134 50708
rect 49420 50652 50764 50708
rect 50820 50652 55580 50708
rect 55636 50652 55646 50708
rect 42924 50596 42980 50652
rect 42690 50540 42700 50596
rect 42756 50540 42980 50596
rect 47506 50540 47516 50596
rect 47572 50540 48076 50596
rect 48132 50540 48142 50596
rect 48290 50540 48300 50596
rect 48356 50540 49308 50596
rect 49364 50540 49374 50596
rect 42914 50428 42924 50484
rect 42980 50428 43652 50484
rect 46162 50428 46172 50484
rect 46228 50428 47292 50484
rect 47348 50428 47740 50484
rect 47796 50428 47806 50484
rect 47954 50428 47964 50484
rect 48020 50428 49980 50484
rect 50036 50428 50046 50484
rect 51314 50428 51324 50484
rect 51380 50428 53452 50484
rect 53508 50428 53518 50484
rect 43596 50372 43652 50428
rect 5954 50316 5964 50372
rect 6020 50316 7420 50372
rect 7476 50316 7486 50372
rect 12562 50316 12572 50372
rect 12628 50316 13916 50372
rect 13972 50316 14812 50372
rect 14868 50316 14878 50372
rect 18610 50316 18620 50372
rect 18676 50316 19068 50372
rect 19124 50316 19134 50372
rect 36418 50316 36428 50372
rect 36484 50316 36652 50372
rect 36708 50316 36718 50372
rect 37324 50316 40012 50372
rect 40068 50316 40078 50372
rect 42354 50316 42364 50372
rect 42420 50316 42430 50372
rect 43586 50316 43596 50372
rect 43652 50316 43662 50372
rect 37324 50260 37380 50316
rect 36866 50204 36876 50260
rect 36932 50204 37324 50260
rect 37380 50204 37390 50260
rect 37548 50204 39508 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 37548 50148 37604 50204
rect 39452 50148 39508 50204
rect 42812 50204 48524 50260
rect 48580 50204 48590 50260
rect 42812 50148 42868 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 5730 50092 5740 50148
rect 5796 50092 6188 50148
rect 6244 50092 6254 50148
rect 36754 50092 36764 50148
rect 36820 50092 37604 50148
rect 37986 50092 37996 50148
rect 38052 50092 39116 50148
rect 39172 50092 39182 50148
rect 39452 50092 42868 50148
rect 43026 50092 43036 50148
rect 43092 50092 43102 50148
rect 18722 49980 18732 50036
rect 18788 49980 18798 50036
rect 38658 49980 38668 50036
rect 38724 49980 40012 50036
rect 40068 49980 41356 50036
rect 41412 49980 41422 50036
rect 12226 49868 12236 49924
rect 12292 49868 13132 49924
rect 13188 49868 15148 49924
rect 16482 49868 16492 49924
rect 16548 49868 17276 49924
rect 17332 49868 17342 49924
rect 15092 49812 15148 49868
rect 18732 49812 18788 49980
rect 43036 49924 43092 50092
rect 22082 49868 22092 49924
rect 22148 49868 22876 49924
rect 22932 49868 23660 49924
rect 23716 49868 23726 49924
rect 30706 49868 30716 49924
rect 30772 49868 31164 49924
rect 31220 49868 32172 49924
rect 32228 49868 32238 49924
rect 37090 49868 37100 49924
rect 37156 49868 43092 49924
rect 47618 49868 47628 49924
rect 47684 49868 48748 49924
rect 48804 49868 48814 49924
rect 12898 49756 12908 49812
rect 12964 49756 13804 49812
rect 13860 49756 14364 49812
rect 14420 49756 14430 49812
rect 15092 49756 16380 49812
rect 16436 49756 16446 49812
rect 18162 49756 18172 49812
rect 18228 49756 19516 49812
rect 19572 49756 19582 49812
rect 22418 49756 22428 49812
rect 22484 49756 23100 49812
rect 23156 49756 23166 49812
rect 34850 49756 34860 49812
rect 34916 49756 35644 49812
rect 35700 49756 35710 49812
rect 36194 49756 36204 49812
rect 36260 49756 37548 49812
rect 37604 49756 37614 49812
rect 39106 49756 39116 49812
rect 39172 49756 39900 49812
rect 39956 49756 42028 49812
rect 42084 49756 42094 49812
rect 43026 49756 43036 49812
rect 43092 49756 43932 49812
rect 43988 49756 49084 49812
rect 49140 49756 49150 49812
rect 11218 49644 11228 49700
rect 11284 49644 11676 49700
rect 11732 49644 13916 49700
rect 13972 49644 13982 49700
rect 19618 49644 19628 49700
rect 19684 49644 22988 49700
rect 23044 49644 23054 49700
rect 30482 49644 30492 49700
rect 30548 49644 30828 49700
rect 30884 49644 31276 49700
rect 31332 49644 31342 49700
rect 40674 49644 40684 49700
rect 40740 49644 41244 49700
rect 41300 49644 42924 49700
rect 42980 49644 42990 49700
rect 44482 49644 44492 49700
rect 44548 49644 44940 49700
rect 44996 49644 45388 49700
rect 45444 49644 45454 49700
rect 14802 49532 14812 49588
rect 14868 49532 15820 49588
rect 15876 49532 15886 49588
rect 21186 49532 21196 49588
rect 21252 49532 21868 49588
rect 21924 49532 21934 49588
rect 36642 49532 36652 49588
rect 36708 49532 41356 49588
rect 41412 49532 41422 49588
rect 4834 49420 4844 49476
rect 4900 49420 4910 49476
rect 20514 49420 20524 49476
rect 20580 49420 21084 49476
rect 21140 49420 34300 49476
rect 34356 49420 34366 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 4844 49140 4900 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 22978 49196 22988 49252
rect 23044 49196 24108 49252
rect 24164 49196 26908 49252
rect 26964 49196 26974 49252
rect 30146 49196 30156 49252
rect 30212 49196 36876 49252
rect 36932 49196 36942 49252
rect 39778 49196 39788 49252
rect 39844 49196 41804 49252
rect 41860 49196 43036 49252
rect 43092 49196 43102 49252
rect 46834 49196 46844 49252
rect 46900 49196 49084 49252
rect 49140 49196 49150 49252
rect 49746 49196 49756 49252
rect 49812 49196 50540 49252
rect 50596 49196 50606 49252
rect 3938 49084 3948 49140
rect 4004 49084 5740 49140
rect 5796 49084 5806 49140
rect 18498 49084 18508 49140
rect 18564 49084 19964 49140
rect 20020 49084 20030 49140
rect 20626 49084 20636 49140
rect 20692 49084 21420 49140
rect 21476 49084 21486 49140
rect 27570 49084 27580 49140
rect 27636 49084 28476 49140
rect 28532 49084 29484 49140
rect 29540 49084 30380 49140
rect 30436 49084 30446 49140
rect 49522 49084 49532 49140
rect 49588 49084 49868 49140
rect 49924 49084 49934 49140
rect 4722 48972 4732 49028
rect 4788 48972 5628 49028
rect 5684 48972 6076 49028
rect 6132 48972 7700 49028
rect 8642 48972 8652 49028
rect 8708 48972 11788 49028
rect 11844 48972 11854 49028
rect 12114 48972 12124 49028
rect 12180 48972 16604 49028
rect 16660 48972 16670 49028
rect 17154 48972 17164 49028
rect 17220 48972 20972 49028
rect 21028 48972 21038 49028
rect 27794 48972 27804 49028
rect 27860 48972 29148 49028
rect 29204 48972 29214 49028
rect 31266 48972 31276 49028
rect 31332 48972 33964 49028
rect 34020 48972 34030 49028
rect 36194 48972 36204 49028
rect 36260 48972 37100 49028
rect 37156 48972 37166 49028
rect 37426 48972 37436 49028
rect 37492 48972 38668 49028
rect 39106 48972 39116 49028
rect 39172 48972 39788 49028
rect 39844 48972 39854 49028
rect 7644 48916 7700 48972
rect 38612 48916 38668 48972
rect 4946 48860 4956 48916
rect 5012 48860 5852 48916
rect 5908 48860 7084 48916
rect 7140 48860 7150 48916
rect 7634 48860 7644 48916
rect 7700 48860 7710 48916
rect 9762 48860 9772 48916
rect 9828 48860 11900 48916
rect 11956 48860 13524 48916
rect 14914 48860 14924 48916
rect 14980 48860 19628 48916
rect 19684 48860 19694 48916
rect 20178 48860 20188 48916
rect 20244 48860 21308 48916
rect 21364 48860 21374 48916
rect 23202 48860 23212 48916
rect 23268 48860 23884 48916
rect 23940 48860 25004 48916
rect 25060 48860 25070 48916
rect 28914 48860 28924 48916
rect 28980 48860 31948 48916
rect 32004 48860 32014 48916
rect 33394 48860 33404 48916
rect 33460 48860 34748 48916
rect 34804 48860 34814 48916
rect 34962 48860 34972 48916
rect 35028 48860 36428 48916
rect 36484 48860 36494 48916
rect 37650 48860 37660 48916
rect 37716 48860 38332 48916
rect 38388 48860 38398 48916
rect 38612 48860 39452 48916
rect 39508 48860 39900 48916
rect 39956 48860 39966 48916
rect 13468 48804 13524 48860
rect 34748 48804 34804 48860
rect 2482 48748 2492 48804
rect 2548 48748 4620 48804
rect 4676 48748 4686 48804
rect 6514 48748 6524 48804
rect 6580 48748 7196 48804
rect 7252 48748 7262 48804
rect 13234 48748 13244 48804
rect 13300 48748 13310 48804
rect 13468 48748 15260 48804
rect 15316 48748 15326 48804
rect 16594 48748 16604 48804
rect 16660 48748 25116 48804
rect 25172 48748 25182 48804
rect 28242 48748 28252 48804
rect 28308 48748 29372 48804
rect 29428 48748 29708 48804
rect 29764 48748 29774 48804
rect 34748 48748 35420 48804
rect 35476 48748 35486 48804
rect 36082 48748 36092 48804
rect 36148 48748 37996 48804
rect 38052 48748 38062 48804
rect 13244 48692 13300 48748
rect 13244 48636 16828 48692
rect 16884 48636 16894 48692
rect 26786 48636 26796 48692
rect 26852 48636 27356 48692
rect 27412 48636 27422 48692
rect 43810 48636 43820 48692
rect 43876 48636 44828 48692
rect 44884 48636 47740 48692
rect 47796 48636 47806 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 25666 48524 25676 48580
rect 25732 48524 26012 48580
rect 26068 48524 27580 48580
rect 27636 48524 27646 48580
rect 11330 48412 11340 48468
rect 11396 48412 15148 48468
rect 15204 48412 15214 48468
rect 17490 48412 17500 48468
rect 17556 48412 17836 48468
rect 17892 48412 17902 48468
rect 19394 48412 19404 48468
rect 19460 48412 20412 48468
rect 20468 48412 20478 48468
rect 24658 48412 24668 48468
rect 24724 48412 25788 48468
rect 25844 48412 26460 48468
rect 26516 48412 30940 48468
rect 30996 48412 31006 48468
rect 43362 48412 43372 48468
rect 43428 48412 49644 48468
rect 49700 48412 49710 48468
rect 50642 48412 50652 48468
rect 50708 48412 51324 48468
rect 51380 48412 51390 48468
rect 3042 48300 3052 48356
rect 3108 48300 6972 48356
rect 7028 48300 7868 48356
rect 7924 48300 7934 48356
rect 11666 48300 11676 48356
rect 11732 48300 15596 48356
rect 15652 48300 15662 48356
rect 22642 48300 22652 48356
rect 22708 48300 23772 48356
rect 23828 48300 23838 48356
rect 33170 48300 33180 48356
rect 33236 48300 34076 48356
rect 34132 48300 34142 48356
rect 44034 48300 44044 48356
rect 44100 48300 46060 48356
rect 46116 48300 46126 48356
rect 46946 48300 46956 48356
rect 47012 48300 50540 48356
rect 50596 48300 51436 48356
rect 51492 48300 51502 48356
rect 4050 48188 4060 48244
rect 4116 48188 8092 48244
rect 8148 48188 8158 48244
rect 8642 48188 8652 48244
rect 8708 48188 9772 48244
rect 9828 48188 10892 48244
rect 10948 48188 10958 48244
rect 12898 48188 12908 48244
rect 12964 48188 14700 48244
rect 14756 48188 14766 48244
rect 16034 48188 16044 48244
rect 16100 48188 17276 48244
rect 17332 48188 17342 48244
rect 18386 48188 18396 48244
rect 18452 48188 20748 48244
rect 20804 48188 20814 48244
rect 23090 48188 23100 48244
rect 23156 48188 24332 48244
rect 24388 48188 26012 48244
rect 26068 48188 28700 48244
rect 28756 48188 28766 48244
rect 31826 48188 31836 48244
rect 31892 48188 32508 48244
rect 32564 48188 33292 48244
rect 33348 48188 36204 48244
rect 36260 48188 38668 48244
rect 43362 48188 43372 48244
rect 43428 48188 44156 48244
rect 44212 48188 44222 48244
rect 47954 48188 47964 48244
rect 48020 48188 48636 48244
rect 48692 48188 48702 48244
rect 4956 48132 5012 48188
rect 38612 48132 38668 48188
rect 4946 48076 4956 48132
rect 5012 48076 5022 48132
rect 8754 48076 8764 48132
rect 8820 48076 9884 48132
rect 9940 48076 9950 48132
rect 17938 48076 17948 48132
rect 18004 48076 21420 48132
rect 21476 48076 21486 48132
rect 22726 48076 22764 48132
rect 22820 48076 22830 48132
rect 23538 48076 23548 48132
rect 23604 48076 26684 48132
rect 26740 48076 27916 48132
rect 27972 48076 27982 48132
rect 28354 48076 28364 48132
rect 28420 48076 29148 48132
rect 29204 48076 29214 48132
rect 38612 48076 45388 48132
rect 45444 48076 45454 48132
rect 46386 48076 46396 48132
rect 46452 48076 48860 48132
rect 48916 48076 48926 48132
rect 51538 48076 51548 48132
rect 51604 48076 53340 48132
rect 53396 48076 53406 48132
rect 27916 48020 27972 48076
rect 8978 47964 8988 48020
rect 9044 47964 9996 48020
rect 10052 47964 10062 48020
rect 12338 47964 12348 48020
rect 12404 47964 13356 48020
rect 13412 47964 13422 48020
rect 22978 47964 22988 48020
rect 23044 47964 23660 48020
rect 23716 47964 23726 48020
rect 27916 47964 29260 48020
rect 29316 47964 29326 48020
rect 43250 47964 43260 48020
rect 43316 47964 47292 48020
rect 47348 47964 47358 48020
rect 48178 47964 48188 48020
rect 48244 47964 49756 48020
rect 49812 47964 50652 48020
rect 50708 47964 50718 48020
rect 16818 47852 16828 47908
rect 16884 47852 17836 47908
rect 17892 47852 18172 47908
rect 18228 47852 18238 47908
rect 28690 47852 28700 47908
rect 28756 47852 33068 47908
rect 33124 47852 33134 47908
rect 46498 47852 46508 47908
rect 46564 47852 49084 47908
rect 49140 47852 50092 47908
rect 50148 47852 50158 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 12674 47740 12684 47796
rect 12740 47740 14140 47796
rect 14196 47740 14588 47796
rect 14644 47740 22764 47796
rect 22820 47740 22830 47796
rect 27234 47740 27244 47796
rect 27300 47740 27356 47796
rect 27412 47740 29708 47796
rect 29764 47740 29774 47796
rect 13570 47628 13580 47684
rect 13636 47628 16492 47684
rect 16548 47628 16558 47684
rect 19506 47628 19516 47684
rect 19572 47628 24332 47684
rect 24388 47628 25340 47684
rect 25396 47628 25406 47684
rect 25666 47628 25676 47684
rect 25732 47628 26684 47684
rect 26740 47628 26750 47684
rect 49634 47628 49644 47684
rect 49700 47628 51548 47684
rect 51604 47628 51614 47684
rect 8866 47516 8876 47572
rect 8932 47516 9660 47572
rect 9716 47516 9726 47572
rect 12114 47516 12124 47572
rect 12180 47516 18396 47572
rect 18452 47516 18462 47572
rect 26852 47516 27244 47572
rect 27300 47516 29820 47572
rect 29876 47516 29886 47572
rect 44258 47516 44268 47572
rect 44324 47516 44716 47572
rect 44772 47516 44782 47572
rect 45378 47516 45388 47572
rect 45444 47516 45836 47572
rect 45892 47516 48524 47572
rect 48580 47516 48590 47572
rect 26852 47460 26908 47516
rect 16706 47404 16716 47460
rect 16772 47404 18508 47460
rect 18564 47404 18574 47460
rect 19618 47404 19628 47460
rect 19684 47404 20412 47460
rect 20468 47404 21308 47460
rect 21364 47404 21374 47460
rect 21746 47404 21756 47460
rect 21812 47404 26908 47460
rect 27682 47404 27692 47460
rect 27748 47404 29036 47460
rect 29092 47404 29102 47460
rect 31378 47404 31388 47460
rect 31444 47404 32732 47460
rect 32788 47404 32798 47460
rect 46050 47404 46060 47460
rect 46116 47404 47180 47460
rect 47236 47404 47246 47460
rect 48290 47404 48300 47460
rect 48356 47404 49868 47460
rect 49924 47404 50316 47460
rect 50372 47404 51212 47460
rect 51268 47404 51278 47460
rect 47180 47348 47236 47404
rect 12562 47292 12572 47348
rect 12628 47292 14140 47348
rect 14196 47292 14206 47348
rect 16482 47292 16492 47348
rect 16548 47292 22540 47348
rect 22596 47292 22606 47348
rect 25974 47292 26012 47348
rect 26068 47292 26078 47348
rect 28018 47292 28028 47348
rect 28084 47292 28756 47348
rect 42130 47292 42140 47348
rect 42196 47292 44828 47348
rect 44884 47292 44894 47348
rect 47180 47292 48748 47348
rect 48804 47292 48814 47348
rect 16716 47236 16772 47292
rect 13906 47180 13916 47236
rect 13972 47180 14756 47236
rect 15026 47180 15036 47236
rect 15092 47180 16044 47236
rect 16100 47180 16110 47236
rect 16706 47180 16716 47236
rect 16772 47180 16782 47236
rect 19628 47180 24108 47236
rect 24164 47180 24556 47236
rect 24612 47180 25676 47236
rect 25732 47180 25742 47236
rect 27682 47180 27692 47236
rect 27748 47180 28476 47236
rect 28532 47180 28542 47236
rect 14700 47124 14756 47180
rect 19628 47124 19684 47180
rect 13458 47068 13468 47124
rect 13524 47068 14140 47124
rect 14196 47068 14206 47124
rect 14700 47068 19684 47124
rect 20738 47068 20748 47124
rect 20804 47068 21196 47124
rect 21252 47068 21262 47124
rect 21410 47068 21420 47124
rect 21476 47068 21532 47124
rect 21588 47068 21598 47124
rect 23426 47068 23436 47124
rect 23492 47068 25452 47124
rect 25508 47068 26236 47124
rect 26292 47068 26302 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 28700 47012 28756 47292
rect 33282 47068 33292 47124
rect 33348 47068 33628 47124
rect 33684 47068 33694 47124
rect 39218 47068 39228 47124
rect 39284 47068 43260 47124
rect 43316 47068 44492 47124
rect 44548 47068 44558 47124
rect 46050 47068 46060 47124
rect 46116 47068 48636 47124
rect 48692 47068 48702 47124
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 12898 46956 12908 47012
rect 12964 46956 13580 47012
rect 13636 46956 14364 47012
rect 14420 46956 15708 47012
rect 15764 46956 15774 47012
rect 16034 46956 16044 47012
rect 16100 46956 17164 47012
rect 17220 46956 17230 47012
rect 28700 46956 28924 47012
rect 28980 46956 28990 47012
rect 29260 46956 32508 47012
rect 32564 46956 33068 47012
rect 33124 46956 33134 47012
rect 34402 46956 34412 47012
rect 34468 46956 34748 47012
rect 34804 46956 35756 47012
rect 35812 46956 36316 47012
rect 36372 46956 37100 47012
rect 37156 46956 37772 47012
rect 37828 46956 37838 47012
rect 50978 46956 50988 47012
rect 51044 46956 51660 47012
rect 51716 46956 51726 47012
rect 16044 46900 16100 46956
rect 14578 46844 14588 46900
rect 14644 46844 16100 46900
rect 19730 46844 19740 46900
rect 19796 46844 20748 46900
rect 20804 46844 23100 46900
rect 23156 46844 24108 46900
rect 24164 46844 24174 46900
rect 25106 46844 25116 46900
rect 25172 46844 27132 46900
rect 27188 46844 27198 46900
rect 29260 46788 29316 46956
rect 29474 46844 29484 46900
rect 29540 46844 29708 46900
rect 29764 46844 29774 46900
rect 30146 46844 30156 46900
rect 30212 46844 30828 46900
rect 30884 46844 30894 46900
rect 16258 46732 16268 46788
rect 16324 46732 16716 46788
rect 16772 46732 16782 46788
rect 17714 46732 17724 46788
rect 17780 46732 26908 46788
rect 28578 46732 28588 46788
rect 28644 46732 29260 46788
rect 29316 46732 29326 46788
rect 29586 46732 29596 46788
rect 29652 46732 30940 46788
rect 30996 46732 31006 46788
rect 31154 46732 31164 46788
rect 31220 46732 32396 46788
rect 32452 46732 32462 46788
rect 47394 46732 47404 46788
rect 47460 46732 49084 46788
rect 49140 46732 49150 46788
rect 26852 46676 26908 46732
rect 6402 46620 6412 46676
rect 6468 46620 7532 46676
rect 7588 46620 7598 46676
rect 11554 46620 11564 46676
rect 11620 46620 13132 46676
rect 13188 46620 13198 46676
rect 13346 46620 13356 46676
rect 13412 46620 17948 46676
rect 18004 46620 18014 46676
rect 18946 46620 18956 46676
rect 19012 46620 19292 46676
rect 19348 46620 19358 46676
rect 20850 46620 20860 46676
rect 20916 46620 21756 46676
rect 21812 46620 21822 46676
rect 22092 46620 25340 46676
rect 25396 46620 25406 46676
rect 26852 46620 28028 46676
rect 28084 46620 31052 46676
rect 31108 46620 31118 46676
rect 31266 46620 31276 46676
rect 31332 46620 32060 46676
rect 32116 46620 32126 46676
rect 33954 46620 33964 46676
rect 34020 46620 34412 46676
rect 34468 46620 39676 46676
rect 39732 46620 39742 46676
rect 44930 46620 44940 46676
rect 44996 46620 45836 46676
rect 45892 46620 50540 46676
rect 50596 46620 50606 46676
rect 22092 46564 22148 46620
rect 13682 46508 13692 46564
rect 13748 46508 14476 46564
rect 14532 46508 14542 46564
rect 16370 46508 16380 46564
rect 16436 46508 22148 46564
rect 22306 46508 22316 46564
rect 22372 46508 29484 46564
rect 29540 46508 31724 46564
rect 31780 46508 31790 46564
rect 40226 46508 40236 46564
rect 40292 46508 41692 46564
rect 41748 46508 41758 46564
rect 46162 46508 46172 46564
rect 46228 46508 46620 46564
rect 46676 46508 48860 46564
rect 48916 46508 48926 46564
rect 3378 46396 3388 46452
rect 3444 46396 4284 46452
rect 4340 46396 4350 46452
rect 15810 46396 15820 46452
rect 15876 46396 25004 46452
rect 25060 46396 25070 46452
rect 26786 46396 26796 46452
rect 26852 46396 27580 46452
rect 27636 46396 27646 46452
rect 35970 46396 35980 46452
rect 36036 46396 37100 46452
rect 37156 46396 37166 46452
rect 45714 46396 45724 46452
rect 45780 46396 47292 46452
rect 47348 46396 47358 46452
rect 11778 46284 11788 46340
rect 11844 46284 16604 46340
rect 16660 46284 16670 46340
rect 18722 46284 18732 46340
rect 18788 46284 19516 46340
rect 19572 46284 19582 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 15138 46172 15148 46228
rect 15204 46172 15316 46228
rect 15922 46172 15932 46228
rect 15988 46172 23212 46228
rect 23268 46172 23278 46228
rect 24882 46172 24892 46228
rect 24948 46172 33404 46228
rect 33460 46172 33470 46228
rect 45042 46172 45052 46228
rect 45108 46172 45836 46228
rect 45892 46172 47068 46228
rect 47124 46172 47134 46228
rect 15260 46116 15316 46172
rect 23212 46116 23268 46172
rect 10546 46060 10556 46116
rect 10612 46060 10892 46116
rect 10948 46060 12460 46116
rect 12516 46060 12526 46116
rect 15260 46060 16492 46116
rect 16548 46060 16558 46116
rect 17154 46060 17164 46116
rect 17220 46060 18060 46116
rect 18116 46060 18126 46116
rect 19030 46060 19068 46116
rect 19124 46060 19134 46116
rect 19282 46060 19292 46116
rect 19348 46060 21980 46116
rect 22036 46060 22046 46116
rect 23212 46060 24052 46116
rect 26562 46060 26572 46116
rect 26628 46060 27020 46116
rect 27076 46060 27468 46116
rect 27524 46060 27534 46116
rect 49298 46060 49308 46116
rect 49364 46060 51548 46116
rect 51604 46060 51614 46116
rect 19404 46004 19460 46060
rect 1810 45948 1820 46004
rect 1876 45948 5068 46004
rect 5124 45948 5134 46004
rect 11218 45948 11228 46004
rect 11284 45948 15036 46004
rect 15092 45948 15484 46004
rect 15540 45948 15550 46004
rect 19394 45948 19404 46004
rect 19460 45948 19470 46004
rect 20626 45948 20636 46004
rect 20692 45948 21756 46004
rect 21812 45948 21822 46004
rect 23996 45892 24052 46060
rect 24210 45948 24220 46004
rect 24276 45948 28140 46004
rect 28196 45948 28206 46004
rect 17714 45836 17724 45892
rect 17780 45836 20356 45892
rect 21634 45836 21644 45892
rect 21700 45836 22988 45892
rect 23044 45836 23054 45892
rect 23996 45836 28028 45892
rect 28084 45836 28094 45892
rect 37538 45836 37548 45892
rect 37604 45836 38332 45892
rect 38388 45836 39228 45892
rect 39284 45836 39294 45892
rect 39890 45836 39900 45892
rect 39956 45836 40460 45892
rect 40516 45836 40526 45892
rect 41458 45836 41468 45892
rect 41524 45836 44044 45892
rect 44100 45836 44492 45892
rect 44548 45836 44940 45892
rect 44996 45836 46620 45892
rect 46676 45836 46686 45892
rect 20300 45780 20356 45836
rect 5842 45724 5852 45780
rect 5908 45724 6524 45780
rect 6580 45724 6590 45780
rect 14690 45724 14700 45780
rect 14756 45724 15708 45780
rect 15764 45724 15774 45780
rect 17042 45724 17052 45780
rect 17108 45724 18284 45780
rect 18340 45724 18350 45780
rect 20290 45724 20300 45780
rect 20356 45724 27692 45780
rect 27748 45724 30156 45780
rect 30212 45724 30222 45780
rect 31154 45724 31164 45780
rect 31220 45724 31724 45780
rect 31780 45724 33292 45780
rect 33348 45724 33358 45780
rect 16034 45612 16044 45668
rect 16100 45612 25900 45668
rect 25956 45612 25966 45668
rect 26852 45612 27244 45668
rect 27300 45612 27310 45668
rect 19366 45500 19404 45556
rect 19460 45500 19470 45556
rect 22978 45500 22988 45556
rect 23044 45500 23884 45556
rect 23940 45500 23950 45556
rect 25554 45500 25564 45556
rect 25620 45500 26012 45556
rect 26068 45500 26078 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 26852 45444 26908 45612
rect 31164 45556 31220 45724
rect 30706 45500 30716 45556
rect 30772 45500 31220 45556
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 14466 45388 14476 45444
rect 14532 45388 15036 45444
rect 15092 45388 15102 45444
rect 24658 45388 24668 45444
rect 24724 45388 25676 45444
rect 25732 45388 26908 45444
rect 27010 45388 27020 45444
rect 27076 45388 28252 45444
rect 28308 45388 29372 45444
rect 29428 45388 29438 45444
rect 39554 45388 39564 45444
rect 39620 45388 39630 45444
rect 39564 45332 39620 45388
rect 17154 45276 17164 45332
rect 17220 45276 24332 45332
rect 24388 45276 24398 45332
rect 26338 45276 26348 45332
rect 26404 45276 29148 45332
rect 29204 45276 29214 45332
rect 29372 45276 31276 45332
rect 31332 45276 31342 45332
rect 39526 45276 39564 45332
rect 39620 45276 40348 45332
rect 40404 45276 44380 45332
rect 44436 45276 44446 45332
rect 29372 45220 29428 45276
rect 2258 45164 2268 45220
rect 2324 45164 2492 45220
rect 2548 45164 3500 45220
rect 3556 45164 4060 45220
rect 4116 45164 4126 45220
rect 6402 45164 6412 45220
rect 6468 45164 8652 45220
rect 8708 45164 10556 45220
rect 10612 45164 10622 45220
rect 18834 45164 18844 45220
rect 18900 45164 23996 45220
rect 24052 45164 24062 45220
rect 26786 45164 26796 45220
rect 26852 45164 29428 45220
rect 30034 45164 30044 45220
rect 30100 45164 31388 45220
rect 31444 45164 32284 45220
rect 32340 45164 32350 45220
rect 39554 45164 39564 45220
rect 39620 45164 41468 45220
rect 41524 45164 42364 45220
rect 42420 45164 42430 45220
rect 2706 45052 2716 45108
rect 2772 45052 3948 45108
rect 4004 45052 4620 45108
rect 4676 45052 4956 45108
rect 5012 45052 5022 45108
rect 11106 45052 11116 45108
rect 11172 45052 12012 45108
rect 12068 45052 12078 45108
rect 12562 45052 12572 45108
rect 12628 45052 14364 45108
rect 14420 45052 14430 45108
rect 17266 45052 17276 45108
rect 17332 45052 17612 45108
rect 17668 45052 17678 45108
rect 17938 45052 17948 45108
rect 18004 45052 19068 45108
rect 19124 45052 19134 45108
rect 23426 45052 23436 45108
rect 23492 45052 23884 45108
rect 23940 45052 23950 45108
rect 26674 45052 26684 45108
rect 26740 45052 29260 45108
rect 29316 45052 29820 45108
rect 29876 45052 29886 45108
rect 30930 45052 30940 45108
rect 30996 45052 33964 45108
rect 34020 45052 34030 45108
rect 41570 45052 41580 45108
rect 41636 45052 42476 45108
rect 42532 45052 42542 45108
rect 12012 44996 12068 45052
rect 11218 44940 11228 44996
rect 11284 44940 11788 44996
rect 11844 44940 11854 44996
rect 12012 44940 12908 44996
rect 12964 44940 12974 44996
rect 15092 44940 18620 44996
rect 18676 44940 18686 44996
rect 20290 44940 20300 44996
rect 20356 44940 22092 44996
rect 22148 44940 22158 44996
rect 34178 44940 34188 44996
rect 34244 44940 35420 44996
rect 35476 44940 35486 44996
rect 51650 44940 51660 44996
rect 51716 44940 52332 44996
rect 52388 44940 52398 44996
rect 15092 44884 15148 44940
rect 10658 44828 10668 44884
rect 10724 44828 15148 44884
rect 16370 44828 16380 44884
rect 16436 44828 17948 44884
rect 18004 44828 19292 44884
rect 19348 44828 19358 44884
rect 27234 44828 27244 44884
rect 27300 44828 28476 44884
rect 28532 44828 28542 44884
rect 33394 44828 33404 44884
rect 33460 44828 33740 44884
rect 33796 44828 33806 44884
rect 39666 44828 39676 44884
rect 39732 44828 42364 44884
rect 42420 44828 42430 44884
rect 27244 44772 27300 44828
rect 17350 44716 17388 44772
rect 17444 44716 17454 44772
rect 19058 44716 19068 44772
rect 19124 44716 27300 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 16818 44604 16828 44660
rect 16884 44604 17724 44660
rect 17780 44604 19852 44660
rect 19908 44604 19918 44660
rect 26898 44604 26908 44660
rect 26964 44604 31612 44660
rect 31668 44604 32508 44660
rect 32564 44604 32574 44660
rect 36866 44604 36876 44660
rect 36932 44604 44828 44660
rect 44884 44604 44894 44660
rect 3378 44492 3388 44548
rect 3444 44492 3668 44548
rect 8754 44492 8764 44548
rect 8820 44492 10108 44548
rect 10164 44492 10174 44548
rect 10994 44492 11004 44548
rect 11060 44492 11452 44548
rect 11508 44492 12572 44548
rect 12628 44492 12638 44548
rect 14140 44492 17276 44548
rect 17332 44492 17342 44548
rect 28578 44492 28588 44548
rect 28644 44492 29596 44548
rect 29652 44492 31276 44548
rect 31332 44492 32956 44548
rect 33012 44492 33516 44548
rect 33572 44492 33582 44548
rect 3612 44100 3668 44492
rect 5954 44380 5964 44436
rect 6020 44380 6030 44436
rect 7298 44380 7308 44436
rect 7364 44380 8540 44436
rect 8596 44380 8606 44436
rect 10210 44380 10220 44436
rect 10276 44380 11788 44436
rect 11844 44380 13468 44436
rect 13524 44380 13534 44436
rect 5964 44100 6020 44380
rect 10658 44268 10668 44324
rect 10724 44268 13692 44324
rect 13748 44268 13758 44324
rect 14140 44212 14196 44492
rect 17042 44380 17052 44436
rect 17108 44380 18172 44436
rect 18228 44380 18238 44436
rect 24994 44380 25004 44436
rect 25060 44380 28364 44436
rect 28420 44380 28430 44436
rect 32834 44380 32844 44436
rect 32900 44380 33740 44436
rect 33796 44380 33806 44436
rect 14466 44268 14476 44324
rect 14532 44268 17948 44324
rect 18004 44268 18014 44324
rect 18274 44268 18284 44324
rect 18340 44268 18956 44324
rect 19012 44268 19022 44324
rect 20066 44268 20076 44324
rect 20132 44268 20524 44324
rect 20580 44268 20590 44324
rect 24210 44268 24220 44324
rect 24276 44268 27356 44324
rect 27412 44268 27422 44324
rect 28242 44268 28252 44324
rect 28308 44268 31276 44324
rect 31332 44268 31342 44324
rect 32386 44268 32396 44324
rect 32452 44268 33404 44324
rect 33460 44268 33470 44324
rect 33740 44268 36092 44324
rect 36148 44268 36158 44324
rect 37986 44268 37996 44324
rect 38052 44268 38780 44324
rect 38836 44268 39788 44324
rect 39844 44268 39854 44324
rect 33740 44212 33796 44268
rect 13234 44156 13244 44212
rect 13300 44156 14140 44212
rect 14196 44156 14206 44212
rect 14354 44156 14364 44212
rect 14420 44156 14924 44212
rect 14980 44156 15484 44212
rect 15540 44156 15932 44212
rect 15988 44156 33796 44212
rect 33954 44156 33964 44212
rect 34020 44156 38444 44212
rect 38500 44156 39116 44212
rect 39172 44156 39182 44212
rect 3602 44044 3612 44100
rect 3668 44044 5068 44100
rect 5124 44044 5134 44100
rect 5282 44044 5292 44100
rect 5348 44044 6020 44100
rect 11116 44044 11676 44100
rect 11732 44044 12012 44100
rect 12068 44044 12078 44100
rect 12338 44044 12348 44100
rect 12404 44044 13804 44100
rect 13860 44044 13870 44100
rect 18834 44044 18844 44100
rect 18900 44044 19740 44100
rect 19796 44044 20636 44100
rect 20692 44044 22988 44100
rect 23044 44044 23054 44100
rect 25890 44044 25900 44100
rect 25956 44044 26908 44100
rect 29922 44044 29932 44100
rect 29988 44044 31052 44100
rect 31108 44044 31118 44100
rect 33394 44044 33404 44100
rect 33460 44044 34076 44100
rect 34132 44044 34142 44100
rect 34626 44044 34636 44100
rect 34692 44044 38668 44100
rect 39218 44044 39228 44100
rect 39284 44044 40124 44100
rect 40180 44044 41804 44100
rect 41860 44044 44156 44100
rect 44212 44044 45836 44100
rect 45892 44044 45902 44100
rect 48178 44044 48188 44100
rect 48244 44044 49084 44100
rect 49140 44044 49150 44100
rect 11116 43876 11172 44044
rect 13010 43932 13020 43988
rect 13076 43932 14476 43988
rect 14532 43932 14542 43988
rect 19282 43932 19292 43988
rect 19348 43932 19684 43988
rect 26226 43932 26236 43988
rect 26292 43932 26684 43988
rect 26740 43932 26750 43988
rect 8978 43820 8988 43876
rect 9044 43820 10332 43876
rect 10388 43820 11116 43876
rect 11172 43820 11182 43876
rect 11778 43820 11788 43876
rect 11844 43820 14700 43876
rect 14756 43820 14766 43876
rect 15138 43820 15148 43876
rect 15204 43820 17724 43876
rect 17780 43820 17790 43876
rect 18274 43820 18284 43876
rect 18340 43820 19404 43876
rect 19460 43820 19470 43876
rect 19628 43764 19684 43932
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 25778 43820 25788 43876
rect 25844 43820 26572 43876
rect 26628 43820 26638 43876
rect 26786 43820 26796 43876
rect 26852 43820 26908 44044
rect 34076 43988 34132 44044
rect 27318 43932 27356 43988
rect 27412 43932 27422 43988
rect 27794 43932 27804 43988
rect 27860 43932 30044 43988
rect 30100 43932 30110 43988
rect 34076 43932 34524 43988
rect 34580 43932 34590 43988
rect 28130 43820 28140 43876
rect 28196 43820 30156 43876
rect 30212 43820 30222 43876
rect 38612 43820 38668 44044
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 38724 43820 39900 43876
rect 39956 43820 39966 43876
rect 4610 43708 4620 43764
rect 4676 43708 4956 43764
rect 5012 43708 5022 43764
rect 5618 43708 5628 43764
rect 5684 43708 5694 43764
rect 14018 43708 14028 43764
rect 14084 43708 14094 43764
rect 17378 43708 17388 43764
rect 17444 43708 19292 43764
rect 19348 43708 19358 43764
rect 19628 43708 21196 43764
rect 21252 43708 22204 43764
rect 22260 43708 22270 43764
rect 22418 43708 22428 43764
rect 22484 43708 26908 43764
rect 26964 43708 27916 43764
rect 27972 43708 27982 43764
rect 30594 43708 30604 43764
rect 30660 43708 32172 43764
rect 32228 43708 32238 43764
rect 39526 43708 39564 43764
rect 39620 43708 39630 43764
rect 5628 43652 5684 43708
rect 14028 43652 14084 43708
rect 4834 43596 4844 43652
rect 4900 43596 7420 43652
rect 7476 43596 9548 43652
rect 9604 43596 9614 43652
rect 10882 43596 10892 43652
rect 10948 43596 11228 43652
rect 11284 43596 11294 43652
rect 13346 43596 13356 43652
rect 13412 43596 15260 43652
rect 15316 43596 15326 43652
rect 18386 43596 18396 43652
rect 18452 43596 19964 43652
rect 20020 43596 24220 43652
rect 24276 43596 24286 43652
rect 25442 43596 25452 43652
rect 25508 43596 27020 43652
rect 27076 43596 27086 43652
rect 28130 43596 28140 43652
rect 28196 43596 29708 43652
rect 29764 43596 29774 43652
rect 36978 43596 36988 43652
rect 37044 43596 37772 43652
rect 37828 43596 40348 43652
rect 40404 43596 40414 43652
rect 44818 43596 44828 43652
rect 44884 43596 46844 43652
rect 46900 43596 46910 43652
rect 3378 43484 3388 43540
rect 3444 43484 5516 43540
rect 5572 43484 5582 43540
rect 6626 43484 6636 43540
rect 6692 43484 9100 43540
rect 9156 43484 9166 43540
rect 13122 43484 13132 43540
rect 13188 43484 13692 43540
rect 13748 43484 16268 43540
rect 16324 43484 16334 43540
rect 16930 43484 16940 43540
rect 16996 43484 18060 43540
rect 18116 43484 18126 43540
rect 19394 43484 19404 43540
rect 19460 43484 20636 43540
rect 20692 43484 20702 43540
rect 23202 43484 23212 43540
rect 23268 43484 26348 43540
rect 26404 43484 26414 43540
rect 26852 43484 28476 43540
rect 28532 43484 28542 43540
rect 28914 43484 28924 43540
rect 28980 43484 30268 43540
rect 30324 43484 30334 43540
rect 38434 43484 38444 43540
rect 38500 43484 38892 43540
rect 38948 43484 38958 43540
rect 41234 43484 41244 43540
rect 41300 43484 42140 43540
rect 42196 43484 43260 43540
rect 43316 43484 43326 43540
rect 26852 43428 26908 43484
rect 4722 43372 4732 43428
rect 4788 43372 5628 43428
rect 5684 43372 10220 43428
rect 10276 43372 10286 43428
rect 17154 43372 17164 43428
rect 17220 43372 17500 43428
rect 17556 43372 20860 43428
rect 20916 43372 20926 43428
rect 21858 43372 21868 43428
rect 21924 43372 24220 43428
rect 24276 43372 24286 43428
rect 24546 43372 24556 43428
rect 24612 43372 26908 43428
rect 27122 43372 27132 43428
rect 27188 43372 28700 43428
rect 28756 43372 28766 43428
rect 34738 43372 34748 43428
rect 34804 43372 35868 43428
rect 35924 43372 35934 43428
rect 39890 43372 39900 43428
rect 39956 43372 41468 43428
rect 41524 43372 41534 43428
rect 45378 43372 45388 43428
rect 45444 43372 46172 43428
rect 46228 43372 46238 43428
rect 48738 43372 48748 43428
rect 48804 43372 51100 43428
rect 51156 43372 51166 43428
rect 5842 43260 5852 43316
rect 5908 43260 7532 43316
rect 7588 43260 7598 43316
rect 8642 43260 8652 43316
rect 8708 43260 11676 43316
rect 11732 43260 11742 43316
rect 16706 43260 16716 43316
rect 16772 43260 17276 43316
rect 17332 43260 17342 43316
rect 18582 43260 18620 43316
rect 18676 43260 18686 43316
rect 25330 43260 25340 43316
rect 25396 43260 25788 43316
rect 25844 43260 26796 43316
rect 26852 43260 26862 43316
rect 28802 43260 28812 43316
rect 28868 43260 34524 43316
rect 34580 43260 34590 43316
rect 38546 43260 38556 43316
rect 38612 43260 40236 43316
rect 40292 43260 40796 43316
rect 40852 43260 40862 43316
rect 46050 43260 46060 43316
rect 46116 43260 47292 43316
rect 47348 43260 47358 43316
rect 51650 43260 51660 43316
rect 51716 43260 53788 43316
rect 53844 43260 53854 43316
rect 11442 43148 11452 43204
rect 11508 43148 12684 43204
rect 12740 43148 13692 43204
rect 13748 43148 13758 43204
rect 17266 43148 17276 43204
rect 17332 43148 18844 43204
rect 18900 43148 20524 43204
rect 20580 43148 23548 43204
rect 23604 43148 24892 43204
rect 24948 43148 24958 43204
rect 25106 43148 25116 43204
rect 25172 43148 25676 43204
rect 25732 43148 25742 43204
rect 28578 43148 28588 43204
rect 28644 43148 31164 43204
rect 31220 43148 31230 43204
rect 51286 43148 51324 43204
rect 51380 43148 51390 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 10210 43036 10220 43092
rect 10276 43036 21868 43092
rect 21924 43036 21934 43092
rect 22092 43036 24388 43092
rect 24658 43036 24668 43092
rect 24724 43036 26012 43092
rect 26068 43036 27468 43092
rect 27524 43036 27534 43092
rect 22092 42980 22148 43036
rect 24332 42980 24388 43036
rect 16034 42924 16044 42980
rect 16100 42924 22148 42980
rect 23538 42924 23548 42980
rect 23604 42924 24108 42980
rect 24164 42924 24174 42980
rect 24332 42924 27356 42980
rect 27412 42924 27422 42980
rect 45238 42924 45276 42980
rect 45332 42924 45342 42980
rect 14018 42812 14028 42868
rect 14084 42812 14812 42868
rect 14868 42812 14878 42868
rect 16594 42812 16604 42868
rect 16660 42812 17052 42868
rect 17108 42812 17948 42868
rect 18004 42812 18014 42868
rect 23762 42812 23772 42868
rect 23828 42812 27916 42868
rect 27972 42812 29148 42868
rect 29204 42812 29708 42868
rect 29764 42812 29774 42868
rect 38994 42812 39004 42868
rect 39060 42812 41132 42868
rect 41188 42812 41198 42868
rect 46610 42812 46620 42868
rect 46676 42812 50428 42868
rect 12786 42700 12796 42756
rect 12852 42700 14140 42756
rect 14196 42700 14206 42756
rect 16258 42700 16268 42756
rect 16324 42700 17724 42756
rect 17780 42700 17790 42756
rect 19842 42700 19852 42756
rect 19908 42700 21308 42756
rect 21364 42700 21374 42756
rect 25442 42700 25452 42756
rect 25508 42700 26124 42756
rect 26180 42700 26460 42756
rect 26516 42700 27132 42756
rect 27188 42700 27198 42756
rect 29474 42700 29484 42756
rect 29540 42700 34748 42756
rect 34804 42700 34814 42756
rect 38770 42700 38780 42756
rect 38836 42700 40348 42756
rect 40404 42700 40414 42756
rect 46274 42700 46284 42756
rect 46340 42700 47404 42756
rect 47460 42700 48188 42756
rect 48244 42700 48254 42756
rect 50372 42700 50428 42812
rect 50484 42700 50494 42756
rect 5618 42588 5628 42644
rect 5684 42588 6412 42644
rect 6468 42588 6478 42644
rect 16146 42588 16156 42644
rect 16212 42588 16716 42644
rect 16772 42588 17164 42644
rect 17220 42588 17276 42644
rect 17332 42588 17342 42644
rect 17490 42588 17500 42644
rect 17556 42588 18508 42644
rect 18564 42588 18574 42644
rect 23202 42588 23212 42644
rect 23268 42588 23660 42644
rect 23716 42588 23726 42644
rect 24434 42588 24444 42644
rect 24500 42588 26236 42644
rect 26292 42588 26302 42644
rect 27570 42588 27580 42644
rect 27636 42588 28476 42644
rect 28532 42588 28542 42644
rect 39890 42588 39900 42644
rect 39956 42588 46844 42644
rect 46900 42588 49084 42644
rect 49140 42588 49150 42644
rect 49746 42588 49756 42644
rect 49812 42588 51660 42644
rect 51716 42588 51726 42644
rect 50988 42532 51044 42588
rect 12002 42476 12012 42532
rect 12068 42476 13356 42532
rect 13412 42476 13422 42532
rect 17714 42476 17724 42532
rect 17780 42476 19404 42532
rect 19460 42476 19470 42532
rect 22082 42476 22092 42532
rect 22148 42476 26012 42532
rect 26068 42476 26078 42532
rect 34962 42476 34972 42532
rect 35028 42476 40124 42532
rect 40180 42476 40190 42532
rect 50306 42476 50316 42532
rect 50372 42476 50764 42532
rect 50820 42476 50830 42532
rect 50978 42476 50988 42532
rect 51044 42476 51054 42532
rect 15362 42364 15372 42420
rect 15428 42364 16044 42420
rect 16100 42364 16110 42420
rect 18050 42364 18060 42420
rect 18116 42364 19180 42420
rect 19236 42364 19246 42420
rect 22194 42364 22204 42420
rect 22260 42364 28028 42420
rect 28084 42364 28364 42420
rect 28420 42364 29932 42420
rect 29988 42364 31388 42420
rect 31444 42364 31454 42420
rect 38612 42364 44380 42420
rect 44436 42364 44446 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 38612 42308 38668 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 16268 42252 16940 42308
rect 16996 42252 17006 42308
rect 18834 42252 18844 42308
rect 18900 42252 18938 42308
rect 19282 42252 19292 42308
rect 19348 42252 19628 42308
rect 19684 42252 19694 42308
rect 26852 42252 34188 42308
rect 34244 42252 35644 42308
rect 35700 42252 38668 42308
rect 41794 42252 41804 42308
rect 41860 42252 45612 42308
rect 45668 42252 45678 42308
rect 14354 42140 14364 42196
rect 14420 42140 15260 42196
rect 15316 42140 15326 42196
rect 8866 42028 8876 42084
rect 8932 42028 13804 42084
rect 13860 42028 13870 42084
rect 14466 42028 14476 42084
rect 14532 42028 14924 42084
rect 14980 42028 14990 42084
rect 16268 41972 16324 42252
rect 17378 42140 17388 42196
rect 17444 42140 18564 42196
rect 21074 42140 21084 42196
rect 21140 42140 22316 42196
rect 22372 42140 22382 42196
rect 18508 42084 18564 42140
rect 17388 42028 17948 42084
rect 18004 42028 18014 42084
rect 18498 42028 18508 42084
rect 18564 42028 19068 42084
rect 19124 42028 19134 42084
rect 19282 42028 19292 42084
rect 19348 42028 20188 42084
rect 20244 42028 20254 42084
rect 21970 42028 21980 42084
rect 22036 42028 23604 42084
rect 17388 41972 17444 42028
rect 23548 41972 23604 42028
rect 26852 41972 26908 42252
rect 27458 42140 27468 42196
rect 27524 42140 28364 42196
rect 28420 42140 28430 42196
rect 31266 42140 31276 42196
rect 31332 42140 32284 42196
rect 32340 42140 35196 42196
rect 35252 42140 35262 42196
rect 36194 42140 36204 42196
rect 36260 42140 37772 42196
rect 37828 42140 37838 42196
rect 27122 42028 27132 42084
rect 27188 42028 30828 42084
rect 30884 42028 30894 42084
rect 32050 42028 32060 42084
rect 32116 42028 32620 42084
rect 32676 42028 34748 42084
rect 34804 42028 34814 42084
rect 35522 42028 35532 42084
rect 35588 42028 36988 42084
rect 37044 42028 37054 42084
rect 40114 42028 40124 42084
rect 40180 42028 46620 42084
rect 46676 42028 46686 42084
rect 51874 42028 51884 42084
rect 51940 42028 53004 42084
rect 53060 42028 53070 42084
rect 2818 41916 2828 41972
rect 2884 41916 3724 41972
rect 3780 41916 3790 41972
rect 4050 41916 4060 41972
rect 4116 41916 4732 41972
rect 4788 41916 5292 41972
rect 5348 41916 5964 41972
rect 6020 41916 6030 41972
rect 8754 41916 8764 41972
rect 8820 41916 9100 41972
rect 9156 41916 9660 41972
rect 9716 41916 9726 41972
rect 11442 41916 11452 41972
rect 11508 41916 12236 41972
rect 12292 41916 12302 41972
rect 16258 41916 16268 41972
rect 16324 41916 16334 41972
rect 16930 41916 16940 41972
rect 16996 41916 17444 41972
rect 18162 41916 18172 41972
rect 18228 41916 18956 41972
rect 19012 41916 19022 41972
rect 20290 41916 20300 41972
rect 20356 41916 21140 41972
rect 21522 41916 21532 41972
rect 21588 41916 21868 41972
rect 21924 41916 23324 41972
rect 23380 41916 23390 41972
rect 23548 41916 26908 41972
rect 30370 41916 30380 41972
rect 30436 41916 30940 41972
rect 30996 41916 31006 41972
rect 31938 41916 31948 41972
rect 32004 41916 33068 41972
rect 33124 41916 33134 41972
rect 33282 41916 33292 41972
rect 33348 41916 33516 41972
rect 33572 41916 33582 41972
rect 35074 41916 35084 41972
rect 35140 41916 35868 41972
rect 35924 41916 35934 41972
rect 43026 41916 43036 41972
rect 43092 41916 44044 41972
rect 44100 41916 44110 41972
rect 52210 41916 52220 41972
rect 52276 41916 53676 41972
rect 53732 41916 53742 41972
rect 3154 41804 3164 41860
rect 3220 41804 3948 41860
rect 4004 41804 4014 41860
rect 13458 41804 13468 41860
rect 13524 41804 16380 41860
rect 16436 41804 16446 41860
rect 19954 41804 19964 41860
rect 20020 41804 20524 41860
rect 20580 41804 20590 41860
rect 21084 41748 21140 41916
rect 22754 41804 22764 41860
rect 22820 41804 22830 41860
rect 26786 41804 26796 41860
rect 26852 41804 27244 41860
rect 27300 41804 27692 41860
rect 27748 41804 27758 41860
rect 29586 41804 29596 41860
rect 29652 41804 35756 41860
rect 35812 41804 35822 41860
rect 38322 41804 38332 41860
rect 38388 41804 39900 41860
rect 39956 41804 48748 41860
rect 48804 41804 48814 41860
rect 22764 41748 22820 41804
rect 14802 41692 14812 41748
rect 14868 41692 15260 41748
rect 15316 41692 15326 41748
rect 20738 41692 20748 41748
rect 20804 41692 22820 41748
rect 23538 41692 23548 41748
rect 23604 41692 28588 41748
rect 28644 41692 30044 41748
rect 30100 41692 30110 41748
rect 32162 41692 32172 41748
rect 32228 41692 33068 41748
rect 33124 41692 33134 41748
rect 35298 41692 35308 41748
rect 35364 41692 38668 41748
rect 46050 41692 46060 41748
rect 46116 41692 49420 41748
rect 49476 41692 51996 41748
rect 52052 41692 52780 41748
rect 52836 41692 52846 41748
rect 38612 41636 38668 41692
rect 13346 41580 13356 41636
rect 13412 41580 13916 41636
rect 13972 41580 13982 41636
rect 16258 41580 16268 41636
rect 16324 41580 19964 41636
rect 20020 41580 21644 41636
rect 21700 41580 21710 41636
rect 23650 41580 23660 41636
rect 23716 41580 23884 41636
rect 23940 41580 26012 41636
rect 26068 41580 26078 41636
rect 30258 41580 30268 41636
rect 30324 41580 30604 41636
rect 30660 41580 30670 41636
rect 38612 41580 39340 41636
rect 39396 41580 39406 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 22530 41468 22540 41524
rect 22596 41468 31948 41524
rect 32004 41468 32014 41524
rect 5618 41356 5628 41412
rect 5684 41356 6860 41412
rect 6916 41356 6926 41412
rect 15586 41356 15596 41412
rect 15652 41356 16044 41412
rect 16100 41356 16492 41412
rect 16548 41356 16558 41412
rect 22614 41356 22652 41412
rect 22708 41356 22718 41412
rect 26226 41356 26236 41412
rect 26292 41356 26908 41412
rect 26964 41356 26974 41412
rect 27570 41356 27580 41412
rect 27636 41356 30828 41412
rect 30884 41356 31836 41412
rect 31892 41356 31902 41412
rect 34850 41356 34860 41412
rect 34916 41356 38332 41412
rect 38388 41356 38398 41412
rect 49970 41356 49980 41412
rect 50036 41356 51324 41412
rect 51380 41356 51390 41412
rect 14242 41244 14252 41300
rect 14308 41244 15764 41300
rect 16146 41244 16156 41300
rect 16212 41244 17388 41300
rect 17444 41244 17454 41300
rect 22194 41244 22204 41300
rect 22260 41244 23100 41300
rect 23156 41244 23324 41300
rect 23380 41244 23390 41300
rect 24098 41244 24108 41300
rect 24164 41244 25788 41300
rect 25844 41244 25854 41300
rect 32050 41244 32060 41300
rect 32116 41244 35084 41300
rect 35140 41244 36204 41300
rect 36260 41244 37100 41300
rect 37156 41244 37166 41300
rect 6178 41132 6188 41188
rect 6244 41132 6972 41188
rect 7028 41132 7038 41188
rect 15334 41132 15372 41188
rect 15428 41132 15438 41188
rect 15708 41076 15764 41244
rect 17938 41132 17948 41188
rect 18004 41132 21308 41188
rect 21364 41132 21374 41188
rect 21970 41132 21980 41188
rect 22036 41132 22876 41188
rect 22932 41132 22942 41188
rect 26562 41132 26572 41188
rect 26628 41132 26908 41188
rect 33506 41132 33516 41188
rect 33572 41132 34636 41188
rect 34692 41132 36092 41188
rect 36148 41132 36158 41188
rect 42018 41132 42028 41188
rect 42084 41132 43372 41188
rect 43428 41132 43438 41188
rect 26852 41076 26908 41132
rect 5842 41020 5852 41076
rect 5908 41020 6636 41076
rect 6692 41020 7084 41076
rect 7140 41020 7150 41076
rect 14914 41020 14924 41076
rect 14980 41020 15484 41076
rect 15540 41020 15550 41076
rect 15698 41020 15708 41076
rect 15764 41020 16156 41076
rect 16212 41020 16222 41076
rect 21746 41020 21756 41076
rect 21812 41020 23436 41076
rect 23492 41020 23502 41076
rect 26852 41020 29484 41076
rect 29540 41020 29550 41076
rect 34962 41020 34972 41076
rect 35028 41020 36652 41076
rect 36708 41020 36718 41076
rect 37202 41020 37212 41076
rect 37268 41020 39116 41076
rect 39172 41020 39788 41076
rect 39844 41020 39854 41076
rect 41570 41020 41580 41076
rect 41636 41020 44268 41076
rect 44324 41020 44334 41076
rect 48850 41020 48860 41076
rect 48916 41020 49980 41076
rect 50036 41020 50046 41076
rect 12562 40908 12572 40964
rect 12628 40908 15148 40964
rect 15362 40908 15372 40964
rect 15428 40908 16268 40964
rect 16324 40908 16334 40964
rect 19058 40908 19068 40964
rect 19124 40908 21644 40964
rect 21700 40908 22092 40964
rect 22148 40908 22158 40964
rect 24994 40908 25004 40964
rect 25060 40908 25340 40964
rect 25396 40908 25406 40964
rect 28578 40908 28588 40964
rect 28644 40908 30268 40964
rect 30324 40908 30334 40964
rect 38098 40908 38108 40964
rect 38164 40908 38668 40964
rect 38882 40908 38892 40964
rect 38948 40908 39340 40964
rect 39396 40908 41692 40964
rect 41748 40908 42476 40964
rect 42532 40908 42542 40964
rect 43698 40908 43708 40964
rect 43764 40908 44156 40964
rect 44212 40908 44222 40964
rect 50754 40908 50764 40964
rect 50820 40908 51884 40964
rect 51940 40908 51950 40964
rect 15092 40852 15148 40908
rect 38612 40852 38668 40908
rect 15092 40796 17108 40852
rect 38612 40796 44828 40852
rect 44884 40796 44894 40852
rect 14354 40684 14364 40740
rect 14420 40684 14812 40740
rect 14868 40684 16828 40740
rect 16884 40684 16894 40740
rect 17052 40628 17108 40796
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 37090 40684 37100 40740
rect 37156 40684 37884 40740
rect 37940 40684 37950 40740
rect 44370 40684 44380 40740
rect 44436 40684 45948 40740
rect 46004 40684 46844 40740
rect 46900 40684 46910 40740
rect 2482 40572 2492 40628
rect 2548 40572 4508 40628
rect 4564 40572 4574 40628
rect 8978 40572 8988 40628
rect 9044 40572 9548 40628
rect 9604 40572 9614 40628
rect 13906 40572 13916 40628
rect 13972 40572 15148 40628
rect 15250 40572 15260 40628
rect 15316 40572 15708 40628
rect 15764 40572 15774 40628
rect 17042 40572 17052 40628
rect 17108 40572 18284 40628
rect 18340 40572 18396 40628
rect 18452 40572 18462 40628
rect 18722 40572 18732 40628
rect 18788 40572 19404 40628
rect 19460 40572 19470 40628
rect 19618 40572 19628 40628
rect 19684 40572 19740 40628
rect 19796 40572 22428 40628
rect 22484 40572 22494 40628
rect 24658 40572 24668 40628
rect 24724 40572 26236 40628
rect 26292 40572 26302 40628
rect 32274 40572 32284 40628
rect 32340 40572 38444 40628
rect 38500 40572 38510 40628
rect 41906 40572 41916 40628
rect 41972 40572 45052 40628
rect 45108 40572 45118 40628
rect 48178 40572 48188 40628
rect 48244 40572 49196 40628
rect 49252 40572 49262 40628
rect 50988 40572 52556 40628
rect 52612 40572 52622 40628
rect 15092 40516 15148 40572
rect 50988 40516 51044 40572
rect 6514 40460 6524 40516
rect 6580 40460 7756 40516
rect 7812 40460 7822 40516
rect 10322 40460 10332 40516
rect 10388 40460 13580 40516
rect 13636 40460 13646 40516
rect 15092 40460 15316 40516
rect 15474 40460 15484 40516
rect 15540 40460 19516 40516
rect 19572 40460 22316 40516
rect 22372 40460 22382 40516
rect 39778 40460 39788 40516
rect 39844 40460 43820 40516
rect 43876 40460 43886 40516
rect 49410 40460 49420 40516
rect 49476 40460 50988 40516
rect 51044 40460 51054 40516
rect 51314 40460 51324 40516
rect 51380 40460 51884 40516
rect 51940 40460 51950 40516
rect 15260 40404 15316 40460
rect 4834 40348 4844 40404
rect 4900 40348 6412 40404
rect 6468 40348 6478 40404
rect 13122 40348 13132 40404
rect 13188 40348 13916 40404
rect 13972 40348 15204 40404
rect 15260 40348 22876 40404
rect 22932 40348 22942 40404
rect 26450 40348 26460 40404
rect 26516 40348 29148 40404
rect 29204 40348 29214 40404
rect 29362 40348 29372 40404
rect 29428 40348 30604 40404
rect 30660 40348 30670 40404
rect 37314 40348 37324 40404
rect 37380 40348 39004 40404
rect 39060 40348 39070 40404
rect 39218 40348 39228 40404
rect 39284 40348 41356 40404
rect 41412 40348 41422 40404
rect 49420 40348 49756 40404
rect 49812 40348 49822 40404
rect 50194 40348 50204 40404
rect 50260 40348 50764 40404
rect 50820 40348 51324 40404
rect 51380 40348 51660 40404
rect 51716 40348 51726 40404
rect 15148 40292 15204 40348
rect 26908 40292 26964 40348
rect 39228 40292 39284 40348
rect 49420 40292 49476 40348
rect 4610 40236 4620 40292
rect 4676 40236 5516 40292
rect 5572 40236 5964 40292
rect 6020 40236 6030 40292
rect 15148 40236 15372 40292
rect 15428 40236 15438 40292
rect 17602 40236 17612 40292
rect 17668 40236 18508 40292
rect 18564 40236 18574 40292
rect 20178 40236 20188 40292
rect 20244 40236 20636 40292
rect 20692 40236 21420 40292
rect 21476 40236 22092 40292
rect 22148 40236 22158 40292
rect 26898 40236 26908 40292
rect 26964 40236 26974 40292
rect 28354 40236 28364 40292
rect 28420 40236 29596 40292
rect 29652 40236 29662 40292
rect 29810 40236 29820 40292
rect 29876 40236 32508 40292
rect 32564 40236 32574 40292
rect 37874 40236 37884 40292
rect 37940 40236 39284 40292
rect 42802 40236 42812 40292
rect 42868 40236 44044 40292
rect 44100 40236 45052 40292
rect 45108 40236 45612 40292
rect 45668 40236 45678 40292
rect 46946 40236 46956 40292
rect 47012 40236 47740 40292
rect 47796 40236 47806 40292
rect 49074 40236 49084 40292
rect 49140 40236 49476 40292
rect 49634 40236 49644 40292
rect 49700 40236 49710 40292
rect 50082 40236 50092 40292
rect 50148 40236 50876 40292
rect 50932 40236 50942 40292
rect 15586 40124 15596 40180
rect 15652 40124 18284 40180
rect 18340 40124 18620 40180
rect 18676 40124 18686 40180
rect 19170 40124 19180 40180
rect 19236 40124 19516 40180
rect 19572 40124 19582 40180
rect 23846 40124 23884 40180
rect 23940 40124 23950 40180
rect 26674 40124 26684 40180
rect 26740 40124 29036 40180
rect 29092 40124 29102 40180
rect 34178 40124 34188 40180
rect 34244 40124 35420 40180
rect 35476 40124 35486 40180
rect 41570 40124 41580 40180
rect 41636 40124 42700 40180
rect 42756 40124 45388 40180
rect 45444 40124 45454 40180
rect 34188 40068 34244 40124
rect 49644 40068 49700 40236
rect 50418 40124 50428 40180
rect 50484 40124 50652 40180
rect 50708 40124 50718 40180
rect 17826 40012 17836 40068
rect 17892 40012 19292 40068
rect 19348 40012 19358 40068
rect 28914 40012 28924 40068
rect 28980 40012 29148 40068
rect 29204 40012 34244 40068
rect 40226 40012 40236 40068
rect 40292 40012 43260 40068
rect 43316 40012 43326 40068
rect 49644 40012 50988 40068
rect 51044 40012 51054 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 13682 39900 13692 39956
rect 13748 39900 26908 39956
rect 26964 39900 26974 39956
rect 39890 39900 39900 39956
rect 39956 39900 41468 39956
rect 41524 39900 41534 39956
rect 46274 39900 46284 39956
rect 46340 39900 50316 39956
rect 50372 39900 50382 39956
rect 15026 39788 15036 39844
rect 15092 39788 15372 39844
rect 15428 39788 15438 39844
rect 17714 39788 17724 39844
rect 17780 39788 18284 39844
rect 18340 39788 18350 39844
rect 20850 39788 20860 39844
rect 20916 39788 21868 39844
rect 21924 39788 25676 39844
rect 25732 39788 25742 39844
rect 28578 39788 28588 39844
rect 28644 39788 28924 39844
rect 28980 39788 31948 39844
rect 32004 39788 32014 39844
rect 38882 39788 38892 39844
rect 38948 39788 47292 39844
rect 47348 39788 47358 39844
rect 47842 39788 47852 39844
rect 47908 39788 49420 39844
rect 49476 39788 49644 39844
rect 49700 39788 49710 39844
rect 50194 39788 50204 39844
rect 50260 39788 50652 39844
rect 50708 39788 50718 39844
rect 11442 39676 11452 39732
rect 11508 39676 12236 39732
rect 12292 39676 12302 39732
rect 12674 39676 12684 39732
rect 12740 39676 21308 39732
rect 21364 39676 21374 39732
rect 23538 39676 23548 39732
rect 23604 39676 23642 39732
rect 36418 39676 36428 39732
rect 36484 39676 37100 39732
rect 37156 39676 37166 39732
rect 41906 39676 41916 39732
rect 41972 39676 42588 39732
rect 42644 39676 42654 39732
rect 49494 39676 49532 39732
rect 49588 39676 49598 39732
rect 15474 39564 15484 39620
rect 15540 39564 16492 39620
rect 16548 39564 16558 39620
rect 17276 39564 17780 39620
rect 18610 39564 18620 39620
rect 18676 39564 22428 39620
rect 22484 39564 22494 39620
rect 25330 39564 25340 39620
rect 25396 39564 26572 39620
rect 26628 39564 27916 39620
rect 27972 39564 28588 39620
rect 28644 39564 28654 39620
rect 39890 39564 39900 39620
rect 39956 39564 41244 39620
rect 41300 39564 41310 39620
rect 45378 39564 45388 39620
rect 45444 39564 46284 39620
rect 46340 39564 46350 39620
rect 47954 39564 47964 39620
rect 48020 39564 48972 39620
rect 49028 39564 49038 39620
rect 49298 39564 49308 39620
rect 49364 39564 49756 39620
rect 49812 39564 49822 39620
rect 13010 39452 13020 39508
rect 13076 39452 17052 39508
rect 17108 39452 17118 39508
rect 17276 39396 17332 39564
rect 17724 39508 17780 39564
rect 17490 39452 17500 39508
rect 17556 39452 17566 39508
rect 17724 39452 19628 39508
rect 19684 39452 19964 39508
rect 20020 39452 20030 39508
rect 20514 39452 20524 39508
rect 20580 39452 21084 39508
rect 21140 39452 21868 39508
rect 21924 39452 21934 39508
rect 26002 39452 26012 39508
rect 26068 39452 28252 39508
rect 28308 39452 28318 39508
rect 40674 39452 40684 39508
rect 40740 39452 44268 39508
rect 44324 39452 44828 39508
rect 44884 39452 44894 39508
rect 45602 39452 45612 39508
rect 45668 39452 45836 39508
rect 45892 39452 45902 39508
rect 46162 39452 46172 39508
rect 46228 39452 49084 39508
rect 49140 39452 49150 39508
rect 49606 39452 49644 39508
rect 49700 39452 49710 39508
rect 4274 39340 4284 39396
rect 4340 39340 5180 39396
rect 5236 39340 5246 39396
rect 6066 39340 6076 39396
rect 6132 39340 6860 39396
rect 6916 39340 6926 39396
rect 13906 39340 13916 39396
rect 13972 39340 14588 39396
rect 14644 39340 17332 39396
rect 17500 39396 17556 39452
rect 17500 39340 21420 39396
rect 21476 39340 22988 39396
rect 23044 39340 23054 39396
rect 29698 39340 29708 39396
rect 29764 39340 33740 39396
rect 33796 39340 33806 39396
rect 43698 39340 43708 39396
rect 43764 39340 44604 39396
rect 44660 39340 44670 39396
rect 45042 39340 45052 39396
rect 45108 39340 45276 39396
rect 45332 39340 45342 39396
rect 45490 39340 45500 39396
rect 45556 39340 45566 39396
rect 3378 39228 3388 39284
rect 3444 39228 4732 39284
rect 4788 39228 6972 39284
rect 7028 39228 7038 39284
rect 14690 39228 14700 39284
rect 14756 39228 15148 39284
rect 15204 39228 15372 39284
rect 15428 39228 15438 39284
rect 17500 39172 17556 39340
rect 45500 39284 45556 39340
rect 22530 39228 22540 39284
rect 22596 39228 23100 39284
rect 23156 39228 26908 39284
rect 33394 39228 33404 39284
rect 33460 39228 35980 39284
rect 36036 39228 36046 39284
rect 45500 39228 47852 39284
rect 47908 39228 47918 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 26852 39172 26908 39228
rect 15250 39116 15260 39172
rect 15316 39116 15708 39172
rect 15764 39116 15774 39172
rect 16482 39116 16492 39172
rect 16548 39116 17556 39172
rect 18610 39116 18620 39172
rect 18676 39116 19292 39172
rect 19348 39116 19358 39172
rect 26852 39116 37548 39172
rect 37604 39116 37614 39172
rect 6514 39004 6524 39060
rect 6580 39004 7532 39060
rect 7588 39004 7598 39060
rect 11890 39004 11900 39060
rect 11956 39004 16268 39060
rect 16324 39004 16334 39060
rect 17378 39004 17388 39060
rect 17444 39004 17724 39060
rect 17780 39004 17790 39060
rect 17938 39004 17948 39060
rect 18004 39004 18042 39060
rect 19730 39004 19740 39060
rect 19796 39004 20860 39060
rect 20916 39004 20926 39060
rect 26674 39004 26684 39060
rect 26740 39004 27692 39060
rect 27748 39004 29036 39060
rect 29092 39004 30156 39060
rect 30212 39004 30222 39060
rect 45500 38948 45556 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 47730 39004 47740 39060
rect 47796 39004 49644 39060
rect 49700 39004 50428 39060
rect 50484 39004 50494 39060
rect 4834 38892 4844 38948
rect 4900 38892 5292 38948
rect 5348 38892 5358 38948
rect 5506 38892 5516 38948
rect 5572 38892 6188 38948
rect 6244 38892 6254 38948
rect 13794 38892 13804 38948
rect 13860 38892 15372 38948
rect 15428 38892 15438 38948
rect 16034 38892 16044 38948
rect 16100 38892 20524 38948
rect 20580 38892 20590 38948
rect 42130 38892 42140 38948
rect 42196 38892 45948 38948
rect 46004 38892 46014 38948
rect 46946 38892 46956 38948
rect 47012 38892 47852 38948
rect 47908 38892 48748 38948
rect 48804 38892 48814 38948
rect 49522 38892 49532 38948
rect 49588 38892 49756 38948
rect 49812 38892 49822 38948
rect 6850 38780 6860 38836
rect 6916 38780 7420 38836
rect 7476 38780 8764 38836
rect 8820 38780 8830 38836
rect 14130 38780 14140 38836
rect 14196 38780 15148 38836
rect 15204 38780 15214 38836
rect 17490 38780 17500 38836
rect 17556 38780 20300 38836
rect 20356 38780 20366 38836
rect 20738 38780 20748 38836
rect 20804 38780 21756 38836
rect 21812 38780 21822 38836
rect 38210 38780 38220 38836
rect 38276 38780 38668 38836
rect 38724 38780 38734 38836
rect 41570 38780 41580 38836
rect 41636 38780 42028 38836
rect 42084 38780 42700 38836
rect 42756 38780 42766 38836
rect 44594 38780 44604 38836
rect 44660 38780 46620 38836
rect 46676 38780 46686 38836
rect 48290 38780 48300 38836
rect 48356 38780 50316 38836
rect 50372 38780 50382 38836
rect 16370 38668 16380 38724
rect 16436 38668 18284 38724
rect 18340 38668 18350 38724
rect 22978 38668 22988 38724
rect 23044 38668 30828 38724
rect 30884 38668 31948 38724
rect 32004 38668 32014 38724
rect 43362 38668 43372 38724
rect 43428 38668 43932 38724
rect 43988 38668 45724 38724
rect 45780 38668 45790 38724
rect 46386 38668 46396 38724
rect 46452 38668 46462 38724
rect 51650 38668 51660 38724
rect 51716 38668 53340 38724
rect 53396 38668 53406 38724
rect 46396 38612 46452 38668
rect 16454 38556 16492 38612
rect 16548 38556 16558 38612
rect 17154 38556 17164 38612
rect 17220 38556 17836 38612
rect 17892 38556 17902 38612
rect 18386 38556 18396 38612
rect 18452 38556 21756 38612
rect 21812 38556 21822 38612
rect 25442 38556 25452 38612
rect 25508 38556 26012 38612
rect 26068 38556 26078 38612
rect 44146 38556 44156 38612
rect 44212 38556 44828 38612
rect 44884 38556 48300 38612
rect 48356 38556 48366 38612
rect 17378 38444 17388 38500
rect 17444 38444 17948 38500
rect 18004 38444 18014 38500
rect 19954 38444 19964 38500
rect 20020 38444 23996 38500
rect 24052 38444 24668 38500
rect 24724 38444 24734 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 9650 38332 9660 38388
rect 9716 38332 12684 38388
rect 12740 38332 12750 38388
rect 15586 38332 15596 38388
rect 15652 38332 17276 38388
rect 17332 38332 17342 38388
rect 22978 38332 22988 38388
rect 23044 38332 27916 38388
rect 27972 38332 28476 38388
rect 28532 38332 28542 38388
rect 36754 38332 36764 38388
rect 36820 38332 37884 38388
rect 37940 38332 37950 38388
rect 38098 38332 38108 38388
rect 38164 38332 38444 38388
rect 38500 38332 38510 38388
rect 14690 38220 14700 38276
rect 14756 38220 16604 38276
rect 16660 38220 27020 38276
rect 27076 38220 27086 38276
rect 33282 38220 33292 38276
rect 33348 38220 34636 38276
rect 34692 38220 34702 38276
rect 38182 38220 38220 38276
rect 38276 38220 38286 38276
rect 4610 38108 4620 38164
rect 4676 38108 5516 38164
rect 5572 38108 5582 38164
rect 17602 38108 17612 38164
rect 17668 38108 18508 38164
rect 18564 38108 20748 38164
rect 20804 38108 20814 38164
rect 21746 38108 21756 38164
rect 21812 38108 22988 38164
rect 23044 38108 23054 38164
rect 38098 38108 38108 38164
rect 38164 38108 38668 38164
rect 45042 38108 45052 38164
rect 45108 38108 45836 38164
rect 45892 38108 45902 38164
rect 1810 37996 1820 38052
rect 1876 37996 5124 38052
rect 10098 37996 10108 38052
rect 10164 37996 15820 38052
rect 15876 37996 15886 38052
rect 28578 37996 28588 38052
rect 28644 37996 29484 38052
rect 29540 37996 30268 38052
rect 30324 37996 30334 38052
rect 37202 37996 37212 38052
rect 37268 37996 38220 38052
rect 38276 37996 38286 38052
rect 2482 37884 2492 37940
rect 2548 37884 3500 37940
rect 3556 37884 3566 37940
rect 5068 37828 5124 37996
rect 11778 37884 11788 37940
rect 11844 37884 14812 37940
rect 14868 37884 14878 37940
rect 23986 37884 23996 37940
rect 24052 37884 25900 37940
rect 25956 37884 25966 37940
rect 29810 37884 29820 37940
rect 29876 37884 30716 37940
rect 30772 37884 31164 37940
rect 31220 37884 31230 37940
rect 36530 37884 36540 37940
rect 36596 37884 37324 37940
rect 37380 37884 37390 37940
rect 5058 37772 5068 37828
rect 5124 37772 5964 37828
rect 6020 37772 8428 37828
rect 8484 37772 8876 37828
rect 8932 37772 9212 37828
rect 9268 37772 9278 37828
rect 17378 37772 17388 37828
rect 17444 37772 19628 37828
rect 19684 37772 19694 37828
rect 35074 37772 35084 37828
rect 35140 37772 36204 37828
rect 36260 37772 36270 37828
rect 16034 37660 16044 37716
rect 16100 37660 18732 37716
rect 18788 37660 18798 37716
rect 33954 37660 33964 37716
rect 34020 37660 34030 37716
rect 37090 37660 37100 37716
rect 37156 37660 37166 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 33964 37604 34020 37660
rect 37100 37604 37156 37660
rect 38612 37604 38668 38108
rect 51762 37996 51772 38052
rect 51828 37996 52780 38052
rect 52836 37996 52846 38052
rect 53554 37996 53564 38052
rect 53620 37996 54572 38052
rect 54628 37996 54638 38052
rect 53564 37940 53620 37996
rect 42802 37884 42812 37940
rect 42868 37884 43708 37940
rect 43764 37884 43774 37940
rect 45126 37884 45164 37940
rect 45220 37884 45230 37940
rect 45378 37884 45388 37940
rect 45444 37884 45612 37940
rect 45668 37884 45678 37940
rect 45826 37884 45836 37940
rect 45892 37884 46396 37940
rect 46452 37884 48188 37940
rect 48244 37884 48254 37940
rect 50978 37884 50988 37940
rect 51044 37884 52556 37940
rect 52612 37884 53620 37940
rect 44482 37772 44492 37828
rect 44548 37772 44828 37828
rect 44884 37772 44894 37828
rect 50306 37772 50316 37828
rect 50372 37772 51100 37828
rect 51156 37772 51166 37828
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 33964 37548 34412 37604
rect 34468 37548 35868 37604
rect 35924 37548 36428 37604
rect 36484 37548 37156 37604
rect 38182 37548 38220 37604
rect 38276 37548 38286 37604
rect 38612 37548 39788 37604
rect 39844 37548 39854 37604
rect 3714 37436 3724 37492
rect 3780 37436 4620 37492
rect 4676 37436 5180 37492
rect 5236 37436 5246 37492
rect 14018 37436 14028 37492
rect 14084 37436 14364 37492
rect 14420 37436 14430 37492
rect 20066 37436 20076 37492
rect 20132 37436 21476 37492
rect 22978 37436 22988 37492
rect 23044 37436 24108 37492
rect 24164 37436 24174 37492
rect 31490 37436 31500 37492
rect 31556 37436 38892 37492
rect 38948 37436 38958 37492
rect 43474 37436 43484 37492
rect 43540 37436 43550 37492
rect 43810 37436 43820 37492
rect 43876 37436 45724 37492
rect 45780 37436 45790 37492
rect 21420 37380 21476 37436
rect 43484 37380 43540 37436
rect 15026 37324 15036 37380
rect 15092 37324 15372 37380
rect 15428 37324 15438 37380
rect 17826 37324 17836 37380
rect 17892 37324 20300 37380
rect 20356 37324 20366 37380
rect 21410 37324 21420 37380
rect 21476 37324 22484 37380
rect 36194 37324 36204 37380
rect 36260 37324 36876 37380
rect 36932 37324 37212 37380
rect 37268 37324 37278 37380
rect 37650 37324 37660 37380
rect 37716 37324 37996 37380
rect 38052 37324 38062 37380
rect 43484 37324 43764 37380
rect 43922 37324 43932 37380
rect 43988 37324 44380 37380
rect 44436 37324 46676 37380
rect 22428 37268 22484 37324
rect 3378 37212 3388 37268
rect 3444 37212 3836 37268
rect 3892 37212 4284 37268
rect 4340 37212 6524 37268
rect 6580 37212 6590 37268
rect 11106 37212 11116 37268
rect 11172 37212 12572 37268
rect 12628 37212 12638 37268
rect 13682 37212 13692 37268
rect 13748 37212 14364 37268
rect 14420 37212 18732 37268
rect 18788 37212 18798 37268
rect 19058 37212 19068 37268
rect 19124 37212 21308 37268
rect 21364 37212 21644 37268
rect 21700 37212 21710 37268
rect 22418 37212 22428 37268
rect 22484 37212 25564 37268
rect 25620 37212 25630 37268
rect 27234 37212 27244 37268
rect 27300 37212 30492 37268
rect 30548 37212 31724 37268
rect 31780 37212 33068 37268
rect 33124 37212 35084 37268
rect 35140 37212 35150 37268
rect 35308 37212 43540 37268
rect 35308 37156 35364 37212
rect 15698 37100 15708 37156
rect 15764 37100 18396 37156
rect 18452 37100 18462 37156
rect 19590 37100 19628 37156
rect 19684 37100 19694 37156
rect 19842 37100 19852 37156
rect 19908 37100 20636 37156
rect 20692 37100 20702 37156
rect 30034 37100 30044 37156
rect 30100 37100 30940 37156
rect 30996 37100 31006 37156
rect 32050 37100 32060 37156
rect 32116 37100 35364 37156
rect 15026 36988 15036 37044
rect 15092 36988 15652 37044
rect 15810 36988 15820 37044
rect 15876 36988 17836 37044
rect 17892 36988 17902 37044
rect 18722 36988 18732 37044
rect 18788 36988 19404 37044
rect 19460 36988 19470 37044
rect 15596 36932 15652 36988
rect 19852 36932 19908 37100
rect 32060 37044 32116 37100
rect 38612 37044 38668 37156
rect 38724 37100 38734 37156
rect 40898 37100 40908 37156
rect 40964 37100 41692 37156
rect 41748 37100 42476 37156
rect 42532 37100 42542 37156
rect 43484 37044 43540 37212
rect 43708 37044 43764 37324
rect 46620 37268 46676 37324
rect 45798 37212 45836 37268
rect 45892 37212 45902 37268
rect 46610 37212 46620 37268
rect 46676 37212 50316 37268
rect 50372 37212 50382 37268
rect 51090 37212 51100 37268
rect 51156 37212 54124 37268
rect 54180 37212 54190 37268
rect 45266 37100 45276 37156
rect 45332 37100 47404 37156
rect 47460 37100 47470 37156
rect 20178 36988 20188 37044
rect 20244 36988 23324 37044
rect 23380 36988 24556 37044
rect 24612 36988 25284 37044
rect 26898 36988 26908 37044
rect 26964 36988 32116 37044
rect 34626 36988 34636 37044
rect 34692 36988 38668 37044
rect 43474 36988 43484 37044
rect 43540 36988 43550 37044
rect 43708 36988 45500 37044
rect 45556 36988 46060 37044
rect 46116 36988 46844 37044
rect 46900 36988 46910 37044
rect 53554 36988 53564 37044
rect 53620 36988 54796 37044
rect 54852 36988 54862 37044
rect 15596 36876 15932 36932
rect 15988 36876 15998 36932
rect 19282 36876 19292 36932
rect 19348 36876 19908 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 25228 36820 25284 36988
rect 28018 36876 28028 36932
rect 28084 36876 33404 36932
rect 33460 36876 33470 36932
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 37324 36820 37380 36988
rect 43708 36932 43764 36988
rect 43362 36876 43372 36932
rect 43428 36876 43764 36932
rect 43922 36876 43932 36932
rect 43988 36876 45276 36932
rect 45332 36876 46172 36932
rect 46228 36876 46238 36932
rect 48850 36876 48860 36932
rect 48916 36876 50428 36932
rect 50484 36876 52556 36932
rect 52612 36876 54684 36932
rect 54740 36876 54750 36932
rect 19170 36764 19180 36820
rect 19236 36764 20636 36820
rect 20692 36764 20702 36820
rect 25218 36764 25228 36820
rect 25284 36764 25294 36820
rect 37314 36764 37324 36820
rect 37380 36764 37390 36820
rect 46386 36764 46396 36820
rect 46452 36764 51660 36820
rect 51716 36764 52332 36820
rect 52388 36764 52398 36820
rect 55458 36764 55468 36820
rect 55524 36764 56364 36820
rect 56420 36764 56430 36820
rect 13794 36652 13804 36708
rect 13860 36652 15820 36708
rect 15876 36652 16156 36708
rect 16212 36652 16222 36708
rect 36530 36652 36540 36708
rect 36596 36652 37212 36708
rect 37268 36652 42476 36708
rect 42532 36652 44156 36708
rect 44212 36652 44222 36708
rect 46274 36652 46284 36708
rect 46340 36652 49868 36708
rect 49924 36652 52892 36708
rect 52948 36652 52958 36708
rect 54562 36652 54572 36708
rect 54628 36652 55468 36708
rect 55412 36596 55468 36652
rect 15092 36540 16716 36596
rect 16772 36540 16782 36596
rect 19180 36540 27356 36596
rect 27412 36540 28140 36596
rect 28196 36540 28588 36596
rect 28644 36540 29484 36596
rect 29540 36540 29550 36596
rect 30034 36540 30044 36596
rect 30100 36540 34300 36596
rect 34356 36540 34366 36596
rect 39442 36540 39452 36596
rect 39508 36540 40348 36596
rect 40404 36540 40414 36596
rect 47618 36540 47628 36596
rect 47684 36540 48972 36596
rect 49028 36540 49038 36596
rect 50194 36540 50204 36596
rect 50260 36540 55020 36596
rect 55076 36540 55086 36596
rect 55402 36540 55412 36596
rect 55468 36540 55478 36596
rect 15092 36484 15148 36540
rect 19180 36484 19236 36540
rect 55580 36484 55636 36764
rect 14018 36428 14028 36484
rect 14084 36428 15148 36484
rect 15250 36428 15260 36484
rect 15316 36428 19236 36484
rect 20514 36428 20524 36484
rect 20580 36428 21756 36484
rect 21812 36428 22204 36484
rect 22260 36428 22270 36484
rect 32498 36428 32508 36484
rect 32564 36428 33516 36484
rect 33572 36428 33964 36484
rect 34020 36428 34030 36484
rect 36082 36428 36092 36484
rect 36148 36428 36988 36484
rect 37044 36428 37054 36484
rect 38612 36428 39676 36484
rect 39732 36428 39742 36484
rect 43474 36428 43484 36484
rect 43540 36428 45276 36484
rect 45332 36428 45342 36484
rect 47170 36428 47180 36484
rect 47236 36428 48748 36484
rect 48804 36428 48814 36484
rect 54002 36428 54012 36484
rect 54068 36428 54572 36484
rect 54628 36428 55636 36484
rect 38612 36372 38668 36428
rect 13794 36316 13804 36372
rect 13860 36316 15932 36372
rect 15988 36316 15998 36372
rect 16482 36316 16492 36372
rect 16548 36316 22428 36372
rect 22484 36316 25900 36372
rect 25956 36316 25966 36372
rect 27682 36316 27692 36372
rect 27748 36316 38668 36372
rect 47058 36316 47068 36372
rect 47124 36316 47516 36372
rect 47572 36316 52668 36372
rect 52724 36316 52734 36372
rect 54114 36316 54124 36372
rect 54180 36316 54460 36372
rect 54516 36316 55580 36372
rect 55636 36316 56028 36372
rect 56084 36316 56094 36372
rect 18946 36204 18956 36260
rect 19012 36204 19516 36260
rect 19572 36204 19582 36260
rect 31826 36204 31836 36260
rect 31892 36204 32396 36260
rect 32452 36204 32462 36260
rect 44930 36204 44940 36260
rect 44996 36204 45500 36260
rect 45556 36204 47740 36260
rect 47796 36204 47806 36260
rect 52098 36204 52108 36260
rect 52164 36204 52174 36260
rect 54226 36204 54236 36260
rect 54292 36204 57260 36260
rect 57316 36204 57820 36260
rect 57876 36204 57886 36260
rect 52108 36148 52164 36204
rect 20290 36092 20300 36148
rect 20356 36092 21308 36148
rect 21364 36092 21374 36148
rect 35746 36092 35756 36148
rect 35812 36092 40684 36148
rect 40740 36092 40750 36148
rect 42802 36092 42812 36148
rect 42868 36092 45164 36148
rect 45220 36092 45230 36148
rect 48066 36092 48076 36148
rect 48132 36092 50204 36148
rect 50260 36092 50270 36148
rect 52108 36092 55580 36148
rect 55636 36092 55646 36148
rect 56130 36092 56140 36148
rect 56196 36092 57036 36148
rect 57092 36092 57102 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 19478 35980 19516 36036
rect 19572 35980 19582 36036
rect 22194 35980 22204 36036
rect 22260 35980 22876 36036
rect 22932 35980 23212 36036
rect 23268 35980 23278 36036
rect 28812 35980 30828 36036
rect 30884 35980 32172 36036
rect 32228 35980 32238 36036
rect 54674 35980 54684 36036
rect 54740 35980 57372 36036
rect 57428 35980 57438 36036
rect 28812 35924 28868 35980
rect 15810 35868 15820 35924
rect 15876 35868 17388 35924
rect 17444 35868 17948 35924
rect 18004 35868 18014 35924
rect 18610 35868 18620 35924
rect 18676 35868 20188 35924
rect 20244 35868 20254 35924
rect 20738 35868 20748 35924
rect 20804 35868 22988 35924
rect 23044 35868 23436 35924
rect 23492 35868 23502 35924
rect 24882 35868 24892 35924
rect 24948 35868 25564 35924
rect 25620 35868 28812 35924
rect 28868 35868 28878 35924
rect 29250 35868 29260 35924
rect 29316 35868 30268 35924
rect 30324 35868 30334 35924
rect 45154 35868 45164 35924
rect 45220 35868 45948 35924
rect 46004 35868 47068 35924
rect 47124 35868 47134 35924
rect 50754 35868 50764 35924
rect 50820 35868 51212 35924
rect 51268 35868 52892 35924
rect 52948 35868 52958 35924
rect 55122 35868 55132 35924
rect 55188 35868 56700 35924
rect 56756 35868 56766 35924
rect 15922 35756 15932 35812
rect 15988 35756 19068 35812
rect 19124 35756 24444 35812
rect 24500 35756 24510 35812
rect 30482 35756 30492 35812
rect 30548 35756 33740 35812
rect 33796 35756 33806 35812
rect 36642 35756 36652 35812
rect 36708 35756 38332 35812
rect 38388 35756 38398 35812
rect 16034 35644 16044 35700
rect 16100 35644 16716 35700
rect 16772 35644 16782 35700
rect 23314 35644 23324 35700
rect 23380 35644 23884 35700
rect 23940 35644 26124 35700
rect 26180 35644 26190 35700
rect 37538 35644 37548 35700
rect 37604 35644 38780 35700
rect 38836 35644 38846 35700
rect 44258 35644 44268 35700
rect 44324 35644 44716 35700
rect 44772 35644 45164 35700
rect 45220 35644 45724 35700
rect 45780 35644 47852 35700
rect 47908 35644 47918 35700
rect 49410 35644 49420 35700
rect 49476 35644 49486 35700
rect 49970 35644 49980 35700
rect 50036 35644 50764 35700
rect 50820 35644 50830 35700
rect 54786 35644 54796 35700
rect 54852 35644 55356 35700
rect 55412 35644 55422 35700
rect 23324 35476 23380 35644
rect 26002 35532 26012 35588
rect 26068 35532 27916 35588
rect 27972 35532 27982 35588
rect 49420 35476 49476 35644
rect 55794 35532 55804 35588
rect 55860 35532 56700 35588
rect 56756 35532 56766 35588
rect 16594 35420 16604 35476
rect 16660 35420 18620 35476
rect 18676 35420 22428 35476
rect 22484 35420 23380 35476
rect 34290 35420 34300 35476
rect 34356 35420 40236 35476
rect 40292 35420 40302 35476
rect 47282 35420 47292 35476
rect 47348 35420 48748 35476
rect 48804 35420 49476 35476
rect 55906 35420 55916 35476
rect 55972 35420 57708 35476
rect 57764 35420 57774 35476
rect 13234 35308 13244 35364
rect 13300 35308 13310 35364
rect 14018 35308 14028 35364
rect 14084 35308 17276 35364
rect 17332 35308 20748 35364
rect 20804 35308 20814 35364
rect 33842 35308 33852 35364
rect 33908 35308 34972 35364
rect 35028 35308 35038 35364
rect 47058 35308 47068 35364
rect 47124 35308 47516 35364
rect 47572 35308 47582 35364
rect 51538 35308 51548 35364
rect 51604 35308 55132 35364
rect 55188 35308 55198 35364
rect 57138 35308 57148 35364
rect 57204 35308 57820 35364
rect 57876 35308 57886 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 13244 35252 13300 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 13244 35196 15036 35252
rect 15092 35196 15102 35252
rect 17154 35196 17164 35252
rect 17220 35196 19628 35252
rect 19684 35196 19694 35252
rect 22754 35196 22764 35252
rect 22820 35196 25228 35252
rect 25284 35196 25294 35252
rect 38770 35196 38780 35252
rect 38836 35196 41020 35252
rect 41076 35196 42140 35252
rect 42196 35196 42206 35252
rect 43698 35196 43708 35252
rect 43764 35196 44380 35252
rect 44436 35196 45276 35252
rect 45332 35196 45342 35252
rect 48962 35196 48972 35252
rect 49028 35196 52892 35252
rect 52948 35196 52958 35252
rect 53330 35196 53340 35252
rect 53396 35196 53676 35252
rect 53732 35196 53742 35252
rect 12674 35084 12684 35140
rect 12740 35084 13580 35140
rect 13636 35084 13646 35140
rect 18498 35084 18508 35140
rect 18564 35084 18956 35140
rect 19012 35084 19022 35140
rect 23762 35084 23772 35140
rect 23828 35084 24556 35140
rect 24612 35084 24622 35140
rect 31266 35084 31276 35140
rect 31332 35084 52668 35140
rect 52724 35084 55580 35140
rect 55636 35084 57036 35140
rect 57092 35084 57102 35140
rect 15362 34972 15372 35028
rect 15428 34972 18732 35028
rect 18788 34972 18798 35028
rect 29250 34972 29260 35028
rect 29316 34972 34860 35028
rect 34916 34972 36428 35028
rect 36484 34972 37884 35028
rect 37940 34972 37950 35028
rect 10546 34860 10556 34916
rect 10612 34860 18844 34916
rect 18900 34860 21308 34916
rect 21364 34860 21374 34916
rect 29138 34860 29148 34916
rect 29204 34860 29484 34916
rect 29540 34860 30268 34916
rect 30324 34860 30334 34916
rect 49298 34860 49308 34916
rect 49364 34860 50428 34916
rect 50484 34860 51772 34916
rect 51828 34860 51838 34916
rect 52322 34860 52332 34916
rect 52388 34860 53508 34916
rect 54450 34860 54460 34916
rect 54516 34860 55356 34916
rect 55412 34860 56812 34916
rect 56868 34860 57260 34916
rect 57316 34860 57326 34916
rect 53452 34804 53508 34860
rect 20738 34748 20748 34804
rect 20804 34748 21980 34804
rect 22036 34748 22046 34804
rect 27010 34748 27020 34804
rect 27076 34748 33180 34804
rect 33236 34748 35756 34804
rect 35812 34748 35822 34804
rect 45714 34748 45724 34804
rect 45780 34748 46396 34804
rect 46452 34748 47628 34804
rect 47684 34748 47694 34804
rect 48738 34748 48748 34804
rect 48804 34748 49420 34804
rect 49476 34748 49486 34804
rect 50082 34748 50092 34804
rect 50148 34748 51100 34804
rect 51156 34748 53228 34804
rect 53284 34748 53294 34804
rect 53442 34748 53452 34804
rect 53508 34748 56588 34804
rect 56644 34748 56654 34804
rect 27122 34636 27132 34692
rect 27188 34636 29372 34692
rect 29428 34636 29438 34692
rect 34066 34636 34076 34692
rect 34132 34636 34300 34692
rect 34356 34636 34366 34692
rect 43922 34636 43932 34692
rect 43988 34636 48972 34692
rect 49028 34636 49038 34692
rect 54674 34636 54684 34692
rect 54740 34636 56812 34692
rect 56868 34636 57708 34692
rect 57764 34636 57774 34692
rect 49074 34524 49084 34580
rect 49140 34524 49756 34580
rect 49812 34524 49822 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 24658 34300 24668 34356
rect 24724 34300 25452 34356
rect 25508 34300 27468 34356
rect 27524 34300 27534 34356
rect 48514 34300 48524 34356
rect 48580 34300 50428 34356
rect 51650 34300 51660 34356
rect 51716 34300 53676 34356
rect 53732 34300 55468 34356
rect 50372 34244 50428 34300
rect 18946 34188 18956 34244
rect 19012 34188 23772 34244
rect 23828 34188 23838 34244
rect 36530 34188 36540 34244
rect 36596 34188 38108 34244
rect 38164 34188 39956 34244
rect 43810 34188 43820 34244
rect 43876 34188 45164 34244
rect 45220 34188 45230 34244
rect 48178 34188 48188 34244
rect 48244 34188 49644 34244
rect 49700 34188 50204 34244
rect 50260 34188 50270 34244
rect 50372 34188 50652 34244
rect 50708 34188 50718 34244
rect 39900 34132 39956 34188
rect 55412 34132 55468 34300
rect 56018 34188 56028 34244
rect 56084 34188 57148 34244
rect 57204 34188 57214 34244
rect 17714 34076 17724 34132
rect 17780 34076 18620 34132
rect 18676 34076 18686 34132
rect 19058 34076 19068 34132
rect 19124 34076 20860 34132
rect 20916 34076 25340 34132
rect 25396 34076 25406 34132
rect 26450 34076 26460 34132
rect 26516 34076 29596 34132
rect 29652 34076 29662 34132
rect 33506 34076 33516 34132
rect 33572 34076 33964 34132
rect 34020 34076 34030 34132
rect 34178 34076 34188 34132
rect 34244 34076 34692 34132
rect 38770 34076 38780 34132
rect 38836 34076 38846 34132
rect 39890 34076 39900 34132
rect 39956 34076 40908 34132
rect 40964 34076 40974 34132
rect 42018 34076 42028 34132
rect 42084 34076 42094 34132
rect 42578 34076 42588 34132
rect 42644 34076 48748 34132
rect 48804 34076 50428 34132
rect 50484 34076 50494 34132
rect 51090 34076 51100 34132
rect 51156 34076 54124 34132
rect 54180 34076 54190 34132
rect 55412 34076 56812 34132
rect 56868 34076 56878 34132
rect 17938 33964 17948 34020
rect 18004 33964 20412 34020
rect 20468 33964 21308 34020
rect 21364 33964 33628 34020
rect 33684 33964 34412 34020
rect 34468 33964 34478 34020
rect 34636 33908 34692 34076
rect 38780 34020 38836 34076
rect 36428 33964 38836 34020
rect 36428 33908 36484 33964
rect 42028 33908 42084 34076
rect 54124 34020 54180 34076
rect 49410 33964 49420 34020
rect 49476 33964 51660 34020
rect 51716 33964 51726 34020
rect 54124 33964 56476 34020
rect 56532 33964 56542 34020
rect 14802 33852 14812 33908
rect 14868 33852 17612 33908
rect 17668 33852 24332 33908
rect 24388 33852 24398 33908
rect 26002 33852 26012 33908
rect 26068 33852 27132 33908
rect 27188 33852 27198 33908
rect 32498 33852 32508 33908
rect 32564 33852 34748 33908
rect 34804 33852 34814 33908
rect 35074 33852 35084 33908
rect 35140 33852 36036 33908
rect 36418 33852 36428 33908
rect 36484 33852 36494 33908
rect 38612 33852 42084 33908
rect 50194 33852 50204 33908
rect 50260 33852 51212 33908
rect 51268 33852 51278 33908
rect 35980 33796 36036 33852
rect 38612 33796 38668 33852
rect 14130 33740 14140 33796
rect 14196 33740 18956 33796
rect 19012 33740 19022 33796
rect 19282 33740 19292 33796
rect 19348 33740 20412 33796
rect 20468 33740 20478 33796
rect 35970 33740 35980 33796
rect 36036 33740 38668 33796
rect 43586 33740 43596 33796
rect 43652 33740 44716 33796
rect 44772 33740 45500 33796
rect 45556 33740 45566 33796
rect 50978 33740 50988 33796
rect 51044 33740 54236 33796
rect 54292 33740 54302 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 18722 33628 18732 33684
rect 18788 33628 19404 33684
rect 19460 33628 19470 33684
rect 20514 33628 20524 33684
rect 20580 33628 21756 33684
rect 21812 33628 21822 33684
rect 34290 33628 34300 33684
rect 34356 33628 34972 33684
rect 35028 33628 35038 33684
rect 41682 33628 41692 33684
rect 41748 33628 47068 33684
rect 47124 33628 47134 33684
rect 51202 33628 51212 33684
rect 51268 33628 53900 33684
rect 53956 33628 53966 33684
rect 43922 33516 43932 33572
rect 43988 33516 45836 33572
rect 45892 33516 45902 33572
rect 30370 33404 30380 33460
rect 30436 33404 32732 33460
rect 32788 33404 33180 33460
rect 33236 33404 33246 33460
rect 36204 33292 36988 33348
rect 37044 33292 37054 33348
rect 46498 33292 46508 33348
rect 46564 33292 47180 33348
rect 47236 33292 47246 33348
rect 50866 33292 50876 33348
rect 50932 33292 54236 33348
rect 54292 33292 57932 33348
rect 57988 33292 57998 33348
rect 36204 33236 36260 33292
rect 15810 33180 15820 33236
rect 15876 33180 16380 33236
rect 16436 33180 16828 33236
rect 16884 33180 18340 33236
rect 23426 33180 23436 33236
rect 23492 33180 30044 33236
rect 30100 33180 30110 33236
rect 35410 33180 35420 33236
rect 35476 33180 36204 33236
rect 36260 33180 36270 33236
rect 36428 33180 37212 33236
rect 37268 33180 37278 33236
rect 52098 33180 52108 33236
rect 52164 33180 53564 33236
rect 53620 33180 53630 33236
rect 18284 33124 18340 33180
rect 36428 33124 36484 33180
rect 11778 33068 11788 33124
rect 11844 33068 17948 33124
rect 18004 33068 18014 33124
rect 18274 33068 18284 33124
rect 18340 33068 19740 33124
rect 19796 33068 20244 33124
rect 20514 33068 20524 33124
rect 20580 33068 24892 33124
rect 24948 33068 24958 33124
rect 36418 33068 36428 33124
rect 36484 33068 36494 33124
rect 37090 33068 37100 33124
rect 37156 33068 39676 33124
rect 39732 33068 40348 33124
rect 40404 33068 40414 33124
rect 47170 33068 47180 33124
rect 47236 33068 49196 33124
rect 49252 33068 49262 33124
rect 20188 33012 20244 33068
rect 20188 32956 21420 33012
rect 21476 32956 21868 33012
rect 21924 32956 22428 33012
rect 22484 32956 23324 33012
rect 23380 32956 23660 33012
rect 23716 32956 24444 33012
rect 24500 32956 24510 33012
rect 45378 32956 45388 33012
rect 45444 32956 46844 33012
rect 46900 32956 46910 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 47954 32844 47964 32900
rect 48020 32844 49084 32900
rect 49140 32844 49150 32900
rect 9426 32732 9436 32788
rect 9492 32732 29708 32788
rect 29764 32732 29774 32788
rect 36418 32732 36428 32788
rect 36484 32732 37100 32788
rect 37156 32732 37166 32788
rect 39116 32732 43372 32788
rect 43428 32732 43820 32788
rect 43876 32732 43886 32788
rect 46386 32732 46396 32788
rect 46452 32732 47516 32788
rect 47572 32732 47582 32788
rect 49186 32732 49196 32788
rect 49252 32732 52220 32788
rect 52276 32732 52286 32788
rect 39116 32676 39172 32732
rect 13346 32620 13356 32676
rect 13412 32620 32396 32676
rect 32452 32620 33292 32676
rect 33348 32620 33358 32676
rect 39106 32620 39116 32676
rect 39172 32620 39182 32676
rect 46918 32620 46956 32676
rect 47012 32620 47022 32676
rect 51650 32620 51660 32676
rect 51716 32620 54796 32676
rect 54852 32620 55244 32676
rect 55300 32620 55310 32676
rect 12450 32508 12460 32564
rect 12516 32508 13580 32564
rect 13636 32508 15708 32564
rect 15764 32508 15774 32564
rect 22306 32508 22316 32564
rect 22372 32508 23660 32564
rect 23716 32508 23726 32564
rect 42914 32508 42924 32564
rect 42980 32508 43708 32564
rect 43764 32508 43774 32564
rect 47730 32508 47740 32564
rect 47796 32508 49532 32564
rect 49588 32508 49756 32564
rect 49812 32508 50204 32564
rect 50260 32508 50764 32564
rect 50820 32508 50830 32564
rect 51762 32508 51772 32564
rect 51828 32508 54012 32564
rect 54068 32508 54078 32564
rect 27234 32396 27244 32452
rect 27300 32396 29148 32452
rect 29204 32396 29214 32452
rect 42802 32396 42812 32452
rect 42868 32396 43820 32452
rect 43876 32396 43886 32452
rect 33506 32284 33516 32340
rect 33572 32284 36652 32340
rect 36708 32284 36718 32340
rect 44818 32284 44828 32340
rect 44884 32284 46284 32340
rect 46340 32284 46350 32340
rect 49746 32284 49756 32340
rect 49812 32284 50316 32340
rect 50372 32284 50382 32340
rect 41458 32172 41468 32228
rect 41524 32172 50988 32228
rect 51044 32172 51054 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 46694 32060 46732 32116
rect 46788 32060 46798 32116
rect 15372 31948 15876 32004
rect 29586 31948 29596 32004
rect 29652 31948 30044 32004
rect 30100 31948 30110 32004
rect 35522 31948 35532 32004
rect 35588 31948 39956 32004
rect 15372 31892 15428 31948
rect 15820 31892 15876 31948
rect 39900 31892 39956 31948
rect 50988 31892 51044 32172
rect 51314 31948 51324 32004
rect 51380 31948 51996 32004
rect 52052 31948 52062 32004
rect 13122 31836 13132 31892
rect 13188 31836 13916 31892
rect 13972 31836 13982 31892
rect 14802 31836 14812 31892
rect 14868 31836 15428 31892
rect 15586 31836 15596 31892
rect 15652 31836 15662 31892
rect 15820 31836 21868 31892
rect 21924 31836 21934 31892
rect 26674 31836 26684 31892
rect 26740 31836 27356 31892
rect 27412 31836 31052 31892
rect 31108 31836 31118 31892
rect 33058 31836 33068 31892
rect 33124 31836 36204 31892
rect 36260 31836 36270 31892
rect 37314 31836 37324 31892
rect 37380 31836 38668 31892
rect 38724 31836 38734 31892
rect 39890 31836 39900 31892
rect 39956 31836 39966 31892
rect 40338 31836 40348 31892
rect 40404 31836 41468 31892
rect 41524 31836 41916 31892
rect 41972 31836 44940 31892
rect 44996 31836 46284 31892
rect 46340 31836 50316 31892
rect 50372 31836 50382 31892
rect 50988 31836 51660 31892
rect 51716 31836 51726 31892
rect 15596 31780 15652 31836
rect 13794 31724 13804 31780
rect 13860 31724 15652 31780
rect 15922 31724 15932 31780
rect 15988 31724 17836 31780
rect 17892 31724 17902 31780
rect 18386 31724 18396 31780
rect 18452 31724 20524 31780
rect 20580 31724 22540 31780
rect 22596 31724 22606 31780
rect 28242 31724 28252 31780
rect 28308 31724 32508 31780
rect 32564 31724 35644 31780
rect 35700 31724 37548 31780
rect 37604 31724 37614 31780
rect 40114 31724 40124 31780
rect 40180 31724 41804 31780
rect 41860 31724 44044 31780
rect 44100 31724 44110 31780
rect 44258 31724 44268 31780
rect 44324 31724 52668 31780
rect 52724 31724 53452 31780
rect 53508 31724 53518 31780
rect 13458 31612 13468 31668
rect 13524 31612 18732 31668
rect 18788 31612 20412 31668
rect 20468 31612 20478 31668
rect 20738 31612 20748 31668
rect 20804 31612 21980 31668
rect 22036 31612 22046 31668
rect 24994 31612 25004 31668
rect 25060 31612 26012 31668
rect 26068 31612 26078 31668
rect 34290 31612 34300 31668
rect 34356 31612 36988 31668
rect 37044 31612 37054 31668
rect 38210 31612 38220 31668
rect 38276 31612 39228 31668
rect 39284 31612 39294 31668
rect 43922 31612 43932 31668
rect 43988 31612 48188 31668
rect 48244 31612 48254 31668
rect 48402 31612 48412 31668
rect 48468 31612 51884 31668
rect 51940 31612 51950 31668
rect 15586 31500 15596 31556
rect 15652 31500 16492 31556
rect 16548 31500 20076 31556
rect 20132 31500 21308 31556
rect 21364 31500 21374 31556
rect 25666 31500 25676 31556
rect 25732 31500 26124 31556
rect 26180 31500 26190 31556
rect 33730 31500 33740 31556
rect 33796 31500 34524 31556
rect 34580 31500 39116 31556
rect 39172 31500 39182 31556
rect 39666 31500 39676 31556
rect 39732 31500 40348 31556
rect 40404 31500 40908 31556
rect 40964 31500 41804 31556
rect 41860 31500 41870 31556
rect 47618 31500 47628 31556
rect 47684 31500 49084 31556
rect 49140 31500 49150 31556
rect 51426 31500 51436 31556
rect 51492 31500 56700 31556
rect 56756 31500 56766 31556
rect 15922 31388 15932 31444
rect 15988 31388 17724 31444
rect 17780 31388 18396 31444
rect 18452 31388 18462 31444
rect 46806 31388 46844 31444
rect 46900 31388 46910 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 43250 31276 43260 31332
rect 43316 31276 43484 31332
rect 43540 31276 45388 31332
rect 45444 31276 48860 31332
rect 48916 31276 49756 31332
rect 49812 31276 49822 31332
rect 52546 31276 52556 31332
rect 52612 31276 53788 31332
rect 53844 31276 54348 31332
rect 54404 31276 54414 31332
rect 13234 31164 13244 31220
rect 13300 31164 14140 31220
rect 14196 31164 14588 31220
rect 14644 31164 14654 31220
rect 17826 31164 17836 31220
rect 17892 31164 18732 31220
rect 18788 31164 18798 31220
rect 24658 31164 24668 31220
rect 24724 31164 28028 31220
rect 28084 31164 28094 31220
rect 29698 31164 29708 31220
rect 29764 31164 31052 31220
rect 31108 31164 31118 31220
rect 44930 31164 44940 31220
rect 44996 31164 45500 31220
rect 45556 31164 49420 31220
rect 49476 31164 49486 31220
rect 51884 31164 52780 31220
rect 52836 31164 52846 31220
rect 51884 31108 51940 31164
rect 39890 31052 39900 31108
rect 39956 31052 41580 31108
rect 41636 31052 44156 31108
rect 44212 31052 44222 31108
rect 48178 31052 48188 31108
rect 48244 31052 51884 31108
rect 51940 31052 51950 31108
rect 52098 31052 52108 31108
rect 52164 31052 53788 31108
rect 53844 31052 54572 31108
rect 54628 31052 54638 31108
rect 29250 30940 29260 30996
rect 29316 30940 29708 30996
rect 29764 30940 29774 30996
rect 44706 30940 44716 30996
rect 44772 30940 45276 30996
rect 45332 30940 45342 30996
rect 46498 30940 46508 30996
rect 46564 30940 47180 30996
rect 47236 30940 47246 30996
rect 50306 30940 50316 30996
rect 50372 30940 54908 30996
rect 54964 30940 55356 30996
rect 55412 30940 57372 30996
rect 57428 30940 58044 30996
rect 58100 30940 58110 30996
rect 16370 30828 16380 30884
rect 16436 30828 17388 30884
rect 17444 30828 17948 30884
rect 18004 30828 18014 30884
rect 18274 30828 18284 30884
rect 18340 30828 19068 30884
rect 19124 30828 21308 30884
rect 21364 30828 21374 30884
rect 26674 30828 26684 30884
rect 26740 30828 27356 30884
rect 27412 30828 27422 30884
rect 46694 30828 46732 30884
rect 46788 30828 46798 30884
rect 49410 30828 49420 30884
rect 49476 30828 50204 30884
rect 50260 30828 52780 30884
rect 52836 30828 52846 30884
rect 55356 30828 55468 30940
rect 16146 30716 16156 30772
rect 16212 30716 16492 30772
rect 16548 30716 18732 30772
rect 18788 30716 18798 30772
rect 29474 30716 29484 30772
rect 29540 30716 30156 30772
rect 30212 30716 30222 30772
rect 32162 30716 32172 30772
rect 32228 30716 38668 30772
rect 40226 30716 40236 30772
rect 40292 30716 41020 30772
rect 41076 30716 41692 30772
rect 41748 30716 42588 30772
rect 42644 30716 42654 30772
rect 45042 30716 45052 30772
rect 45108 30716 45612 30772
rect 45668 30716 45678 30772
rect 38612 30660 38668 30716
rect 38612 30604 40572 30660
rect 40628 30604 50988 30660
rect 51044 30604 51054 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 32162 30492 32172 30548
rect 32228 30492 33404 30548
rect 33460 30492 33470 30548
rect 21858 30380 21868 30436
rect 21924 30380 22428 30436
rect 22484 30380 23324 30436
rect 23380 30380 25228 30436
rect 25284 30380 27132 30436
rect 27188 30380 27198 30436
rect 38994 30380 39004 30436
rect 39060 30380 46508 30436
rect 46564 30380 46574 30436
rect 49186 30380 49196 30436
rect 49252 30380 49262 30436
rect 49196 30324 49252 30380
rect 26114 30268 26124 30324
rect 26180 30268 26908 30324
rect 26964 30268 26974 30324
rect 46806 30268 46844 30324
rect 46900 30268 46910 30324
rect 47702 30268 47740 30324
rect 47796 30268 47806 30324
rect 47954 30268 47964 30324
rect 48020 30268 49084 30324
rect 49140 30268 49252 30324
rect 53666 30268 53676 30324
rect 53732 30268 54572 30324
rect 54628 30268 54638 30324
rect 18386 30156 18396 30212
rect 18452 30156 19516 30212
rect 19572 30156 19582 30212
rect 21634 30156 21644 30212
rect 21700 30156 22316 30212
rect 22372 30156 22988 30212
rect 23044 30156 23054 30212
rect 26562 30156 26572 30212
rect 26628 30156 28140 30212
rect 28196 30156 28206 30212
rect 35186 30156 35196 30212
rect 35252 30156 35756 30212
rect 35812 30156 38220 30212
rect 38276 30156 38286 30212
rect 42018 30156 42028 30212
rect 42084 30156 42364 30212
rect 42420 30156 42430 30212
rect 46386 30156 46396 30212
rect 46452 30156 46956 30212
rect 47012 30156 47022 30212
rect 48738 30156 48748 30212
rect 48804 30156 48972 30212
rect 49028 30156 49038 30212
rect 51874 30156 51884 30212
rect 51940 30156 53116 30212
rect 53172 30156 53182 30212
rect 15698 30044 15708 30100
rect 15764 30044 16604 30100
rect 16660 30044 16670 30100
rect 22866 30044 22876 30100
rect 22932 30044 24108 30100
rect 24164 30044 24174 30100
rect 28466 30044 28476 30100
rect 28532 30044 29372 30100
rect 29428 30044 30604 30100
rect 30660 30044 30670 30100
rect 34626 30044 34636 30100
rect 34692 30044 43372 30100
rect 43428 30044 43438 30100
rect 45602 30044 45612 30100
rect 45668 30044 51548 30100
rect 51604 30044 51614 30100
rect 52994 30044 53004 30100
rect 53060 30044 53788 30100
rect 53844 30044 53854 30100
rect 16034 29932 16044 29988
rect 16100 29932 17388 29988
rect 17444 29932 17454 29988
rect 20066 29932 20076 29988
rect 20132 29932 25340 29988
rect 25396 29932 25406 29988
rect 43250 29932 43260 29988
rect 43316 29932 48076 29988
rect 48132 29932 48524 29988
rect 48580 29932 49420 29988
rect 49476 29932 49486 29988
rect 49634 29932 49644 29988
rect 49700 29932 51436 29988
rect 51492 29932 51502 29988
rect 52770 29932 52780 29988
rect 52836 29932 53564 29988
rect 53620 29932 53630 29988
rect 16146 29820 16156 29876
rect 16212 29820 17948 29876
rect 18004 29820 18014 29876
rect 38098 29820 38108 29876
rect 38164 29820 39228 29876
rect 39284 29820 45724 29876
rect 45780 29820 47292 29876
rect 47348 29820 50204 29876
rect 50260 29820 50270 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 18050 29708 18060 29764
rect 18116 29708 18844 29764
rect 18900 29708 18910 29764
rect 21858 29708 21868 29764
rect 21924 29708 23436 29764
rect 23492 29708 23502 29764
rect 26674 29708 26684 29764
rect 26740 29708 27020 29764
rect 27076 29708 27086 29764
rect 45798 29708 45836 29764
rect 45892 29708 45902 29764
rect 21746 29596 21756 29652
rect 21812 29596 28252 29652
rect 28308 29596 28318 29652
rect 33730 29596 33740 29652
rect 33796 29596 34076 29652
rect 34132 29596 35196 29652
rect 35252 29596 35262 29652
rect 46050 29596 46060 29652
rect 46116 29596 46956 29652
rect 47012 29596 47022 29652
rect 47394 29596 47404 29652
rect 47460 29596 49868 29652
rect 49924 29596 49934 29652
rect 15922 29484 15932 29540
rect 15988 29484 18060 29540
rect 18116 29484 18126 29540
rect 39106 29484 39116 29540
rect 39172 29484 39900 29540
rect 39956 29484 39966 29540
rect 45826 29484 45836 29540
rect 45892 29484 52892 29540
rect 52948 29484 52958 29540
rect 12226 29372 12236 29428
rect 12292 29372 13468 29428
rect 13524 29372 13534 29428
rect 24658 29372 24668 29428
rect 24724 29372 25452 29428
rect 25508 29372 25518 29428
rect 32274 29372 32284 29428
rect 32340 29372 33068 29428
rect 33124 29372 33134 29428
rect 33954 29372 33964 29428
rect 34020 29372 35308 29428
rect 35364 29372 35374 29428
rect 42242 29372 42252 29428
rect 42308 29372 43484 29428
rect 43540 29372 44716 29428
rect 44772 29372 45164 29428
rect 45220 29372 45724 29428
rect 45780 29372 45790 29428
rect 46610 29372 46620 29428
rect 46676 29372 47068 29428
rect 47124 29372 47134 29428
rect 53106 29372 53116 29428
rect 53172 29372 54796 29428
rect 54852 29372 54862 29428
rect 4274 29260 4284 29316
rect 4340 29260 5740 29316
rect 5796 29260 8316 29316
rect 8372 29260 8988 29316
rect 9044 29260 9054 29316
rect 15474 29260 15484 29316
rect 15540 29260 16828 29316
rect 16884 29260 16894 29316
rect 32498 29260 32508 29316
rect 32564 29260 33516 29316
rect 33572 29260 34524 29316
rect 34580 29260 34590 29316
rect 41682 29260 41692 29316
rect 41748 29260 44492 29316
rect 44548 29260 47404 29316
rect 47460 29260 47470 29316
rect 48290 29260 48300 29316
rect 48356 29260 49644 29316
rect 49700 29260 49710 29316
rect 53890 29260 53900 29316
rect 53956 29260 54460 29316
rect 54516 29260 54526 29316
rect 24658 29148 24668 29204
rect 24724 29148 27580 29204
rect 27636 29148 27646 29204
rect 45154 29148 45164 29204
rect 45220 29148 46396 29204
rect 46452 29148 47180 29204
rect 47236 29148 49756 29204
rect 49812 29148 49822 29204
rect 17154 29036 17164 29092
rect 17220 29036 17836 29092
rect 17892 29036 18620 29092
rect 18676 29036 18686 29092
rect 36978 29036 36988 29092
rect 37044 29036 37660 29092
rect 37716 29036 44268 29092
rect 44324 29036 44334 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 33058 28924 33068 28980
rect 33124 28924 33348 28980
rect 41122 28924 41132 28980
rect 41188 28924 43596 28980
rect 43652 28924 50428 28980
rect 53554 28924 53564 28980
rect 53620 28924 54236 28980
rect 54292 28924 54302 28980
rect 33292 28868 33348 28924
rect 50372 28868 50428 28924
rect 24322 28812 24332 28868
rect 24388 28812 25228 28868
rect 25284 28812 25294 28868
rect 26450 28812 26460 28868
rect 26516 28812 27804 28868
rect 27860 28812 27870 28868
rect 28242 28812 28252 28868
rect 28308 28812 29148 28868
rect 29204 28812 29214 28868
rect 33282 28812 33292 28868
rect 33348 28812 33358 28868
rect 43810 28812 43820 28868
rect 43876 28812 45500 28868
rect 45556 28812 46620 28868
rect 46676 28812 46686 28868
rect 50372 28812 51212 28868
rect 51268 28812 51772 28868
rect 51828 28812 51838 28868
rect 52780 28812 53676 28868
rect 53732 28812 55356 28868
rect 55412 28812 56252 28868
rect 56308 28812 56318 28868
rect 33842 28700 33852 28756
rect 33908 28700 34748 28756
rect 34804 28700 38668 28756
rect 41458 28700 41468 28756
rect 41524 28700 41916 28756
rect 41972 28700 41982 28756
rect 43362 28700 43372 28756
rect 43428 28700 44044 28756
rect 44100 28700 44828 28756
rect 44884 28700 44894 28756
rect 45378 28700 45388 28756
rect 45444 28700 46396 28756
rect 46452 28700 46462 28756
rect 38612 28644 38668 28700
rect 7858 28588 7868 28644
rect 7924 28588 8540 28644
rect 8596 28588 8606 28644
rect 12898 28588 12908 28644
rect 12964 28588 13468 28644
rect 13524 28588 13804 28644
rect 13860 28588 15484 28644
rect 15540 28588 15550 28644
rect 22754 28588 22764 28644
rect 22820 28588 23436 28644
rect 23492 28588 23502 28644
rect 24098 28588 24108 28644
rect 24164 28588 25228 28644
rect 25284 28588 25294 28644
rect 25442 28588 25452 28644
rect 25508 28588 27356 28644
rect 27412 28588 27422 28644
rect 33506 28588 33516 28644
rect 33572 28588 34076 28644
rect 34132 28588 34142 28644
rect 37202 28588 37212 28644
rect 37268 28588 38108 28644
rect 38164 28588 38174 28644
rect 38612 28588 39340 28644
rect 39396 28588 40572 28644
rect 40628 28588 40638 28644
rect 42578 28588 42588 28644
rect 42644 28588 46172 28644
rect 46228 28588 46238 28644
rect 52780 28532 52836 28812
rect 53778 28700 53788 28756
rect 53844 28700 54908 28756
rect 54964 28700 54974 28756
rect 54002 28588 54012 28644
rect 54068 28588 56476 28644
rect 56532 28588 56542 28644
rect 8642 28476 8652 28532
rect 8708 28476 10892 28532
rect 10948 28476 10958 28532
rect 18386 28476 18396 28532
rect 18452 28476 19180 28532
rect 19236 28476 19246 28532
rect 32946 28476 32956 28532
rect 33012 28476 33740 28532
rect 33796 28476 33806 28532
rect 44258 28476 44268 28532
rect 44324 28476 47292 28532
rect 47348 28476 47358 28532
rect 49970 28476 49980 28532
rect 50036 28476 51660 28532
rect 51716 28476 51726 28532
rect 52770 28476 52780 28532
rect 52836 28476 52846 28532
rect 19058 28364 19068 28420
rect 19124 28364 21420 28420
rect 21476 28364 21756 28420
rect 21812 28364 21822 28420
rect 32386 28364 32396 28420
rect 32452 28364 35308 28420
rect 35364 28364 36428 28420
rect 36484 28364 36494 28420
rect 42438 28364 42476 28420
rect 42532 28364 42542 28420
rect 43260 28364 45836 28420
rect 45892 28364 45902 28420
rect 46946 28364 46956 28420
rect 47012 28364 55468 28420
rect 55524 28364 55534 28420
rect 43260 28308 43316 28364
rect 45836 28308 45892 28364
rect 43250 28252 43260 28308
rect 43316 28252 43326 28308
rect 45836 28252 48860 28308
rect 48916 28252 49532 28308
rect 49588 28252 49598 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 55010 28140 55020 28196
rect 55076 28140 55692 28196
rect 55748 28140 55758 28196
rect 16818 28028 16828 28084
rect 16884 28028 17500 28084
rect 17556 28028 17566 28084
rect 38546 28028 38556 28084
rect 38612 28028 40348 28084
rect 40404 28028 40414 28084
rect 44930 28028 44940 28084
rect 44996 28028 50428 28084
rect 50484 28028 50494 28084
rect 50642 28028 50652 28084
rect 50708 28028 51660 28084
rect 51716 28028 51726 28084
rect 54114 28028 54124 28084
rect 54180 28028 56812 28084
rect 56868 28028 56878 28084
rect 31826 27916 31836 27972
rect 31892 27916 32284 27972
rect 32340 27916 35084 27972
rect 35140 27916 36540 27972
rect 36596 27916 36606 27972
rect 46722 27916 46732 27972
rect 46788 27916 46956 27972
rect 47012 27916 47022 27972
rect 51762 27916 51772 27972
rect 51828 27916 53788 27972
rect 53844 27916 54460 27972
rect 54516 27916 56588 27972
rect 56644 27916 56654 27972
rect 23986 27804 23996 27860
rect 24052 27804 26236 27860
rect 26292 27804 26302 27860
rect 32498 27804 32508 27860
rect 32564 27804 35532 27860
rect 35588 27804 35598 27860
rect 36082 27804 36092 27860
rect 36148 27804 37324 27860
rect 37380 27804 38556 27860
rect 38612 27804 38622 27860
rect 47842 27804 47852 27860
rect 47908 27804 52332 27860
rect 52388 27804 55020 27860
rect 55076 27804 55086 27860
rect 4722 27692 4732 27748
rect 4788 27692 5628 27748
rect 5684 27692 5694 27748
rect 18610 27692 18620 27748
rect 18676 27692 19740 27748
rect 19796 27692 22988 27748
rect 23044 27692 23436 27748
rect 23492 27692 28364 27748
rect 28420 27692 28812 27748
rect 28868 27692 28878 27748
rect 54226 27692 54236 27748
rect 54292 27692 55580 27748
rect 55636 27692 57708 27748
rect 57764 27692 57774 27748
rect 5954 27580 5964 27636
rect 6020 27580 7308 27636
rect 7364 27580 7374 27636
rect 17154 27580 17164 27636
rect 17220 27580 18956 27636
rect 19012 27580 19022 27636
rect 41234 27580 41244 27636
rect 41300 27580 41804 27636
rect 41860 27580 41870 27636
rect 49186 27580 49196 27636
rect 49252 27580 49980 27636
rect 50036 27580 50046 27636
rect 50418 27580 50428 27636
rect 50484 27580 51436 27636
rect 51492 27580 51660 27636
rect 51716 27580 54348 27636
rect 54404 27580 54414 27636
rect 21522 27468 21532 27524
rect 21588 27468 22092 27524
rect 22148 27468 22540 27524
rect 22596 27468 22606 27524
rect 33618 27468 33628 27524
rect 33684 27468 33964 27524
rect 34020 27468 34030 27524
rect 42018 27468 42028 27524
rect 42084 27468 42094 27524
rect 43026 27468 43036 27524
rect 43092 27468 43596 27524
rect 43652 27468 43662 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 42028 27412 42084 27468
rect 38882 27356 38892 27412
rect 38948 27356 40012 27412
rect 40068 27356 48188 27412
rect 48244 27356 48254 27412
rect 50754 27356 50764 27412
rect 50820 27356 51660 27412
rect 51716 27356 53228 27412
rect 53284 27356 53294 27412
rect 33702 27244 33740 27300
rect 33796 27244 34188 27300
rect 34244 27244 34254 27300
rect 37762 27244 37772 27300
rect 37828 27244 39564 27300
rect 39620 27244 39630 27300
rect 42130 27244 42140 27300
rect 42196 27244 42924 27300
rect 42980 27244 42990 27300
rect 45042 27244 45052 27300
rect 45108 27244 45836 27300
rect 45892 27244 45902 27300
rect 6962 27132 6972 27188
rect 7028 27132 8204 27188
rect 8260 27132 11116 27188
rect 11172 27132 11182 27188
rect 38322 27132 38332 27188
rect 38388 27132 40460 27188
rect 40516 27132 45276 27188
rect 45332 27132 45342 27188
rect 47394 27132 47404 27188
rect 47460 27132 48188 27188
rect 48244 27132 48254 27188
rect 50978 27132 50988 27188
rect 51044 27132 52780 27188
rect 52836 27132 52846 27188
rect 10210 27020 10220 27076
rect 10276 27020 10780 27076
rect 10836 27020 10846 27076
rect 20514 27020 20524 27076
rect 20580 27020 22540 27076
rect 22596 27020 22606 27076
rect 31602 27020 31612 27076
rect 31668 27020 32284 27076
rect 32340 27020 33292 27076
rect 33348 27020 33358 27076
rect 36418 27020 36428 27076
rect 36484 27020 36988 27076
rect 37044 27020 37054 27076
rect 38892 27020 40012 27076
rect 40068 27020 40078 27076
rect 40338 27020 40348 27076
rect 40404 27020 41916 27076
rect 41972 27020 41982 27076
rect 42242 27020 42252 27076
rect 42308 27020 42812 27076
rect 42868 27020 42878 27076
rect 44034 27020 44044 27076
rect 44100 27020 45724 27076
rect 45780 27020 45790 27076
rect 46610 27020 46620 27076
rect 46676 27020 48748 27076
rect 48804 27020 48814 27076
rect 51202 27020 51212 27076
rect 51268 27020 52332 27076
rect 52388 27020 53340 27076
rect 53396 27020 53406 27076
rect 33618 26908 33628 26964
rect 33684 26908 34524 26964
rect 34580 26908 34590 26964
rect 36194 26908 36204 26964
rect 36260 26908 37212 26964
rect 37268 26908 37436 26964
rect 37492 26908 37502 26964
rect 38892 26852 38948 27020
rect 43250 26908 43260 26964
rect 43316 26908 43484 26964
rect 43540 26908 43550 26964
rect 53676 26908 54460 26964
rect 54516 26908 54908 26964
rect 54964 26908 54974 26964
rect 53676 26852 53732 26908
rect 19516 26796 20076 26852
rect 20132 26796 20142 26852
rect 21746 26796 21756 26852
rect 21812 26796 22652 26852
rect 22708 26796 22718 26852
rect 29586 26796 29596 26852
rect 29652 26796 33180 26852
rect 33236 26796 33246 26852
rect 33506 26796 33516 26852
rect 33572 26796 33740 26852
rect 33796 26796 33806 26852
rect 34066 26796 34076 26852
rect 34132 26796 35644 26852
rect 35700 26796 35710 26852
rect 38630 26796 38668 26852
rect 38724 26796 38734 26852
rect 38882 26796 38892 26852
rect 38948 26796 38958 26852
rect 41234 26796 41244 26852
rect 41300 26796 43932 26852
rect 43988 26796 43998 26852
rect 46834 26796 46844 26852
rect 46900 26796 48524 26852
rect 48580 26796 48590 26852
rect 50372 26796 51996 26852
rect 52052 26796 52062 26852
rect 53666 26796 53676 26852
rect 53732 26796 53742 26852
rect 19516 26740 19572 26796
rect 50372 26740 50428 26796
rect 19506 26684 19516 26740
rect 19572 26684 19582 26740
rect 49858 26684 49868 26740
rect 49924 26684 50428 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 7074 26572 7084 26628
rect 7140 26572 8316 26628
rect 8372 26572 10108 26628
rect 10164 26572 10174 26628
rect 22418 26572 22428 26628
rect 22484 26572 23212 26628
rect 23268 26572 23278 26628
rect 41122 26572 41132 26628
rect 41188 26572 42476 26628
rect 42532 26572 42588 26628
rect 42644 26572 42654 26628
rect 11106 26460 11116 26516
rect 11172 26460 13916 26516
rect 13972 26460 13982 26516
rect 20626 26460 20636 26516
rect 20692 26460 21644 26516
rect 21700 26460 23548 26516
rect 23604 26460 23614 26516
rect 33618 26460 33628 26516
rect 33684 26460 34412 26516
rect 34468 26460 34478 26516
rect 45266 26460 45276 26516
rect 45332 26460 48636 26516
rect 48692 26460 48860 26516
rect 48916 26460 48926 26516
rect 51538 26460 51548 26516
rect 51604 26460 51884 26516
rect 51940 26460 51950 26516
rect 22530 26348 22540 26404
rect 22596 26348 22606 26404
rect 46050 26348 46060 26404
rect 46116 26348 46732 26404
rect 46788 26348 46798 26404
rect 47618 26348 47628 26404
rect 47684 26348 50316 26404
rect 50372 26348 53900 26404
rect 53956 26348 53966 26404
rect 22540 26292 22596 26348
rect 9650 26236 9660 26292
rect 9716 26236 12348 26292
rect 12404 26236 12414 26292
rect 22540 26236 23100 26292
rect 23156 26236 24332 26292
rect 24388 26236 25116 26292
rect 25172 26236 25182 26292
rect 28466 26236 28476 26292
rect 28532 26236 28700 26292
rect 28756 26236 28766 26292
rect 31602 26236 31612 26292
rect 31668 26236 32060 26292
rect 32116 26236 33516 26292
rect 33572 26236 33582 26292
rect 35298 26236 35308 26292
rect 35364 26236 35980 26292
rect 36036 26236 37100 26292
rect 37156 26236 37166 26292
rect 40114 26236 40124 26292
rect 40180 26236 41356 26292
rect 41412 26236 41916 26292
rect 41972 26236 41982 26292
rect 45378 26236 45388 26292
rect 45444 26236 46844 26292
rect 46900 26236 48972 26292
rect 49028 26236 49038 26292
rect 50950 26236 50988 26292
rect 51044 26236 51054 26292
rect 51314 26236 51324 26292
rect 51380 26236 52556 26292
rect 52612 26236 52622 26292
rect 51324 26180 51380 26236
rect 19506 26124 19516 26180
rect 19572 26124 21196 26180
rect 21252 26124 21262 26180
rect 23874 26124 23884 26180
rect 23940 26124 25340 26180
rect 25396 26124 25406 26180
rect 30482 26124 30492 26180
rect 30548 26124 33180 26180
rect 33236 26124 33246 26180
rect 37202 26124 37212 26180
rect 37268 26124 39900 26180
rect 39956 26124 39966 26180
rect 45938 26124 45948 26180
rect 46004 26124 51380 26180
rect 21634 26012 21644 26068
rect 21700 26012 22988 26068
rect 23044 26012 24892 26068
rect 24948 26012 26124 26068
rect 26180 26012 26190 26068
rect 32498 26012 32508 26068
rect 32564 26012 33068 26068
rect 33124 26012 33134 26068
rect 34514 26012 34524 26068
rect 34580 26012 35532 26068
rect 35588 26012 35598 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 42466 25788 42476 25844
rect 42532 25788 43484 25844
rect 43540 25788 45388 25844
rect 45444 25788 46172 25844
rect 46228 25788 47516 25844
rect 47572 25788 47582 25844
rect 50866 25788 50876 25844
rect 50932 25788 50942 25844
rect 7410 25676 7420 25732
rect 7476 25676 11452 25732
rect 11508 25676 11518 25732
rect 12226 25676 12236 25732
rect 12292 25676 12796 25732
rect 12852 25676 26908 25732
rect 8866 25564 8876 25620
rect 8932 25564 9884 25620
rect 9940 25564 11228 25620
rect 11284 25564 11294 25620
rect 13906 25564 13916 25620
rect 13972 25564 15484 25620
rect 15540 25564 15550 25620
rect 23538 25564 23548 25620
rect 23604 25564 24444 25620
rect 24500 25564 26684 25620
rect 26740 25564 26750 25620
rect 23986 25452 23996 25508
rect 24052 25452 25564 25508
rect 25620 25452 25630 25508
rect 10658 25340 10668 25396
rect 10724 25340 11564 25396
rect 11620 25340 11900 25396
rect 11956 25340 11966 25396
rect 12114 25340 12124 25396
rect 12180 25340 12908 25396
rect 12964 25340 14140 25396
rect 14196 25340 14206 25396
rect 14690 25340 14700 25396
rect 14756 25340 15260 25396
rect 15316 25340 15326 25396
rect 20290 25340 20300 25396
rect 20356 25340 22540 25396
rect 22596 25340 22606 25396
rect 24322 25340 24332 25396
rect 24388 25340 25340 25396
rect 25396 25340 25406 25396
rect 8082 25228 8092 25284
rect 8148 25228 10332 25284
rect 10388 25228 10398 25284
rect 11442 25228 11452 25284
rect 11508 25228 15148 25284
rect 18162 25228 18172 25284
rect 18228 25228 18732 25284
rect 18788 25228 18798 25284
rect 19628 25228 19964 25284
rect 20020 25228 20244 25284
rect 20738 25228 20748 25284
rect 20804 25228 21196 25284
rect 21252 25228 21262 25284
rect 21410 25228 21420 25284
rect 21476 25228 21980 25284
rect 22036 25228 22046 25284
rect 25106 25228 25116 25284
rect 25172 25228 25676 25284
rect 25732 25228 25742 25284
rect 15092 24836 15148 25228
rect 19628 25172 19684 25228
rect 16146 25116 16156 25172
rect 16212 25116 18396 25172
rect 18452 25116 18462 25172
rect 19058 25116 19068 25172
rect 19124 25116 19684 25172
rect 20188 25172 20244 25228
rect 20188 25116 26124 25172
rect 26180 25116 26190 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 26852 25060 26908 25676
rect 50876 25620 50932 25788
rect 52546 25676 52556 25732
rect 52612 25676 53900 25732
rect 53956 25676 53966 25732
rect 40114 25564 40124 25620
rect 40180 25564 42868 25620
rect 43586 25564 43596 25620
rect 43652 25564 44996 25620
rect 45826 25564 45836 25620
rect 45892 25564 46956 25620
rect 47012 25564 47516 25620
rect 47572 25564 47582 25620
rect 50866 25564 50876 25620
rect 50932 25564 51324 25620
rect 51380 25564 51390 25620
rect 52882 25564 52892 25620
rect 52948 25564 52958 25620
rect 42812 25508 42868 25564
rect 44940 25508 44996 25564
rect 52892 25508 52948 25564
rect 39890 25452 39900 25508
rect 39956 25452 40796 25508
rect 40852 25452 40862 25508
rect 41682 25452 41692 25508
rect 41748 25452 42252 25508
rect 42308 25452 42318 25508
rect 42802 25452 42812 25508
rect 42868 25452 43708 25508
rect 43764 25452 43774 25508
rect 44930 25452 44940 25508
rect 44996 25452 47292 25508
rect 47348 25452 47358 25508
rect 50642 25452 50652 25508
rect 50708 25452 51548 25508
rect 51604 25452 52948 25508
rect 28578 25340 28588 25396
rect 28644 25340 29372 25396
rect 29428 25340 29596 25396
rect 29652 25340 29662 25396
rect 32610 25340 32620 25396
rect 32676 25340 33628 25396
rect 33684 25340 33694 25396
rect 38658 25340 38668 25396
rect 38724 25340 41244 25396
rect 41300 25340 41310 25396
rect 44034 25340 44044 25396
rect 44100 25340 45724 25396
rect 45780 25340 45790 25396
rect 51650 25340 51660 25396
rect 51716 25340 51996 25396
rect 52052 25340 54460 25396
rect 54516 25340 54526 25396
rect 32050 25228 32060 25284
rect 32116 25228 33068 25284
rect 33124 25228 33134 25284
rect 41346 25228 41356 25284
rect 41412 25228 42028 25284
rect 42084 25228 42476 25284
rect 42532 25228 42542 25284
rect 44146 25228 44156 25284
rect 44212 25228 47740 25284
rect 47796 25228 47806 25284
rect 51426 25228 51436 25284
rect 51492 25228 52668 25284
rect 52724 25228 52734 25284
rect 33842 25116 33852 25172
rect 33908 25116 34972 25172
rect 35028 25116 36988 25172
rect 37044 25116 37884 25172
rect 37940 25116 37950 25172
rect 40898 25116 40908 25172
rect 40964 25116 42140 25172
rect 42196 25116 42206 25172
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 26852 25004 28924 25060
rect 28980 25004 28990 25060
rect 34290 25004 34300 25060
rect 34356 25004 41132 25060
rect 41188 25004 41198 25060
rect 47170 25004 47180 25060
rect 47236 25004 49196 25060
rect 49252 25004 49262 25060
rect 49410 25004 49420 25060
rect 49476 25004 50204 25060
rect 50260 25004 50270 25060
rect 16258 24892 16268 24948
rect 16324 24892 20748 24948
rect 20804 24892 20814 24948
rect 24658 24892 24668 24948
rect 24724 24892 26348 24948
rect 26404 24892 26414 24948
rect 32498 24892 32508 24948
rect 32564 24892 34636 24948
rect 34692 24892 34702 24948
rect 49522 24892 49532 24948
rect 49588 24892 50988 24948
rect 51044 24892 51054 24948
rect 15092 24780 18508 24836
rect 18564 24780 18574 24836
rect 23090 24780 23100 24836
rect 23156 24780 23548 24836
rect 23604 24780 23614 24836
rect 24546 24780 24556 24836
rect 24612 24780 25452 24836
rect 25508 24780 26684 24836
rect 26740 24780 26750 24836
rect 34402 24780 34412 24836
rect 34468 24780 35420 24836
rect 35476 24780 35486 24836
rect 38210 24780 38220 24836
rect 38276 24780 38556 24836
rect 38612 24780 38892 24836
rect 38948 24780 38958 24836
rect 40796 24780 41244 24836
rect 41300 24780 41310 24836
rect 49532 24780 49980 24836
rect 50036 24780 51100 24836
rect 51156 24780 51166 24836
rect 52546 24780 52556 24836
rect 52612 24780 53340 24836
rect 53396 24780 53406 24836
rect 40796 24724 40852 24780
rect 49532 24724 49588 24780
rect 15810 24668 15820 24724
rect 15876 24668 16268 24724
rect 16324 24668 29148 24724
rect 29204 24668 29214 24724
rect 33282 24668 33292 24724
rect 33348 24668 34076 24724
rect 34132 24668 34142 24724
rect 37986 24668 37996 24724
rect 38052 24668 40012 24724
rect 40068 24668 40078 24724
rect 40786 24668 40796 24724
rect 40852 24668 40862 24724
rect 41010 24668 41020 24724
rect 41076 24668 42700 24724
rect 42756 24668 42766 24724
rect 44940 24668 46508 24724
rect 46564 24668 46574 24724
rect 49074 24668 49084 24724
rect 49140 24668 49532 24724
rect 49588 24668 49598 24724
rect 50278 24668 50316 24724
rect 50372 24668 50382 24724
rect 50950 24668 50988 24724
rect 51044 24668 51054 24724
rect 51986 24668 51996 24724
rect 52052 24668 53676 24724
rect 53732 24668 53742 24724
rect 44940 24612 44996 24668
rect 51996 24612 52052 24668
rect 32274 24556 32284 24612
rect 32340 24556 33516 24612
rect 33572 24556 33582 24612
rect 38630 24556 38668 24612
rect 38724 24556 38734 24612
rect 44258 24556 44268 24612
rect 44324 24556 44940 24612
rect 44996 24556 45006 24612
rect 45938 24556 45948 24612
rect 46004 24556 47964 24612
rect 48020 24556 48030 24612
rect 48626 24556 48636 24612
rect 48692 24556 50092 24612
rect 50148 24556 52052 24612
rect 17938 24444 17948 24500
rect 18004 24444 18956 24500
rect 19012 24444 19628 24500
rect 19684 24444 19694 24500
rect 23650 24444 23660 24500
rect 23716 24444 25788 24500
rect 25844 24444 25854 24500
rect 48178 24444 48188 24500
rect 48244 24444 49084 24500
rect 49140 24444 50428 24500
rect 50484 24444 50494 24500
rect 39078 24332 39116 24388
rect 39172 24332 39182 24388
rect 47842 24332 47852 24388
rect 47908 24332 50204 24388
rect 50260 24332 50270 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 29138 24220 29148 24276
rect 29204 24220 30156 24276
rect 30212 24220 30222 24276
rect 46722 24220 46732 24276
rect 46788 24220 47180 24276
rect 47236 24220 47628 24276
rect 47684 24220 49196 24276
rect 49252 24220 49262 24276
rect 49858 24220 49868 24276
rect 49924 24220 53228 24276
rect 53284 24220 53294 24276
rect 35410 24108 35420 24164
rect 35476 24108 36316 24164
rect 36372 24108 36652 24164
rect 36708 24108 41804 24164
rect 41860 24108 41870 24164
rect 45602 24108 45612 24164
rect 45668 24108 47348 24164
rect 47292 24052 47348 24108
rect 7074 23996 7084 24052
rect 7140 23996 7532 24052
rect 7588 23996 8652 24052
rect 8708 23996 8718 24052
rect 9202 23996 9212 24052
rect 9268 23996 25340 24052
rect 25396 23996 26796 24052
rect 26852 23996 26862 24052
rect 35522 23996 35532 24052
rect 35588 23996 37324 24052
rect 37380 23996 37390 24052
rect 46386 23996 46396 24052
rect 46452 23996 47068 24052
rect 47124 23996 47134 24052
rect 47282 23996 47292 24052
rect 47348 23996 50764 24052
rect 50820 23996 50830 24052
rect 9212 23940 9268 23996
rect 7298 23884 7308 23940
rect 7364 23884 7756 23940
rect 7812 23884 9268 23940
rect 23090 23884 23100 23940
rect 23156 23884 24220 23940
rect 24276 23884 24892 23940
rect 24948 23884 25228 23940
rect 25284 23884 25294 23940
rect 37202 23884 37212 23940
rect 37268 23884 38332 23940
rect 38388 23884 38398 23940
rect 38612 23884 45164 23940
rect 45220 23884 45230 23940
rect 47394 23884 47404 23940
rect 47460 23884 49420 23940
rect 49476 23884 49486 23940
rect 50866 23884 50876 23940
rect 50932 23884 51436 23940
rect 51492 23884 51502 23940
rect 38612 23828 38668 23884
rect 17266 23772 17276 23828
rect 17332 23772 17724 23828
rect 17780 23772 18732 23828
rect 18788 23772 18798 23828
rect 19618 23772 19628 23828
rect 19684 23772 21532 23828
rect 21588 23772 21868 23828
rect 21924 23772 22764 23828
rect 22820 23772 22830 23828
rect 29362 23772 29372 23828
rect 29428 23772 31276 23828
rect 31332 23772 31342 23828
rect 35858 23772 35868 23828
rect 35924 23772 36204 23828
rect 36260 23772 37100 23828
rect 37156 23772 37166 23828
rect 37324 23772 38668 23828
rect 40898 23772 40908 23828
rect 40964 23772 41356 23828
rect 41412 23772 42028 23828
rect 42084 23772 42094 23828
rect 46498 23772 46508 23828
rect 46564 23772 48300 23828
rect 48356 23772 48366 23828
rect 48934 23772 48972 23828
rect 49028 23772 49038 23828
rect 49270 23772 49308 23828
rect 49364 23772 49374 23828
rect 49634 23772 49644 23828
rect 49700 23772 52780 23828
rect 52836 23772 52846 23828
rect 37324 23716 37380 23772
rect 48300 23716 48356 23772
rect 19282 23660 19292 23716
rect 19348 23660 19964 23716
rect 20020 23660 20300 23716
rect 20356 23660 20366 23716
rect 22866 23660 22876 23716
rect 22932 23660 24444 23716
rect 24500 23660 24510 23716
rect 34738 23660 34748 23716
rect 34804 23660 35644 23716
rect 35700 23660 37380 23716
rect 38434 23660 38444 23716
rect 38500 23660 40684 23716
rect 40740 23660 40750 23716
rect 41794 23660 41804 23716
rect 41860 23660 45388 23716
rect 45444 23660 45454 23716
rect 48300 23660 49868 23716
rect 49924 23660 49934 23716
rect 33842 23548 33852 23604
rect 33908 23548 36428 23604
rect 36484 23548 36494 23604
rect 38994 23548 39004 23604
rect 39060 23548 39564 23604
rect 39620 23548 40236 23604
rect 40292 23548 41692 23604
rect 41748 23548 43484 23604
rect 43540 23548 43550 23604
rect 48150 23548 48188 23604
rect 48244 23548 48254 23604
rect 49298 23548 49308 23604
rect 49364 23548 49532 23604
rect 49588 23548 49598 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 49970 23492 49980 23548
rect 50036 23492 50046 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 13682 23436 13692 23492
rect 13748 23436 18284 23492
rect 18340 23436 18350 23492
rect 20402 23436 20412 23492
rect 20468 23436 21308 23492
rect 21364 23436 22652 23492
rect 22708 23436 22718 23492
rect 23100 23436 23996 23492
rect 24052 23436 24062 23492
rect 38658 23436 38668 23492
rect 38724 23436 40012 23492
rect 40068 23436 40078 23492
rect 47058 23436 47068 23492
rect 47124 23436 47628 23492
rect 47684 23436 47694 23492
rect 47954 23436 47964 23492
rect 48020 23436 48524 23492
rect 48580 23436 48590 23492
rect 48962 23436 48972 23492
rect 49028 23436 49038 23492
rect 49980 23436 50092 23492
rect 50148 23436 50158 23492
rect 23100 23380 23156 23436
rect 4610 23324 4620 23380
rect 4676 23324 6524 23380
rect 6580 23324 6590 23380
rect 17490 23324 17500 23380
rect 17556 23324 18172 23380
rect 18228 23324 18620 23380
rect 18676 23324 18686 23380
rect 19506 23324 19516 23380
rect 19572 23324 19852 23380
rect 19908 23324 19918 23380
rect 20178 23324 20188 23380
rect 20244 23324 20748 23380
rect 20804 23324 20814 23380
rect 21186 23324 21196 23380
rect 21252 23324 21756 23380
rect 21812 23324 23100 23380
rect 23156 23324 23166 23380
rect 23314 23324 23324 23380
rect 23380 23324 25340 23380
rect 25396 23324 25406 23380
rect 34290 23324 34300 23380
rect 34356 23324 37772 23380
rect 37828 23324 37838 23380
rect 38546 23324 38556 23380
rect 38612 23324 39564 23380
rect 39620 23324 39630 23380
rect 39778 23324 39788 23380
rect 39844 23324 40796 23380
rect 40852 23324 42812 23380
rect 42868 23324 42878 23380
rect 48972 23268 49028 23436
rect 49634 23324 49644 23380
rect 49700 23324 50316 23380
rect 50372 23324 50382 23380
rect 50754 23324 50764 23380
rect 50820 23324 51660 23380
rect 51716 23324 52332 23380
rect 52388 23324 52398 23380
rect 12338 23212 12348 23268
rect 12404 23212 13916 23268
rect 13972 23212 13982 23268
rect 20066 23212 20076 23268
rect 20132 23212 20300 23268
rect 20356 23212 22204 23268
rect 22260 23212 22270 23268
rect 34178 23212 34188 23268
rect 34244 23212 36540 23268
rect 36596 23212 37212 23268
rect 37268 23212 37278 23268
rect 39666 23212 39676 23268
rect 39732 23212 41244 23268
rect 41300 23212 41310 23268
rect 42242 23212 42252 23268
rect 42308 23212 46060 23268
rect 46116 23212 46126 23268
rect 48626 23212 48636 23268
rect 48692 23212 49028 23268
rect 50372 23212 51436 23268
rect 51492 23212 51502 23268
rect 51874 23212 51884 23268
rect 51940 23212 53004 23268
rect 53060 23212 53070 23268
rect 50372 23156 50428 23212
rect 3266 23100 3276 23156
rect 3332 23100 5068 23156
rect 5124 23100 6412 23156
rect 6468 23100 9660 23156
rect 9716 23100 9726 23156
rect 18050 23100 18060 23156
rect 18116 23100 19516 23156
rect 19572 23100 22540 23156
rect 22596 23100 22606 23156
rect 33506 23100 33516 23156
rect 33572 23100 34748 23156
rect 34804 23100 35756 23156
rect 35812 23100 36652 23156
rect 36708 23100 38220 23156
rect 38276 23100 38286 23156
rect 43026 23100 43036 23156
rect 43092 23100 43820 23156
rect 43876 23100 43886 23156
rect 45378 23100 45388 23156
rect 45444 23100 49084 23156
rect 49140 23100 49150 23156
rect 49298 23100 49308 23156
rect 49364 23100 50428 23156
rect 50530 23100 50540 23156
rect 50596 23100 52108 23156
rect 52164 23100 52174 23156
rect 12562 22988 12572 23044
rect 12628 22988 13804 23044
rect 13860 22988 13870 23044
rect 15474 22988 15484 23044
rect 15540 22988 16716 23044
rect 16772 22988 16782 23044
rect 25666 22988 25676 23044
rect 25732 22988 26460 23044
rect 26516 22988 26526 23044
rect 28578 22988 28588 23044
rect 28644 22988 30716 23044
rect 30772 22988 30782 23044
rect 34626 22988 34636 23044
rect 34692 22988 35084 23044
rect 35140 22988 42140 23044
rect 42196 22988 42206 23044
rect 49858 22988 49868 23044
rect 49924 22988 50316 23044
rect 50372 22988 50382 23044
rect 50754 22988 50764 23044
rect 50820 22988 53340 23044
rect 53396 22988 53406 23044
rect 7970 22876 7980 22932
rect 8036 22876 13468 22932
rect 13524 22876 13534 22932
rect 42466 22876 42476 22932
rect 42532 22876 46284 22932
rect 46340 22876 46350 22932
rect 49074 22876 49084 22932
rect 49140 22876 50092 22932
rect 50148 22876 50158 22932
rect 51090 22876 51100 22932
rect 51156 22876 51772 22932
rect 51828 22876 51838 22932
rect 8978 22764 8988 22820
rect 9044 22764 9324 22820
rect 9380 22764 15148 22820
rect 15204 22764 16156 22820
rect 16212 22764 16222 22820
rect 49074 22764 49084 22820
rect 49140 22764 49756 22820
rect 49812 22764 49822 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 41122 22652 41132 22708
rect 41188 22652 42028 22708
rect 42084 22652 44828 22708
rect 44884 22652 44894 22708
rect 2706 22540 2716 22596
rect 2772 22540 5740 22596
rect 5796 22540 5806 22596
rect 6066 22540 6076 22596
rect 6132 22540 6860 22596
rect 6916 22540 8652 22596
rect 8708 22540 8718 22596
rect 13794 22540 13804 22596
rect 13860 22540 14252 22596
rect 14308 22540 23996 22596
rect 24052 22540 24444 22596
rect 24500 22540 24510 22596
rect 34962 22540 34972 22596
rect 35028 22540 36204 22596
rect 36260 22540 36270 22596
rect 36418 22540 36428 22596
rect 36484 22540 37436 22596
rect 37492 22540 38556 22596
rect 38612 22540 39116 22596
rect 39172 22540 39182 22596
rect 41234 22540 41244 22596
rect 41300 22540 42644 22596
rect 46050 22540 46060 22596
rect 46116 22540 50764 22596
rect 50820 22540 50830 22596
rect 42588 22484 42644 22540
rect 19842 22428 19852 22484
rect 19908 22428 23100 22484
rect 23156 22428 23166 22484
rect 32722 22428 32732 22484
rect 32788 22428 34188 22484
rect 34244 22428 35532 22484
rect 35588 22428 35598 22484
rect 37314 22428 37324 22484
rect 37380 22428 38892 22484
rect 38948 22428 39900 22484
rect 39956 22428 39966 22484
rect 40114 22428 40124 22484
rect 40180 22428 42028 22484
rect 42084 22428 42094 22484
rect 42578 22428 42588 22484
rect 42644 22428 46508 22484
rect 46564 22428 46574 22484
rect 47058 22428 47068 22484
rect 47124 22428 47852 22484
rect 47908 22428 48692 22484
rect 48850 22428 48860 22484
rect 48916 22428 51212 22484
rect 51268 22428 51278 22484
rect 42028 22372 42084 22428
rect 48636 22372 48692 22428
rect 6850 22316 6860 22372
rect 6916 22316 7644 22372
rect 7700 22316 7710 22372
rect 17714 22316 17724 22372
rect 17780 22316 18732 22372
rect 18788 22316 20412 22372
rect 20468 22316 20478 22372
rect 26450 22316 26460 22372
rect 26516 22316 27692 22372
rect 27748 22316 27758 22372
rect 40002 22316 40012 22372
rect 40068 22316 40684 22372
rect 40740 22316 40750 22372
rect 42028 22316 43148 22372
rect 43204 22316 43214 22372
rect 45500 22316 46060 22372
rect 46116 22316 46126 22372
rect 47618 22316 47628 22372
rect 47684 22316 48412 22372
rect 48468 22316 48478 22372
rect 48636 22316 50428 22372
rect 50484 22316 51996 22372
rect 52052 22316 52062 22372
rect 45500 22260 45556 22316
rect 12898 22204 12908 22260
rect 12964 22204 13468 22260
rect 13524 22204 15372 22260
rect 15428 22204 15438 22260
rect 17938 22204 17948 22260
rect 18004 22204 19068 22260
rect 19124 22204 19134 22260
rect 27010 22204 27020 22260
rect 27076 22204 28476 22260
rect 28532 22204 29820 22260
rect 29876 22204 29886 22260
rect 40226 22204 40236 22260
rect 40292 22204 43372 22260
rect 43428 22204 44268 22260
rect 44324 22204 45276 22260
rect 45332 22204 45342 22260
rect 45490 22204 45500 22260
rect 45556 22204 45566 22260
rect 47954 22204 47964 22260
rect 48020 22204 49420 22260
rect 49476 22204 49980 22260
rect 50036 22204 50046 22260
rect 26898 22092 26908 22148
rect 26964 22092 27580 22148
rect 27636 22092 27646 22148
rect 41010 22092 41020 22148
rect 41076 22092 42252 22148
rect 42308 22092 42318 22148
rect 42802 22092 42812 22148
rect 42868 22092 44044 22148
rect 44100 22092 45388 22148
rect 45444 22092 45454 22148
rect 46050 22092 46060 22148
rect 46116 22092 48636 22148
rect 48692 22092 48702 22148
rect 6850 21980 6860 22036
rect 6916 21980 15932 22036
rect 15988 21980 18284 22036
rect 18340 21980 18350 22036
rect 40114 21980 40124 22036
rect 40180 21980 42476 22036
rect 42532 21980 42542 22036
rect 47506 21980 47516 22036
rect 47572 21980 48748 22036
rect 48804 21980 49756 22036
rect 49812 21980 49822 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 4610 21868 4620 21924
rect 4676 21868 6076 21924
rect 6132 21868 7532 21924
rect 7588 21868 7598 21924
rect 20514 21868 20524 21924
rect 20580 21868 21532 21924
rect 21588 21868 21598 21924
rect 22306 21868 22316 21924
rect 22372 21868 23324 21924
rect 23380 21868 26684 21924
rect 26740 21868 26750 21924
rect 33282 21868 33292 21924
rect 33348 21868 34972 21924
rect 35028 21868 36988 21924
rect 37044 21868 37772 21924
rect 37828 21868 37838 21924
rect 24556 21812 24612 21868
rect 8754 21756 8764 21812
rect 8820 21756 9884 21812
rect 9940 21756 9950 21812
rect 24546 21756 24556 21812
rect 24612 21756 24622 21812
rect 26562 21756 26572 21812
rect 26628 21756 27524 21812
rect 29698 21756 29708 21812
rect 29764 21756 30492 21812
rect 30548 21756 30558 21812
rect 47842 21756 47852 21812
rect 47908 21756 49644 21812
rect 49700 21756 49710 21812
rect 27468 21700 27524 21756
rect 8866 21644 8876 21700
rect 8932 21644 10108 21700
rect 10164 21644 10174 21700
rect 11218 21644 11228 21700
rect 11284 21644 11900 21700
rect 11956 21644 11966 21700
rect 18386 21644 18396 21700
rect 18452 21644 19964 21700
rect 20020 21644 20030 21700
rect 23174 21644 23212 21700
rect 23268 21644 23278 21700
rect 24658 21644 24668 21700
rect 24724 21644 26908 21700
rect 27458 21644 27468 21700
rect 27524 21644 27534 21700
rect 30034 21644 30044 21700
rect 30100 21644 30380 21700
rect 30436 21644 30446 21700
rect 39890 21644 39900 21700
rect 39956 21644 46172 21700
rect 46228 21644 46238 21700
rect 47282 21644 47292 21700
rect 47348 21644 47740 21700
rect 47796 21644 47806 21700
rect 26852 21588 26908 21644
rect 8530 21532 8540 21588
rect 8596 21532 9772 21588
rect 9828 21532 9838 21588
rect 12226 21532 12236 21588
rect 12292 21532 12572 21588
rect 12628 21532 14476 21588
rect 14532 21532 14542 21588
rect 20178 21532 20188 21588
rect 20244 21532 20860 21588
rect 20916 21532 21868 21588
rect 21924 21532 21934 21588
rect 24882 21532 24892 21588
rect 24948 21532 25452 21588
rect 25508 21532 25518 21588
rect 26852 21532 33740 21588
rect 33796 21532 35644 21588
rect 35700 21532 35710 21588
rect 41234 21532 41244 21588
rect 41300 21532 43036 21588
rect 43092 21532 43102 21588
rect 47730 21532 47740 21588
rect 47796 21532 48972 21588
rect 49028 21532 49644 21588
rect 49700 21532 49710 21588
rect 7858 21420 7868 21476
rect 7924 21420 8652 21476
rect 8708 21420 8718 21476
rect 9650 21420 9660 21476
rect 9716 21420 12348 21476
rect 12404 21420 12414 21476
rect 14690 21420 14700 21476
rect 14756 21420 15260 21476
rect 15316 21420 15326 21476
rect 16706 21420 16716 21476
rect 16772 21420 16940 21476
rect 16996 21420 17500 21476
rect 17556 21420 25116 21476
rect 25172 21420 25182 21476
rect 25452 21420 26572 21476
rect 26628 21420 26638 21476
rect 40226 21420 40236 21476
rect 40292 21420 41804 21476
rect 41860 21420 41870 21476
rect 43922 21420 43932 21476
rect 43988 21420 49084 21476
rect 49140 21420 49150 21476
rect 14700 21364 14756 21420
rect 25452 21364 25508 21420
rect 4610 21308 4620 21364
rect 4676 21308 7644 21364
rect 7700 21308 7710 21364
rect 11554 21308 11564 21364
rect 11620 21308 14756 21364
rect 21634 21308 21644 21364
rect 21700 21308 22092 21364
rect 22148 21308 22158 21364
rect 25442 21308 25452 21364
rect 25508 21308 25518 21364
rect 25778 21308 25788 21364
rect 25844 21308 26124 21364
rect 26180 21308 26190 21364
rect 28690 21308 28700 21364
rect 28756 21308 29036 21364
rect 29092 21308 29102 21364
rect 32386 21308 32396 21364
rect 32452 21308 33516 21364
rect 33572 21308 33582 21364
rect 44258 21308 44268 21364
rect 44324 21308 49532 21364
rect 49588 21308 49598 21364
rect 7410 21196 7420 21252
rect 7476 21196 12796 21252
rect 12852 21196 17612 21252
rect 17668 21196 17678 21252
rect 18050 21196 18060 21252
rect 18116 21196 18508 21252
rect 18564 21196 28588 21252
rect 28644 21196 28654 21252
rect 48262 21196 48300 21252
rect 48356 21196 48366 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 18946 21084 18956 21140
rect 19012 21084 22204 21140
rect 22260 21084 23324 21140
rect 23380 21084 23390 21140
rect 7970 20972 7980 21028
rect 8036 20972 8540 21028
rect 8596 20972 8606 21028
rect 8978 20972 8988 21028
rect 9044 20972 14364 21028
rect 14420 20972 14430 21028
rect 17378 20972 17388 21028
rect 17444 20972 17836 21028
rect 17892 20972 18172 21028
rect 18228 20972 29708 21028
rect 29764 20972 29774 21028
rect 8866 20860 8876 20916
rect 8932 20860 8942 20916
rect 28578 20860 28588 20916
rect 28644 20860 29148 20916
rect 29204 20860 29214 20916
rect 44930 20860 44940 20916
rect 44996 20860 46844 20916
rect 46900 20860 47180 20916
rect 47236 20860 48636 20916
rect 48692 20860 49868 20916
rect 49924 20860 49934 20916
rect 8876 20804 8932 20860
rect 8530 20748 8540 20804
rect 8596 20748 8932 20804
rect 12898 20748 12908 20804
rect 12964 20748 13580 20804
rect 13636 20748 13646 20804
rect 14354 20748 14364 20804
rect 14420 20748 15260 20804
rect 15316 20748 15326 20804
rect 20290 20748 20300 20804
rect 20356 20748 24556 20804
rect 24612 20748 24622 20804
rect 14364 20692 14420 20748
rect 2706 20636 2716 20692
rect 2772 20636 3836 20692
rect 3892 20636 3902 20692
rect 4722 20636 4732 20692
rect 4788 20636 6748 20692
rect 6804 20636 6814 20692
rect 12338 20636 12348 20692
rect 12404 20636 12572 20692
rect 12628 20636 14420 20692
rect 19954 20636 19964 20692
rect 20020 20636 21308 20692
rect 21364 20636 21374 20692
rect 12674 20524 12684 20580
rect 12740 20524 14700 20580
rect 14756 20524 14766 20580
rect 15092 20524 18620 20580
rect 18676 20524 18686 20580
rect 39106 20524 39116 20580
rect 39172 20524 41580 20580
rect 41636 20524 41646 20580
rect 15092 20468 15148 20524
rect 4946 20412 4956 20468
rect 5012 20412 7756 20468
rect 7812 20412 15148 20468
rect 18274 20412 18284 20468
rect 18340 20412 19628 20468
rect 19684 20412 19694 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 23426 20300 23436 20356
rect 23492 20300 27132 20356
rect 27188 20300 27198 20356
rect 28242 20300 28252 20356
rect 28308 20300 29484 20356
rect 29540 20300 29550 20356
rect 29810 20300 29820 20356
rect 29876 20300 35532 20356
rect 35588 20300 35598 20356
rect 29484 20244 29540 20300
rect 14802 20188 14812 20244
rect 14868 20188 14878 20244
rect 17602 20188 17612 20244
rect 17668 20188 20860 20244
rect 20916 20188 20926 20244
rect 21074 20188 21084 20244
rect 21140 20188 22204 20244
rect 22260 20188 22764 20244
rect 22820 20188 23212 20244
rect 23268 20188 23548 20244
rect 25666 20188 25676 20244
rect 25732 20188 26236 20244
rect 26292 20188 26302 20244
rect 29484 20188 30044 20244
rect 30100 20188 34076 20244
rect 34132 20188 34142 20244
rect 14812 20132 14868 20188
rect 23492 20132 23548 20188
rect 14812 20076 15484 20132
rect 15540 20076 15550 20132
rect 20178 20076 20188 20132
rect 20244 20076 21308 20132
rect 21364 20076 21980 20132
rect 22036 20076 22046 20132
rect 22390 20076 22428 20132
rect 22484 20076 22494 20132
rect 23492 20076 23772 20132
rect 23828 20076 23838 20132
rect 25218 20076 25228 20132
rect 25284 20076 26124 20132
rect 26180 20076 26190 20132
rect 27010 20076 27020 20132
rect 27076 20076 28924 20132
rect 28980 20076 28990 20132
rect 8978 19964 8988 20020
rect 9044 19964 14588 20020
rect 14644 19964 14654 20020
rect 15026 19964 15036 20020
rect 15092 19964 15708 20020
rect 15764 19964 15774 20020
rect 16594 19964 16604 20020
rect 16660 19964 17388 20020
rect 17444 19964 17454 20020
rect 21746 19964 21756 20020
rect 21812 19964 22988 20020
rect 23044 19964 23054 20020
rect 23426 19964 23436 20020
rect 23492 19964 29484 20020
rect 29540 19964 29550 20020
rect 6850 19852 6860 19908
rect 6916 19852 7644 19908
rect 7700 19852 9548 19908
rect 9604 19852 9614 19908
rect 21970 19852 21980 19908
rect 22036 19852 22652 19908
rect 22708 19852 22718 19908
rect 24658 19852 24668 19908
rect 24724 19852 25564 19908
rect 25620 19852 25630 19908
rect 35410 19852 35420 19908
rect 35476 19852 37100 19908
rect 37156 19852 37166 19908
rect 38546 19852 38556 19908
rect 38612 19852 39788 19908
rect 39844 19852 42140 19908
rect 42196 19852 42206 19908
rect 7522 19740 7532 19796
rect 7588 19740 7980 19796
rect 8036 19740 11564 19796
rect 11620 19740 13692 19796
rect 13748 19740 13758 19796
rect 14914 19740 14924 19796
rect 14980 19740 15932 19796
rect 15988 19740 17612 19796
rect 17668 19740 17678 19796
rect 19394 19740 19404 19796
rect 19460 19740 20412 19796
rect 20468 19740 20478 19796
rect 28466 19740 28476 19796
rect 28532 19740 29260 19796
rect 29316 19740 29326 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 22166 19516 22204 19572
rect 22260 19516 22270 19572
rect 12786 19404 12796 19460
rect 12852 19404 14476 19460
rect 14532 19404 14542 19460
rect 16482 19404 16492 19460
rect 16548 19404 20300 19460
rect 20356 19404 20366 19460
rect 8194 19292 8204 19348
rect 8260 19292 21084 19348
rect 21140 19292 21150 19348
rect 21634 19292 21644 19348
rect 21700 19292 24220 19348
rect 24276 19292 24286 19348
rect 25442 19292 25452 19348
rect 25508 19292 27580 19348
rect 27636 19292 27646 19348
rect 33506 19292 33516 19348
rect 33572 19292 34636 19348
rect 34692 19292 34702 19348
rect 15026 19180 15036 19236
rect 15092 19180 15708 19236
rect 15764 19180 15774 19236
rect 16706 19180 16716 19236
rect 16772 19180 25004 19236
rect 25060 19180 25070 19236
rect 7298 19068 7308 19124
rect 7364 19068 8316 19124
rect 8372 19068 8652 19124
rect 8708 19068 8718 19124
rect 22082 19068 22092 19124
rect 22148 19068 22428 19124
rect 22484 19068 22494 19124
rect 25218 19068 25228 19124
rect 25284 19068 25676 19124
rect 25732 19068 26404 19124
rect 26348 19012 26404 19068
rect 5058 18956 5068 19012
rect 5124 18956 5740 19012
rect 5796 18956 8092 19012
rect 8148 18956 8158 19012
rect 10098 18956 10108 19012
rect 10164 18956 13804 19012
rect 13860 18956 13870 19012
rect 26338 18956 26348 19012
rect 26404 18956 26414 19012
rect 27010 18956 27020 19012
rect 27076 18956 33740 19012
rect 33796 18956 35308 19012
rect 35364 18956 35374 19012
rect 36978 18956 36988 19012
rect 37044 18956 37548 19012
rect 37604 18956 38220 19012
rect 38276 18956 38286 19012
rect 25666 18844 25676 18900
rect 25732 18844 26460 18900
rect 26516 18844 26526 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 24210 18732 24220 18788
rect 24276 18732 27804 18788
rect 27860 18732 27870 18788
rect 6850 18620 6860 18676
rect 6916 18620 9548 18676
rect 9604 18620 9614 18676
rect 21186 18620 21196 18676
rect 21252 18620 27692 18676
rect 27748 18620 27758 18676
rect 28914 18620 28924 18676
rect 28980 18620 30156 18676
rect 30212 18620 30222 18676
rect 6738 18508 6748 18564
rect 6804 18508 7980 18564
rect 8036 18508 8046 18564
rect 9426 18508 9436 18564
rect 9492 18508 13356 18564
rect 13412 18508 13422 18564
rect 13570 18508 13580 18564
rect 13636 18508 13646 18564
rect 26852 18508 33292 18564
rect 33348 18508 33358 18564
rect 13580 18452 13636 18508
rect 26852 18452 26908 18508
rect 2818 18396 2828 18452
rect 2884 18396 5628 18452
rect 5684 18396 5694 18452
rect 5954 18396 5964 18452
rect 6020 18396 8876 18452
rect 8932 18396 8942 18452
rect 9090 18396 9100 18452
rect 9156 18396 9996 18452
rect 10052 18396 10062 18452
rect 10210 18396 10220 18452
rect 10276 18396 11116 18452
rect 11172 18396 11182 18452
rect 11442 18396 11452 18452
rect 11508 18396 12460 18452
rect 12516 18396 12526 18452
rect 12786 18396 12796 18452
rect 12852 18396 13636 18452
rect 17490 18396 17500 18452
rect 17556 18396 18284 18452
rect 18340 18396 21308 18452
rect 21364 18396 21644 18452
rect 21700 18396 21710 18452
rect 22092 18396 25228 18452
rect 25284 18396 25294 18452
rect 26450 18396 26460 18452
rect 26516 18396 26908 18452
rect 27682 18396 27692 18452
rect 27748 18396 28028 18452
rect 28084 18396 28094 18452
rect 5964 18340 6020 18396
rect 22092 18340 22148 18396
rect 4946 18284 4956 18340
rect 5012 18284 6020 18340
rect 12898 18284 12908 18340
rect 12964 18284 14476 18340
rect 14532 18284 14542 18340
rect 16146 18284 16156 18340
rect 16212 18284 17948 18340
rect 18004 18284 18396 18340
rect 18452 18284 22148 18340
rect 24658 18284 24668 18340
rect 24724 18284 31668 18340
rect 31826 18284 31836 18340
rect 31892 18284 32284 18340
rect 32340 18284 33628 18340
rect 33684 18284 34300 18340
rect 34356 18284 34860 18340
rect 34916 18284 36988 18340
rect 37044 18284 37054 18340
rect 31612 18228 31668 18284
rect 9650 18172 9660 18228
rect 9716 18172 13244 18228
rect 13300 18172 13310 18228
rect 21186 18172 21196 18228
rect 21252 18172 24892 18228
rect 24948 18172 24958 18228
rect 25442 18172 25452 18228
rect 25508 18172 26348 18228
rect 26404 18172 27244 18228
rect 27300 18172 27310 18228
rect 31612 18172 32732 18228
rect 32788 18172 32798 18228
rect 10434 18060 10444 18116
rect 10500 18060 18172 18116
rect 18228 18060 18238 18116
rect 21970 18060 21980 18116
rect 22036 18060 25900 18116
rect 25956 18060 26796 18116
rect 26852 18060 26862 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 11106 17948 11116 18004
rect 11172 17948 13468 18004
rect 13524 17948 13534 18004
rect 15586 17948 15596 18004
rect 15652 17948 16044 18004
rect 16100 17948 16110 18004
rect 3602 17836 3612 17892
rect 3668 17836 5740 17892
rect 5796 17836 5806 17892
rect 11890 17836 11900 17892
rect 11956 17836 12572 17892
rect 12628 17836 12638 17892
rect 15138 17836 15148 17892
rect 15204 17836 16940 17892
rect 16996 17836 23212 17892
rect 23268 17836 23884 17892
rect 23940 17836 23950 17892
rect 25554 17836 25564 17892
rect 25620 17836 26012 17892
rect 26068 17836 26078 17892
rect 6402 17724 6412 17780
rect 6468 17724 7084 17780
rect 7140 17724 9548 17780
rect 9604 17724 9614 17780
rect 12898 17724 12908 17780
rect 12964 17724 15372 17780
rect 15428 17724 15438 17780
rect 16146 17724 16156 17780
rect 16212 17724 18060 17780
rect 18116 17724 18126 17780
rect 14690 17612 14700 17668
rect 14756 17612 15148 17668
rect 15204 17612 15214 17668
rect 15586 17612 15596 17668
rect 15652 17612 16604 17668
rect 16660 17612 25788 17668
rect 25844 17612 26572 17668
rect 26628 17612 26638 17668
rect 6402 17500 6412 17556
rect 6468 17500 7868 17556
rect 7924 17500 7934 17556
rect 8082 17500 8092 17556
rect 8148 17500 8988 17556
rect 9044 17500 9054 17556
rect 9202 17500 9212 17556
rect 9268 17500 10668 17556
rect 10724 17500 15148 17556
rect 15204 17500 15214 17556
rect 15596 17444 15652 17612
rect 23538 17500 23548 17556
rect 23604 17500 27916 17556
rect 27972 17500 27982 17556
rect 36082 17500 36092 17556
rect 36148 17500 37436 17556
rect 37492 17500 37502 17556
rect 8306 17388 8316 17444
rect 8372 17388 14364 17444
rect 14420 17388 14430 17444
rect 14690 17388 14700 17444
rect 14756 17388 15652 17444
rect 25106 17388 25116 17444
rect 25172 17388 27356 17444
rect 27412 17388 27422 17444
rect 27794 17388 27804 17444
rect 27860 17388 29820 17444
rect 29876 17388 29886 17444
rect 9202 17276 9212 17332
rect 9268 17276 16156 17332
rect 16212 17276 16222 17332
rect 21634 17276 21644 17332
rect 21700 17276 21980 17332
rect 22036 17276 22046 17332
rect 24658 17276 24668 17332
rect 24724 17276 25508 17332
rect 27122 17276 27132 17332
rect 27188 17276 28252 17332
rect 28308 17276 28318 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 25452 17220 25508 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 13906 17164 13916 17220
rect 13972 17164 14924 17220
rect 14980 17164 19684 17220
rect 19628 17108 19684 17164
rect 21644 17164 23772 17220
rect 23828 17164 23838 17220
rect 24322 17164 24332 17220
rect 24388 17164 25228 17220
rect 25284 17164 25294 17220
rect 25452 17164 26908 17220
rect 26964 17164 26974 17220
rect 27206 17164 27244 17220
rect 27300 17164 27310 17220
rect 21644 17108 21700 17164
rect 15092 17052 16492 17108
rect 16548 17052 16558 17108
rect 19628 17052 21700 17108
rect 21858 17052 21868 17108
rect 21924 17052 22652 17108
rect 22708 17052 25340 17108
rect 25396 17052 26460 17108
rect 26516 17052 26526 17108
rect 27458 17052 27468 17108
rect 27524 17052 27580 17108
rect 27636 17052 27646 17108
rect 15092 16996 15148 17052
rect 6962 16940 6972 16996
rect 7028 16940 7868 16996
rect 7924 16940 7934 16996
rect 14802 16940 14812 16996
rect 14868 16940 15148 16996
rect 16594 16940 16604 16996
rect 16660 16940 17500 16996
rect 17556 16940 17566 16996
rect 17826 16940 17836 16996
rect 17892 16940 20356 16996
rect 21522 16940 21532 16996
rect 21588 16940 23884 16996
rect 23940 16940 24668 16996
rect 24724 16940 24734 16996
rect 26002 16940 26012 16996
rect 26068 16940 31276 16996
rect 31332 16940 31342 16996
rect 20300 16884 20356 16940
rect 6066 16828 6076 16884
rect 6132 16828 7308 16884
rect 7364 16828 7644 16884
rect 7700 16828 7710 16884
rect 10322 16828 10332 16884
rect 10388 16828 11116 16884
rect 11172 16828 11182 16884
rect 12450 16828 12460 16884
rect 12516 16828 13020 16884
rect 13076 16828 13916 16884
rect 13972 16828 13982 16884
rect 14242 16828 14252 16884
rect 14308 16828 15484 16884
rect 15540 16828 17948 16884
rect 18004 16828 20244 16884
rect 20300 16828 24556 16884
rect 24612 16828 24622 16884
rect 25218 16828 25228 16884
rect 25284 16828 25294 16884
rect 25638 16828 25676 16884
rect 25732 16828 25742 16884
rect 26898 16828 26908 16884
rect 26964 16828 27002 16884
rect 27542 16828 27580 16884
rect 27636 16828 27646 16884
rect 29810 16828 29820 16884
rect 29876 16828 31948 16884
rect 32004 16828 32014 16884
rect 20188 16772 20244 16828
rect 25228 16772 25284 16828
rect 5954 16716 5964 16772
rect 6020 16716 7420 16772
rect 7476 16716 7486 16772
rect 14578 16716 14588 16772
rect 14644 16716 15148 16772
rect 15204 16716 15214 16772
rect 16818 16716 16828 16772
rect 16884 16716 17612 16772
rect 17668 16716 17678 16772
rect 18162 16716 18172 16772
rect 18228 16716 18956 16772
rect 19012 16716 19022 16772
rect 20188 16716 23660 16772
rect 23716 16716 23726 16772
rect 23996 16716 26124 16772
rect 26180 16716 26190 16772
rect 23996 16660 24052 16716
rect 2706 16604 2716 16660
rect 2772 16604 5740 16660
rect 5796 16604 5806 16660
rect 12898 16604 12908 16660
rect 12964 16604 14364 16660
rect 14420 16604 14430 16660
rect 16706 16604 16716 16660
rect 16772 16604 24052 16660
rect 24210 16604 24220 16660
rect 24276 16604 25676 16660
rect 25732 16604 25742 16660
rect 26786 16604 26796 16660
rect 26852 16604 27468 16660
rect 27524 16604 27534 16660
rect 31602 16604 31612 16660
rect 31668 16604 35084 16660
rect 35140 16604 36428 16660
rect 36484 16604 36494 16660
rect 9314 16492 9324 16548
rect 9380 16492 9772 16548
rect 9828 16492 17388 16548
rect 17444 16492 17454 16548
rect 19842 16492 19852 16548
rect 19908 16492 21196 16548
rect 21252 16492 29596 16548
rect 29652 16492 29662 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 17388 16436 17444 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 13794 16380 13804 16436
rect 13860 16380 14588 16436
rect 14644 16380 14654 16436
rect 17388 16380 22764 16436
rect 22820 16380 23436 16436
rect 23492 16380 23502 16436
rect 24994 16380 25004 16436
rect 25060 16380 25676 16436
rect 25732 16380 25742 16436
rect 30818 16380 30828 16436
rect 30884 16380 32956 16436
rect 33012 16380 33022 16436
rect 4610 16268 4620 16324
rect 4676 16268 6076 16324
rect 6132 16268 6142 16324
rect 11666 16268 11676 16324
rect 11732 16268 12124 16324
rect 12180 16268 12190 16324
rect 16034 16268 16044 16324
rect 16100 16268 16380 16324
rect 16436 16268 16446 16324
rect 18274 16268 18284 16324
rect 18340 16268 20972 16324
rect 21028 16268 21038 16324
rect 25452 16268 26684 16324
rect 26740 16268 26750 16324
rect 28130 16268 28140 16324
rect 28196 16268 30044 16324
rect 30100 16268 30110 16324
rect 13346 16156 13356 16212
rect 13412 16156 15820 16212
rect 15876 16156 19012 16212
rect 20626 16156 20636 16212
rect 20692 16156 21420 16212
rect 21476 16156 21486 16212
rect 13570 16044 13580 16100
rect 13636 16044 14140 16100
rect 14196 16044 14644 16100
rect 14802 16044 14812 16100
rect 14868 16044 16828 16100
rect 16884 16044 18060 16100
rect 18116 16044 18126 16100
rect 14588 15988 14644 16044
rect 18956 15988 19012 16156
rect 25452 16100 25508 16268
rect 26114 16156 26124 16212
rect 26180 16156 26190 16212
rect 30370 16156 30380 16212
rect 30436 16156 30828 16212
rect 30884 16156 31836 16212
rect 31892 16156 31902 16212
rect 26124 16100 26180 16156
rect 23762 16044 23772 16100
rect 23828 16044 25004 16100
rect 25060 16044 25070 16100
rect 25442 16044 25452 16100
rect 25508 16044 25518 16100
rect 25666 16044 25676 16100
rect 25732 16044 25788 16100
rect 25844 16044 25854 16100
rect 26124 16044 26684 16100
rect 26740 16044 26750 16100
rect 27010 16044 27020 16100
rect 27076 16044 27804 16100
rect 27860 16044 27870 16100
rect 32722 16044 32732 16100
rect 32788 16044 34748 16100
rect 34804 16044 35532 16100
rect 35588 16044 35598 16100
rect 6850 15932 6860 15988
rect 6916 15932 7420 15988
rect 7476 15932 7486 15988
rect 7746 15932 7756 15988
rect 7812 15932 10444 15988
rect 10500 15932 10892 15988
rect 10948 15932 11844 15988
rect 12450 15932 12460 15988
rect 12516 15932 14364 15988
rect 14420 15932 14430 15988
rect 14588 15932 15260 15988
rect 15316 15932 15326 15988
rect 18946 15932 18956 15988
rect 19012 15932 20412 15988
rect 20468 15932 20478 15988
rect 24210 15932 24220 15988
rect 24276 15932 24556 15988
rect 24612 15932 24622 15988
rect 25330 15932 25340 15988
rect 25396 15932 27356 15988
rect 27412 15932 28028 15988
rect 28084 15932 28094 15988
rect 11788 15876 11844 15932
rect 8306 15820 8316 15876
rect 8372 15820 11564 15876
rect 11620 15820 11630 15876
rect 11788 15820 15148 15876
rect 15204 15820 15214 15876
rect 16482 15820 16492 15876
rect 16548 15820 17164 15876
rect 17220 15820 22148 15876
rect 24770 15820 24780 15876
rect 24836 15820 26684 15876
rect 26740 15820 26750 15876
rect 36082 15820 36092 15876
rect 36148 15820 37548 15876
rect 37604 15820 37614 15876
rect 22092 15764 22148 15820
rect 14354 15708 14364 15764
rect 14420 15708 18732 15764
rect 18788 15708 19180 15764
rect 19236 15708 19246 15764
rect 22092 15708 24892 15764
rect 24948 15708 25676 15764
rect 25732 15708 25742 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 15138 15596 15148 15652
rect 15204 15596 16380 15652
rect 16436 15596 17052 15652
rect 17108 15596 17118 15652
rect 23314 15596 23324 15652
rect 23380 15596 25788 15652
rect 25844 15596 25854 15652
rect 26114 15596 26124 15652
rect 26180 15596 26684 15652
rect 26740 15596 26750 15652
rect 27458 15596 27468 15652
rect 27524 15596 33852 15652
rect 33908 15596 33918 15652
rect 7634 15484 7644 15540
rect 7700 15484 12796 15540
rect 12852 15484 13468 15540
rect 13524 15484 13534 15540
rect 23650 15484 23660 15540
rect 23716 15484 25004 15540
rect 25060 15484 25070 15540
rect 25452 15484 28364 15540
rect 28420 15484 28430 15540
rect 32498 15484 32508 15540
rect 32564 15484 33404 15540
rect 33460 15484 33628 15540
rect 33684 15484 33694 15540
rect 12002 15372 12012 15428
rect 12068 15372 13356 15428
rect 13412 15372 13422 15428
rect 19170 15372 19180 15428
rect 19236 15372 20524 15428
rect 20580 15372 20590 15428
rect 2370 15260 2380 15316
rect 2436 15260 2940 15316
rect 2996 15260 5068 15316
rect 5124 15260 5134 15316
rect 6962 15260 6972 15316
rect 7028 15260 8540 15316
rect 8596 15260 8606 15316
rect 10322 15260 10332 15316
rect 10388 15260 12796 15316
rect 12852 15260 12862 15316
rect 19842 15260 19852 15316
rect 19908 15260 21644 15316
rect 21700 15260 21710 15316
rect 24546 15260 24556 15316
rect 24612 15260 25228 15316
rect 25284 15260 25294 15316
rect 25452 15204 25508 15484
rect 25890 15372 25900 15428
rect 25956 15372 26460 15428
rect 26516 15372 27132 15428
rect 27188 15372 27198 15428
rect 27458 15372 27468 15428
rect 27524 15372 29260 15428
rect 29316 15372 29326 15428
rect 26338 15260 26348 15316
rect 26404 15260 26796 15316
rect 26852 15260 26862 15316
rect 28354 15260 28364 15316
rect 28420 15260 28430 15316
rect 31266 15260 31276 15316
rect 31332 15260 34524 15316
rect 34580 15260 34590 15316
rect 28364 15204 28420 15260
rect 15586 15148 15596 15204
rect 15652 15148 21980 15204
rect 22036 15148 22046 15204
rect 23090 15148 23100 15204
rect 23156 15148 25452 15204
rect 25508 15148 25518 15204
rect 26646 15148 26684 15204
rect 26740 15148 28420 15204
rect 34178 15148 34188 15204
rect 34244 15148 35084 15204
rect 35140 15148 35420 15204
rect 35476 15148 35486 15204
rect 25190 15036 25228 15092
rect 25284 15036 25294 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 15922 14700 15932 14756
rect 15988 14700 16828 14756
rect 16884 14700 16894 14756
rect 24658 14700 24668 14756
rect 24724 14700 26124 14756
rect 26180 14700 26348 14756
rect 26404 14700 26414 14756
rect 26786 14700 26796 14756
rect 26852 14700 31500 14756
rect 31556 14700 31566 14756
rect 9874 14588 9884 14644
rect 9940 14588 10892 14644
rect 10948 14588 11900 14644
rect 11956 14588 11966 14644
rect 20066 14588 20076 14644
rect 20132 14588 22092 14644
rect 22148 14588 22158 14644
rect 22866 14588 22876 14644
rect 22932 14588 26124 14644
rect 26180 14588 26190 14644
rect 5058 14476 5068 14532
rect 5124 14476 5964 14532
rect 6020 14476 7084 14532
rect 7140 14476 8204 14532
rect 8260 14476 8270 14532
rect 12898 14476 12908 14532
rect 12964 14476 13804 14532
rect 13860 14476 18508 14532
rect 18564 14476 18574 14532
rect 21298 14476 21308 14532
rect 21364 14476 24220 14532
rect 24276 14476 27692 14532
rect 27748 14476 27758 14532
rect 4162 14364 4172 14420
rect 4228 14364 6188 14420
rect 6244 14364 6254 14420
rect 8978 14364 8988 14420
rect 9044 14364 10220 14420
rect 10276 14364 10286 14420
rect 14130 14364 14140 14420
rect 14196 14364 14924 14420
rect 14980 14364 14990 14420
rect 11218 14252 11228 14308
rect 11284 14252 13580 14308
rect 13636 14252 13646 14308
rect 30594 14252 30604 14308
rect 30660 14252 31612 14308
rect 31668 14252 31678 14308
rect 24210 14140 24220 14196
rect 24276 14140 25116 14196
rect 25172 14140 25182 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 12786 14028 12796 14084
rect 12852 14028 13468 14084
rect 13524 14028 13534 14084
rect 25554 14028 25564 14084
rect 25620 14028 28364 14084
rect 28420 14028 34972 14084
rect 35028 14028 35756 14084
rect 35812 14028 35822 14084
rect 8372 13916 9100 13972
rect 9156 13916 11788 13972
rect 11844 13916 11854 13972
rect 13122 13916 13132 13972
rect 13188 13916 13804 13972
rect 13860 13916 13870 13972
rect 25302 13916 25340 13972
rect 25396 13916 25406 13972
rect 27122 13916 27132 13972
rect 27188 13916 27244 13972
rect 27300 13916 27310 13972
rect 2482 13804 2492 13860
rect 2548 13804 3724 13860
rect 3780 13804 3790 13860
rect 8372 13636 8428 13916
rect 12226 13804 12236 13860
rect 12292 13804 13916 13860
rect 13972 13804 14476 13860
rect 14532 13804 14542 13860
rect 23426 13804 23436 13860
rect 23492 13804 24108 13860
rect 24164 13804 24174 13860
rect 26852 13804 33236 13860
rect 26786 13692 26796 13748
rect 26852 13692 26908 13804
rect 33180 13748 33236 13804
rect 27122 13692 27132 13748
rect 27188 13692 27198 13748
rect 27906 13692 27916 13748
rect 27972 13692 33012 13748
rect 33170 13692 33180 13748
rect 33236 13692 33246 13748
rect 27132 13636 27188 13692
rect 32956 13636 33012 13692
rect 5282 13580 5292 13636
rect 5348 13580 5358 13636
rect 8194 13580 8204 13636
rect 8260 13580 8428 13636
rect 8866 13580 8876 13636
rect 8932 13580 10668 13636
rect 10724 13580 10734 13636
rect 16594 13580 16604 13636
rect 16660 13580 18284 13636
rect 18340 13580 18350 13636
rect 19618 13580 19628 13636
rect 19684 13580 21420 13636
rect 21476 13580 22316 13636
rect 22372 13580 24444 13636
rect 24500 13580 24510 13636
rect 26012 13580 27188 13636
rect 27458 13580 27468 13636
rect 27524 13580 29932 13636
rect 29988 13580 29998 13636
rect 32956 13580 35084 13636
rect 35140 13580 35150 13636
rect 5292 13524 5348 13580
rect 8876 13524 8932 13580
rect 5292 13468 8932 13524
rect 11330 13468 11340 13524
rect 11396 13468 14140 13524
rect 14196 13468 14206 13524
rect 15092 13468 21196 13524
rect 21252 13468 21868 13524
rect 21924 13468 21934 13524
rect 24098 13468 24108 13524
rect 24164 13468 25564 13524
rect 25620 13468 25630 13524
rect 15092 13412 15148 13468
rect 26012 13412 26068 13580
rect 26338 13468 26348 13524
rect 26404 13468 26908 13524
rect 26964 13468 26974 13524
rect 28466 13468 28476 13524
rect 28532 13468 29596 13524
rect 29652 13468 31276 13524
rect 31332 13468 31342 13524
rect 8530 13356 8540 13412
rect 8596 13356 9996 13412
rect 10052 13356 12460 13412
rect 12516 13356 15148 13412
rect 24434 13356 24444 13412
rect 24500 13356 26012 13412
rect 26068 13356 26078 13412
rect 27346 13356 27356 13412
rect 27412 13356 27524 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 8194 13244 8204 13300
rect 8260 13244 9772 13300
rect 9828 13244 9838 13300
rect 21858 13244 21868 13300
rect 21924 13244 23548 13300
rect 23604 13244 23614 13300
rect 3266 13132 3276 13188
rect 3332 13132 5740 13188
rect 5796 13132 5806 13188
rect 11666 13132 11676 13188
rect 11732 13132 12572 13188
rect 12628 13132 12638 13188
rect 20850 13132 20860 13188
rect 20916 13132 22092 13188
rect 22148 13132 22158 13188
rect 22306 13132 22316 13188
rect 22372 13132 26908 13188
rect 26964 13132 27244 13188
rect 27300 13132 27310 13188
rect 27468 13076 27524 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 6402 13020 6412 13076
rect 6468 13020 11228 13076
rect 11284 13020 11294 13076
rect 17154 13020 17164 13076
rect 17220 13020 24444 13076
rect 24500 13020 24510 13076
rect 25554 13020 25564 13076
rect 25620 13020 26236 13076
rect 26292 13020 26302 13076
rect 26852 13020 29764 13076
rect 22764 12964 22820 13020
rect 26852 12964 26908 13020
rect 29708 12964 29764 13020
rect 4946 12908 4956 12964
rect 5012 12908 6076 12964
rect 6132 12908 12012 12964
rect 12068 12908 12078 12964
rect 13906 12908 13916 12964
rect 13972 12908 14700 12964
rect 14756 12908 14766 12964
rect 22754 12908 22764 12964
rect 22820 12908 22830 12964
rect 24322 12908 24332 12964
rect 24388 12908 25116 12964
rect 25172 12908 25182 12964
rect 25666 12908 25676 12964
rect 25732 12908 26908 12964
rect 27542 12908 27580 12964
rect 27636 12908 27646 12964
rect 27990 12908 28028 12964
rect 28084 12908 28094 12964
rect 29362 12908 29372 12964
rect 29428 12908 29438 12964
rect 29698 12908 29708 12964
rect 29764 12908 29774 12964
rect 29372 12852 29428 12908
rect 12898 12796 12908 12852
rect 12964 12796 14140 12852
rect 14196 12796 14206 12852
rect 22978 12796 22988 12852
rect 23044 12796 25004 12852
rect 25060 12796 25070 12852
rect 25330 12796 25340 12852
rect 25396 12796 29428 12852
rect 10882 12684 10892 12740
rect 10948 12684 13580 12740
rect 13636 12684 13646 12740
rect 18610 12684 18620 12740
rect 18676 12684 19404 12740
rect 19460 12684 26124 12740
rect 26180 12684 26190 12740
rect 4610 12572 4620 12628
rect 4676 12572 5404 12628
rect 5460 12572 11340 12628
rect 11396 12572 11406 12628
rect 21970 12572 21980 12628
rect 22036 12572 23772 12628
rect 23828 12572 27020 12628
rect 27076 12572 27086 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 16370 12460 16380 12516
rect 16436 12460 17388 12516
rect 17444 12460 17454 12516
rect 4050 12348 4060 12404
rect 4116 12348 5068 12404
rect 5124 12348 5134 12404
rect 23426 12348 23436 12404
rect 23492 12348 23884 12404
rect 23940 12348 23950 12404
rect 29922 12348 29932 12404
rect 29988 12348 30716 12404
rect 30772 12348 30782 12404
rect 6066 12236 6076 12292
rect 6132 12236 7196 12292
rect 7252 12236 8316 12292
rect 8372 12236 8382 12292
rect 10210 12124 10220 12180
rect 10276 12124 12348 12180
rect 12404 12124 12414 12180
rect 18386 12124 18396 12180
rect 18452 12124 20524 12180
rect 20580 12124 20590 12180
rect 24770 12124 24780 12180
rect 24836 12124 27020 12180
rect 27076 12124 27916 12180
rect 27972 12124 27982 12180
rect 37090 12124 37100 12180
rect 37156 12124 39116 12180
rect 39172 12124 39182 12180
rect 12450 12012 12460 12068
rect 12516 12012 12684 12068
rect 12740 12012 12750 12068
rect 26310 12012 26348 12068
rect 26404 12012 26908 12068
rect 26964 12012 26974 12068
rect 34290 12012 34300 12068
rect 34356 12012 35980 12068
rect 36036 12012 36046 12068
rect 19282 11900 19292 11956
rect 19348 11900 20076 11956
rect 20132 11900 20748 11956
rect 20804 11900 20814 11956
rect 25330 11900 25340 11956
rect 25396 11900 26460 11956
rect 26516 11900 29596 11956
rect 29652 11900 33964 11956
rect 34020 11900 34030 11956
rect 12450 11788 12460 11844
rect 12516 11788 13916 11844
rect 13972 11788 13982 11844
rect 20290 11788 20300 11844
rect 20356 11788 21924 11844
rect 26338 11788 26348 11844
rect 26404 11788 26414 11844
rect 35970 11788 35980 11844
rect 36036 11788 38444 11844
rect 38500 11788 38510 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 21868 11732 21924 11788
rect 21868 11676 22092 11732
rect 22148 11676 23996 11732
rect 24052 11676 24062 11732
rect 26348 11620 26404 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 31490 11676 31500 11732
rect 31556 11676 33628 11732
rect 33684 11676 34524 11732
rect 34580 11676 34590 11732
rect 7410 11564 7420 11620
rect 7476 11564 8540 11620
rect 8596 11564 8606 11620
rect 14802 11564 14812 11620
rect 14868 11564 15372 11620
rect 15428 11564 15438 11620
rect 23492 11564 24332 11620
rect 24388 11564 26404 11620
rect 30370 11564 30380 11620
rect 30436 11564 30716 11620
rect 30772 11564 35532 11620
rect 35588 11564 35598 11620
rect 1810 11452 1820 11508
rect 1876 11452 4844 11508
rect 4900 11452 5628 11508
rect 5684 11452 6076 11508
rect 6132 11452 8876 11508
rect 8932 11452 9548 11508
rect 9604 11452 9614 11508
rect 15698 11452 15708 11508
rect 15764 11452 16604 11508
rect 16660 11452 17276 11508
rect 17332 11452 17836 11508
rect 17892 11452 19964 11508
rect 20020 11452 20030 11508
rect 23426 11452 23436 11508
rect 23492 11452 23548 11564
rect 24546 11452 24556 11508
rect 24612 11452 30604 11508
rect 30660 11452 30670 11508
rect 14578 11340 14588 11396
rect 14644 11340 15484 11396
rect 15540 11340 15550 11396
rect 25442 11340 25452 11396
rect 25508 11340 26684 11396
rect 26740 11340 26750 11396
rect 27458 11340 27468 11396
rect 27524 11340 33852 11396
rect 33908 11340 35756 11396
rect 35812 11340 35822 11396
rect 8530 11228 8540 11284
rect 8596 11228 14028 11284
rect 14084 11228 14094 11284
rect 20626 11228 20636 11284
rect 20692 11228 22876 11284
rect 22932 11228 22942 11284
rect 29250 11228 29260 11284
rect 29316 11228 30940 11284
rect 30996 11228 31006 11284
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 18946 10780 18956 10836
rect 19012 10780 20300 10836
rect 20356 10780 20366 10836
rect 24658 10780 24668 10836
rect 24724 10780 29596 10836
rect 29652 10780 29662 10836
rect 30258 10780 30268 10836
rect 30324 10780 31500 10836
rect 31556 10780 31566 10836
rect 12562 10668 12572 10724
rect 12628 10668 15372 10724
rect 15428 10668 15438 10724
rect 28242 10668 28252 10724
rect 28308 10668 30828 10724
rect 30884 10668 30894 10724
rect 27682 10444 27692 10500
rect 27748 10444 28588 10500
rect 28644 10444 28654 10500
rect 20066 10332 20076 10388
rect 20132 10332 21532 10388
rect 21588 10332 21598 10388
rect 19058 10220 19068 10276
rect 19124 10220 25228 10276
rect 25284 10220 25294 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 20178 9996 20188 10052
rect 20244 9996 23324 10052
rect 23380 9996 24556 10052
rect 24612 9996 24622 10052
rect 26002 9996 26012 10052
rect 26068 9996 26796 10052
rect 26852 9996 26862 10052
rect 15026 9884 15036 9940
rect 15092 9884 16380 9940
rect 16436 9884 16446 9940
rect 16930 9884 16940 9940
rect 16996 9884 24668 9940
rect 24724 9884 25004 9940
rect 25060 9884 25070 9940
rect 19618 9772 19628 9828
rect 19684 9772 20412 9828
rect 20468 9772 20478 9828
rect 22306 9772 22316 9828
rect 22372 9772 24332 9828
rect 24388 9772 24398 9828
rect 6626 9660 6636 9716
rect 6692 9660 7308 9716
rect 7364 9660 7374 9716
rect 8978 9660 8988 9716
rect 9044 9660 11900 9716
rect 11956 9660 11966 9716
rect 25218 9548 25228 9604
rect 25284 9548 25564 9604
rect 25620 9548 25630 9604
rect 30146 9548 30156 9604
rect 30212 9548 31388 9604
rect 31444 9548 31454 9604
rect 26226 9436 26236 9492
rect 26292 9436 26572 9492
rect 26628 9436 26638 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 15138 9324 15148 9380
rect 15204 9324 15484 9380
rect 15540 9324 15550 9380
rect 26002 9212 26012 9268
rect 26068 9212 29148 9268
rect 29204 9212 29214 9268
rect 25890 9100 25900 9156
rect 25956 9100 25966 9156
rect 26450 9100 26460 9156
rect 26516 9100 27580 9156
rect 27636 9100 27646 9156
rect 25900 9044 25956 9100
rect 24546 8988 24556 9044
rect 24612 8988 25228 9044
rect 25284 8988 25294 9044
rect 25900 8988 26460 9044
rect 26516 8988 26526 9044
rect 26674 8988 26684 9044
rect 26740 8988 27804 9044
rect 27860 8988 27870 9044
rect 7634 8876 7644 8932
rect 7700 8876 8988 8932
rect 9044 8876 9054 8932
rect 19282 8876 19292 8932
rect 19348 8876 20076 8932
rect 20132 8876 21308 8932
rect 21364 8876 22316 8932
rect 22372 8876 22382 8932
rect 26852 8820 26908 8932
rect 26964 8876 26974 8932
rect 14690 8764 14700 8820
rect 14756 8764 16268 8820
rect 16324 8764 18060 8820
rect 18116 8764 18732 8820
rect 18788 8764 18798 8820
rect 20402 8764 20412 8820
rect 20468 8764 21980 8820
rect 22036 8764 22046 8820
rect 24322 8764 24332 8820
rect 24388 8764 26908 8820
rect 12898 8652 12908 8708
rect 12964 8652 13692 8708
rect 13748 8652 25564 8708
rect 25620 8652 25630 8708
rect 26422 8652 26460 8708
rect 26516 8652 26526 8708
rect 26674 8652 26684 8708
rect 26740 8652 26778 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 26852 8484 26908 8764
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 21746 8428 21756 8484
rect 21812 8428 23772 8484
rect 23828 8428 23838 8484
rect 25330 8428 25340 8484
rect 25396 8428 25406 8484
rect 26562 8428 26572 8484
rect 26628 8428 26908 8484
rect 9762 8316 9772 8372
rect 9828 8316 13580 8372
rect 13636 8316 13646 8372
rect 11890 8204 11900 8260
rect 11956 8204 12572 8260
rect 12628 8204 13132 8260
rect 13188 8204 17836 8260
rect 17892 8204 17902 8260
rect 18274 8204 18284 8260
rect 18340 8204 19180 8260
rect 19236 8204 19246 8260
rect 22876 8148 22932 8428
rect 25340 8372 25396 8428
rect 23650 8316 23660 8372
rect 23716 8316 27132 8372
rect 27188 8316 27198 8372
rect 27906 8316 27916 8372
rect 27972 8316 28588 8372
rect 28644 8316 28654 8372
rect 31266 8316 31276 8372
rect 31332 8316 32844 8372
rect 32900 8316 32910 8372
rect 23986 8204 23996 8260
rect 24052 8204 24668 8260
rect 24724 8204 24734 8260
rect 12226 8092 12236 8148
rect 12292 8092 14140 8148
rect 14196 8092 14206 8148
rect 14802 8092 14812 8148
rect 14868 8092 17724 8148
rect 17780 8092 17790 8148
rect 22866 8092 22876 8148
rect 22932 8092 22942 8148
rect 23874 8092 23884 8148
rect 23940 8092 24444 8148
rect 24500 8092 24510 8148
rect 18498 7980 18508 8036
rect 18564 7980 19180 8036
rect 19236 7980 19246 8036
rect 20066 7980 20076 8036
rect 20132 7980 22148 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 22092 7700 22148 7980
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 22306 7756 22316 7812
rect 22372 7756 24220 7812
rect 24276 7756 24286 7812
rect 19170 7644 19180 7700
rect 19236 7644 21868 7700
rect 21924 7644 21934 7700
rect 22092 7644 23996 7700
rect 24052 7644 24668 7700
rect 24724 7644 24734 7700
rect 12898 7532 12908 7588
rect 12964 7532 13356 7588
rect 13412 7532 13916 7588
rect 13972 7532 13982 7588
rect 14690 7532 14700 7588
rect 14756 7532 18508 7588
rect 18564 7532 18574 7588
rect 13234 7420 13244 7476
rect 13300 7420 14812 7476
rect 14868 7420 14878 7476
rect 16818 7420 16828 7476
rect 16884 7420 17500 7476
rect 17556 7420 17566 7476
rect 17826 7420 17836 7476
rect 17892 7420 19404 7476
rect 19460 7420 19470 7476
rect 11442 7196 11452 7252
rect 11508 7196 12236 7252
rect 12292 7196 12302 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 23090 6860 23100 6916
rect 23156 6860 23548 6916
rect 23604 6860 23614 6916
rect 21858 6748 21868 6804
rect 21924 6748 22764 6804
rect 22820 6748 22830 6804
rect 24210 6748 24220 6804
rect 24276 6748 24892 6804
rect 24948 6748 24958 6804
rect 10098 6636 10108 6692
rect 10164 6636 12236 6692
rect 12292 6636 12684 6692
rect 12740 6636 12750 6692
rect 15698 6636 15708 6692
rect 15764 6636 16604 6692
rect 16660 6636 18956 6692
rect 19012 6636 19628 6692
rect 19684 6636 20300 6692
rect 20356 6636 20366 6692
rect 23986 6636 23996 6692
rect 24052 6636 26124 6692
rect 26180 6636 26190 6692
rect 15026 6524 15036 6580
rect 15092 6524 15260 6580
rect 15316 6524 15326 6580
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 22642 6188 22652 6244
rect 22708 6188 23884 6244
rect 23940 6188 24332 6244
rect 24388 6188 24398 6244
rect 16034 5964 16044 6020
rect 16100 5964 18508 6020
rect 18564 5964 19404 6020
rect 19460 5964 19470 6020
rect 22642 5964 22652 6020
rect 22708 5964 24220 6020
rect 24276 5964 24286 6020
rect 16482 5852 16492 5908
rect 16548 5852 17612 5908
rect 17668 5852 17678 5908
rect 26226 5740 26236 5796
rect 26292 5740 27020 5796
rect 27076 5740 28252 5796
rect 28308 5740 28318 5796
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 21522 5292 21532 5348
rect 21588 5292 23212 5348
rect 23268 5292 23278 5348
rect 19842 5180 19852 5236
rect 19908 5180 20860 5236
rect 20916 5180 22092 5236
rect 22148 5180 23492 5236
rect 21746 5068 21756 5124
rect 21812 5068 22876 5124
rect 22932 5068 22942 5124
rect 23436 5012 23492 5180
rect 23436 4956 24220 5012
rect 24276 4956 25340 5012
rect 25396 4956 25406 5012
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 25666 4508 25676 4564
rect 25732 4508 26684 4564
rect 26740 4508 26750 4564
rect 27906 4172 27916 4228
rect 27972 4172 29596 4228
rect 29652 4172 29662 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 39228 53340 39284 53396
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 35644 52780 35700 52836
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 35644 51884 35700 51940
rect 38780 51772 38836 51828
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 42140 51212 42196 51268
rect 38780 51100 38836 51156
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 39228 50652 39284 50708
rect 42140 50540 42196 50596
rect 22652 50428 22708 50484
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 26908 49196 26964 49252
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 26012 48524 26068 48580
rect 16044 48188 16100 48244
rect 22764 48076 22820 48132
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 27356 47740 27412 47796
rect 26012 47292 26068 47348
rect 15036 47180 15092 47236
rect 16044 47180 16100 47236
rect 21420 47068 21476 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 24892 46172 24948 46228
rect 19068 46060 19124 46116
rect 19404 45948 19460 46004
rect 19404 45500 19460 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 39564 45276 39620 45332
rect 17388 44716 17444 44772
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 45836 44044 45892 44100
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 27356 43932 27412 43988
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 39564 43708 39620 43764
rect 18620 43260 18676 43316
rect 17276 43148 17332 43204
rect 18844 43148 18900 43204
rect 23548 43148 23604 43204
rect 24892 43148 24948 43204
rect 51324 43148 51380 43204
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 45276 42924 45332 42980
rect 17276 42588 17332 42644
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 18844 42252 18900 42308
rect 19628 42252 19684 42308
rect 19068 42028 19124 42084
rect 22764 41804 22820 41860
rect 23884 41580 23940 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 16492 41356 16548 41412
rect 22652 41356 22708 41412
rect 26908 41356 26964 41412
rect 17388 41244 17444 41300
rect 15372 41132 15428 41188
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 18396 40572 18452 40628
rect 19628 40572 19684 40628
rect 51324 40348 51380 40404
rect 18620 40124 18676 40180
rect 19516 40124 19572 40180
rect 23884 40124 23940 40180
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 15036 39788 15092 39844
rect 49644 39788 49700 39844
rect 23548 39676 23604 39732
rect 49532 39676 49588 39732
rect 19628 39452 19684 39508
rect 49644 39452 49700 39508
rect 21420 39340 21476 39396
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 17388 39004 17444 39060
rect 17948 39004 18004 39060
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 15372 38892 15428 38948
rect 49532 38892 49588 38948
rect 16492 38556 16548 38612
rect 18396 38556 18452 38612
rect 17948 38444 18004 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 38220 38220 38276 38276
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 45164 37884 45220 37940
rect 50316 37772 50372 37828
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 38220 37548 38276 37604
rect 19628 37100 19684 37156
rect 45836 37212 45892 37268
rect 50316 37212 50372 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 45276 36876 45332 36932
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 19516 35980 19572 36036
rect 23436 35868 23492 35924
rect 45164 35644 45220 35700
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 23436 33180 23492 33236
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 39116 32620 39172 32676
rect 46956 32620 47012 32676
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 46732 32060 46788 32116
rect 50316 31836 50372 31892
rect 39116 31500 39172 31556
rect 46844 31388 46900 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 50316 30940 50372 30996
rect 46732 30828 46788 30884
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 46844 30268 46900 30324
rect 47740 30268 47796 30324
rect 49084 30268 49140 30324
rect 48972 30156 49028 30212
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 45836 29708 45892 29764
rect 39116 29484 39172 29540
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 42476 28364 42532 28420
rect 45836 28364 45892 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 46956 27916 47012 27972
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 48188 27356 48244 27412
rect 33740 27244 33796 27300
rect 33740 26796 33796 26852
rect 38668 26796 38724 26852
rect 46844 26796 46900 26852
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 42476 26572 42532 26628
rect 50988 26236 51044 26292
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 38668 25340 38724 25396
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 50316 24668 50372 24724
rect 50988 24668 51044 24724
rect 38668 24556 38724 24612
rect 39116 24332 39172 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 48300 23772 48356 23828
rect 48972 23772 49028 23828
rect 49308 23772 49364 23828
rect 48188 23548 48244 23604
rect 49308 23548 49364 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 50092 23436 50148 23492
rect 49084 23100 49140 23156
rect 50316 22988 50372 23044
rect 50092 22876 50148 22932
rect 49084 22764 49140 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 23212 21644 23268 21700
rect 47740 21644 47796 21700
rect 26124 21308 26180 21364
rect 48300 21196 48356 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 22204 21084 22260 21140
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 23212 20188 23268 20244
rect 22428 20076 22484 20132
rect 25228 20076 25284 20132
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 22204 19516 22260 19572
rect 22428 19068 22484 19124
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 28028 18396 28084 18452
rect 26348 18172 26404 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 15148 17836 15204 17892
rect 25788 17612 25844 17668
rect 15148 17500 15204 17556
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 26908 17164 26964 17220
rect 27244 17164 27300 17220
rect 25340 17052 25396 17108
rect 27468 17052 27524 17108
rect 25676 16828 25732 16884
rect 26908 16828 26964 16884
rect 27580 16828 27636 16884
rect 25676 16604 25732 16660
rect 27468 16604 27524 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 25788 16044 25844 16100
rect 26684 16044 26740 16100
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 26684 15148 26740 15204
rect 25228 15036 25284 15092
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 26124 14700 26180 14756
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 25340 13916 25396 13972
rect 27244 13916 27300 13972
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 26908 13132 26964 13188
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 27580 12908 27636 12964
rect 28028 12908 28084 12964
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 26348 12012 26404 12068
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 26460 9100 26516 9156
rect 26684 8988 26740 9044
rect 26460 8652 26516 8708
rect 26684 8652 26740 8708
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 39228 53396 39284 53406
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35644 52836 35700 52846
rect 35644 51940 35700 52780
rect 35644 51874 35700 51884
rect 38780 51828 38836 51838
rect 38780 51156 38836 51772
rect 38780 51090 38836 51100
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 16044 48244 16100 48254
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 15036 47236 15092 47246
rect 15036 39844 15092 47180
rect 16044 47236 16100 48188
rect 16044 47170 16100 47180
rect 19808 47068 20128 48580
rect 22652 50484 22708 50494
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19068 46116 19124 46126
rect 17388 44772 17444 44782
rect 17276 43204 17332 43214
rect 17276 42644 17332 43148
rect 17276 42578 17332 42588
rect 16492 41412 16548 41422
rect 15036 39778 15092 39788
rect 15372 41188 15428 41198
rect 15372 38948 15428 41132
rect 15372 38882 15428 38892
rect 16492 38612 16548 41356
rect 17388 41300 17444 44716
rect 17388 39060 17444 41244
rect 18620 43316 18676 43326
rect 18396 40628 18452 40638
rect 17388 38994 17444 39004
rect 17948 39060 18004 39070
rect 16492 38546 16548 38556
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 17948 38500 18004 39004
rect 18396 38612 18452 40572
rect 18620 40180 18676 43260
rect 18844 43204 18900 43214
rect 18844 42308 18900 43148
rect 18844 42242 18900 42252
rect 19068 42084 19124 46060
rect 19404 46004 19460 46014
rect 19404 45556 19460 45948
rect 19404 45490 19460 45500
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19068 42018 19124 42028
rect 19628 42308 19684 42318
rect 19628 40628 19684 42252
rect 19628 40562 19684 40572
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 18620 40114 18676 40124
rect 19516 40180 19572 40190
rect 18396 38546 18452 38556
rect 17948 38434 18004 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 19516 36036 19572 40124
rect 19628 39508 19684 39518
rect 19628 37156 19684 39452
rect 19628 37090 19684 37100
rect 19808 39228 20128 40740
rect 21420 47124 21476 47134
rect 21420 39396 21476 47068
rect 22652 41412 22708 50428
rect 35168 49420 35488 50932
rect 39228 50708 39284 53340
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 39228 50642 39284 50652
rect 42140 51268 42196 51278
rect 42140 50596 42196 51212
rect 42140 50530 42196 50540
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 26908 49252 26964 49262
rect 26012 48580 26068 48590
rect 22764 48132 22820 48142
rect 22764 41860 22820 48076
rect 26012 47348 26068 48524
rect 26012 47282 26068 47292
rect 24892 46228 24948 46238
rect 22764 41794 22820 41804
rect 23548 43204 23604 43214
rect 22652 41346 22708 41356
rect 23548 39732 23604 43148
rect 24892 43204 24948 46172
rect 24892 43138 24948 43148
rect 23884 41636 23940 41646
rect 23884 40180 23940 41580
rect 26908 41412 26964 49196
rect 35168 47852 35488 49364
rect 27356 47796 27412 47806
rect 27356 43988 27412 47740
rect 27356 43922 27412 43932
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 26908 41346 26964 41356
rect 35168 43148 35488 44660
rect 39564 45332 39620 45342
rect 39564 43764 39620 45276
rect 39564 43698 39620 43708
rect 45836 44100 45892 44110
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 23884 40114 23940 40124
rect 23548 39666 23604 39676
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 21420 39330 21476 39340
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19516 35970 19572 35980
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 19808 34524 20128 36036
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 45276 42980 45332 42990
rect 38220 38276 38276 38286
rect 38220 37604 38276 38220
rect 38220 37538 38276 37548
rect 45164 37940 45220 37950
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 23436 35924 23492 35934
rect 23436 33236 23492 35868
rect 23436 33170 23492 33180
rect 35168 35308 35488 36820
rect 45164 35700 45220 37884
rect 45276 36932 45332 42924
rect 45836 37268 45892 44044
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 49644 39844 49700 39854
rect 49532 39732 49588 39742
rect 49532 38948 49588 39676
rect 49644 39508 49700 39788
rect 49644 39442 49700 39452
rect 49532 38882 49588 38892
rect 50528 39228 50848 40740
rect 51324 43204 51380 43214
rect 51324 40404 51380 43148
rect 51324 40338 51380 40348
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 45836 37202 45892 37212
rect 50316 37828 50372 37838
rect 50316 37268 50372 37772
rect 45276 36866 45332 36876
rect 45164 35634 45220 35644
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 33740 27300 33796 27310
rect 33740 26852 33796 27244
rect 33740 26786 33796 26796
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 35168 25900 35488 27412
rect 39116 32676 39172 32686
rect 39116 31556 39172 32620
rect 46956 32676 47012 32686
rect 39116 29540 39172 31500
rect 46732 32116 46788 32126
rect 46732 30884 46788 32060
rect 46732 30818 46788 30828
rect 46844 31444 46900 31454
rect 46844 30324 46900 31388
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 38668 26852 38724 26862
rect 38668 25396 38724 26796
rect 38668 24612 38724 25340
rect 38668 24546 38724 24556
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 39116 24388 39172 29484
rect 45836 29764 45892 29774
rect 42476 28420 42532 28430
rect 42476 26628 42532 28364
rect 45836 28420 45892 29708
rect 45836 28354 45892 28364
rect 46844 26852 46900 30268
rect 46956 27972 47012 32620
rect 50316 31892 50372 37212
rect 50316 30996 50372 31836
rect 50316 30930 50372 30940
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 46956 27906 47012 27916
rect 47740 30324 47796 30334
rect 46844 26786 46900 26796
rect 42476 26562 42532 26572
rect 39116 24322 39172 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 23212 21700 23268 21710
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 22204 21140 22260 21150
rect 22204 19572 22260 21084
rect 23212 20244 23268 21644
rect 23212 20178 23268 20188
rect 26124 21364 26180 21374
rect 22204 19506 22260 19516
rect 22428 20132 22484 20142
rect 22428 19124 22484 20076
rect 22428 19058 22484 19068
rect 25228 20132 25284 20142
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 15148 17892 15204 17902
rect 15148 17556 15204 17836
rect 15148 17490 15204 17500
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 25228 15092 25284 20076
rect 25788 17668 25844 17678
rect 25228 15026 25284 15036
rect 25340 17108 25396 17118
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 25340 13972 25396 17052
rect 25676 16884 25732 16894
rect 25676 16660 25732 16828
rect 25676 16594 25732 16604
rect 25788 16100 25844 17612
rect 25788 16034 25844 16044
rect 26124 14756 26180 21308
rect 35168 21196 35488 22708
rect 47740 21700 47796 30268
rect 49084 30324 49140 30334
rect 48972 30212 49028 30222
rect 48188 27412 48244 27422
rect 48188 23604 48244 27356
rect 48188 23538 48244 23548
rect 48300 23828 48356 23838
rect 47740 21634 47796 21644
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 48300 21252 48356 23772
rect 48972 23828 49028 30156
rect 48972 23762 49028 23772
rect 49084 23156 49140 30268
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50316 24724 50372 24734
rect 49308 23828 49364 23838
rect 49308 23604 49364 23772
rect 49308 23538 49364 23548
rect 49084 22820 49140 23100
rect 50092 23492 50148 23502
rect 50092 22932 50148 23436
rect 50316 23044 50372 24668
rect 50316 22978 50372 22988
rect 50528 23548 50848 25060
rect 50988 26292 51044 26302
rect 50988 24724 51044 26236
rect 50988 24658 51044 24668
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50092 22866 50148 22876
rect 49084 22754 49140 22764
rect 48300 21186 48356 21196
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 28028 18452 28084 18462
rect 26124 14690 26180 14700
rect 26348 18228 26404 18238
rect 25340 13906 25396 13916
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 26348 12068 26404 18172
rect 26908 17220 26964 17230
rect 26908 16884 26964 17164
rect 26684 16100 26740 16110
rect 26684 15204 26740 16044
rect 26684 15138 26740 15148
rect 26908 13188 26964 16828
rect 27244 17220 27300 17230
rect 27244 13972 27300 17164
rect 27468 17108 27524 17118
rect 27468 16660 27524 17052
rect 27468 16594 27524 16604
rect 27580 16884 27636 16894
rect 27244 13906 27300 13916
rect 26908 13122 26964 13132
rect 27580 12964 27636 16828
rect 27580 12898 27636 12908
rect 28028 12964 28084 18396
rect 28028 12898 28084 12908
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 26348 12002 26404 12012
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 26460 9156 26516 9166
rect 26460 8708 26516 9100
rect 26460 8642 26516 8652
rect 26684 9044 26740 9054
rect 26684 8708 26740 8988
rect 26684 8642 26740 8652
rect 35168 8652 35488 10164
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1287_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42112 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1288_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1289_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 47600 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1290_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47376 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1291_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 50624 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1292_
timestamp 1698431365
transform -1 0 44128 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1293_
timestamp 1698431365
transform -1 0 48048 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1294_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45472 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1295_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46480 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1296_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 49616 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1297_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47936 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1298_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46368 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1299_
timestamp 1698431365
transform -1 0 43904 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1300_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42000 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1301_
timestamp 1698431365
transform 1 0 41776 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1302_
timestamp 1698431365
transform -1 0 41888 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1303_
timestamp 1698431365
transform -1 0 46928 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1304_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42784 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1305_
timestamp 1698431365
transform -1 0 39984 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1306_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41664 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1307_
timestamp 1698431365
transform 1 0 42336 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1308_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42560 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1309_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37072 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1310_
timestamp 1698431365
transform 1 0 44800 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1311_
timestamp 1698431365
transform 1 0 41664 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1312_
timestamp 1698431365
transform -1 0 41776 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1313_
timestamp 1698431365
transform 1 0 41104 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1314_
timestamp 1698431365
transform -1 0 41888 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1315_
timestamp 1698431365
transform -1 0 43456 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1316_
timestamp 1698431365
transform -1 0 40880 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1317_
timestamp 1698431365
transform -1 0 39312 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1318_
timestamp 1698431365
transform 1 0 39536 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1319_
timestamp 1698431365
transform 1 0 39760 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1320_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35280 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1321_
timestamp 1698431365
transform 1 0 37072 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1322_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40432 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1323_
timestamp 1698431365
transform -1 0 40320 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1324_
timestamp 1698431365
transform 1 0 37744 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1325_
timestamp 1698431365
transform 1 0 41888 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1326_
timestamp 1698431365
transform -1 0 41328 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1327_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform 1 0 43456 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1329_
timestamp 1698431365
transform 1 0 37632 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1330_
timestamp 1698431365
transform 1 0 39424 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1331_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39648 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1332_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38304 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1333_
timestamp 1698431365
transform -1 0 32480 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1334_
timestamp 1698431365
transform -1 0 38304 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1335_
timestamp 1698431365
transform -1 0 36400 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1336_
timestamp 1698431365
transform -1 0 35728 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1337_
timestamp 1698431365
transform -1 0 39424 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1338_
timestamp 1698431365
transform -1 0 38528 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1339_
timestamp 1698431365
transform -1 0 41440 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1340_
timestamp 1698431365
transform 1 0 34496 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1341_
timestamp 1698431365
transform -1 0 34720 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1342_
timestamp 1698431365
transform 1 0 35728 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1343_
timestamp 1698431365
transform 1 0 41888 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1344_
timestamp 1698431365
transform -1 0 36400 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1345_
timestamp 1698431365
transform 1 0 36624 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1346_
timestamp 1698431365
transform 1 0 35840 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1347_
timestamp 1698431365
transform -1 0 36176 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1348_
timestamp 1698431365
transform 1 0 12096 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1349_
timestamp 1698431365
transform 1 0 29344 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1350_
timestamp 1698431365
transform 1 0 31360 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1351_
timestamp 1698431365
transform -1 0 32704 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1352_
timestamp 1698431365
transform 1 0 12656 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1353_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1354_
timestamp 1698431365
transform 1 0 11648 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1355_
timestamp 1698431365
transform 1 0 13888 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1356_
timestamp 1698431365
transform -1 0 19264 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1357_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17136 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1358_
timestamp 1698431365
transform 1 0 11088 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1359_
timestamp 1698431365
transform -1 0 11536 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1360_
timestamp 1698431365
transform -1 0 15232 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1361_
timestamp 1698431365
transform 1 0 12432 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1362_
timestamp 1698431365
transform -1 0 11984 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1363_
timestamp 1698431365
transform -1 0 15344 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1364_
timestamp 1698431365
transform 1 0 14560 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1365_
timestamp 1698431365
transform 1 0 12656 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1366_
timestamp 1698431365
transform 1 0 12096 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1367_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1368_
timestamp 1698431365
transform -1 0 24192 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1369_
timestamp 1698431365
transform 1 0 20272 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1370_
timestamp 1698431365
transform 1 0 21056 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1371_
timestamp 1698431365
transform 1 0 18144 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1372_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19152 0 -1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1373_
timestamp 1698431365
transform -1 0 19936 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1374_
timestamp 1698431365
transform -1 0 18816 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1375_
timestamp 1698431365
transform 1 0 16128 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1376_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1377_
timestamp 1698431365
transform -1 0 18368 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1378_
timestamp 1698431365
transform -1 0 14672 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1379_
timestamp 1698431365
transform 1 0 11312 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1380_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16912 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1381_
timestamp 1698431365
transform -1 0 13104 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1382_
timestamp 1698431365
transform -1 0 18816 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1383_
timestamp 1698431365
transform -1 0 11648 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1384_
timestamp 1698431365
transform 1 0 10416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1385_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10864 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1386_
timestamp 1698431365
transform 1 0 11760 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1387_
timestamp 1698431365
transform 1 0 31696 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1388_
timestamp 1698431365
transform 1 0 30800 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1389_
timestamp 1698431365
transform -1 0 18144 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1390_
timestamp 1698431365
transform -1 0 18144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1391_
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1392_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18368 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1393_
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1394_
timestamp 1698431365
transform -1 0 22064 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1395_
timestamp 1698431365
transform -1 0 19264 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1396_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 -1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1397_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1398_
timestamp 1698431365
transform -1 0 27440 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1399_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26432 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1400_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1401_
timestamp 1698431365
transform -1 0 22624 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1402_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21056 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1403_
timestamp 1698431365
transform 1 0 21616 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1404_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26992 0 1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1405_
timestamp 1698431365
transform -1 0 18592 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1406_
timestamp 1698431365
transform -1 0 18592 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1407_
timestamp 1698431365
transform 1 0 16352 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1408_
timestamp 1698431365
transform -1 0 16352 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1409_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1410_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 29792
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1411_
timestamp 1698431365
transform -1 0 17920 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1412_
timestamp 1698431365
transform 1 0 17472 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1413_
timestamp 1698431365
transform 1 0 24864 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1414_
timestamp 1698431365
transform -1 0 17696 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1415_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24864 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1416_
timestamp 1698431365
transform 1 0 27104 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1417_
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1418_
timestamp 1698431365
transform -1 0 17920 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1419_
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1420_
timestamp 1698431365
transform 1 0 28336 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1421_
timestamp 1698431365
transform 1 0 25648 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1422_
timestamp 1698431365
transform -1 0 30352 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1423_
timestamp 1698431365
transform -1 0 17472 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1424_
timestamp 1698431365
transform 1 0 23072 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1425_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1426_
timestamp 1698431365
transform 1 0 16240 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1427_
timestamp 1698431365
transform 1 0 27664 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1428_
timestamp 1698431365
transform 1 0 34944 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1429_
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1430_
timestamp 1698431365
transform -1 0 25984 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1431_
timestamp 1698431365
transform 1 0 29120 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1432_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1433_
timestamp 1698431365
transform -1 0 16240 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1434_
timestamp 1698431365
transform 1 0 16688 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1435_
timestamp 1698431365
transform -1 0 28112 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1436_
timestamp 1698431365
transform -1 0 16912 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1437_
timestamp 1698431365
transform -1 0 27440 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1438_
timestamp 1698431365
transform 1 0 33600 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1439_
timestamp 1698431365
transform -1 0 29344 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1440_
timestamp 1698431365
transform 1 0 27440 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1441_
timestamp 1698431365
transform -1 0 28896 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1442_
timestamp 1698431365
transform -1 0 27664 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1443_
timestamp 1698431365
transform 1 0 23184 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1444_
timestamp 1698431365
transform 1 0 22736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1445_
timestamp 1698431365
transform 1 0 25984 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1446_
timestamp 1698431365
transform 1 0 24864 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1447_
timestamp 1698431365
transform 1 0 23744 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1448_
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1449_
timestamp 1698431365
transform -1 0 24864 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1450_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1451_
timestamp 1698431365
transform -1 0 14448 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1452_
timestamp 1698431365
transform -1 0 14672 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1453_
timestamp 1698431365
transform 1 0 13552 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1454_
timestamp 1698431365
transform 1 0 9520 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1455_
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1456_
timestamp 1698431365
transform -1 0 16688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1457_
timestamp 1698431365
transform -1 0 11984 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1458_
timestamp 1698431365
transform -1 0 10864 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1459_
timestamp 1698431365
transform 1 0 10864 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1698431365
transform -1 0 15792 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1461_
timestamp 1698431365
transform -1 0 13216 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1462_
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1463_
timestamp 1698431365
transform 1 0 6608 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1464_
timestamp 1698431365
transform -1 0 16912 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1465_
timestamp 1698431365
transform 1 0 8848 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1466_
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1467_
timestamp 1698431365
transform -1 0 15792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1468_
timestamp 1698431365
transform 1 0 12656 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1469_
timestamp 1698431365
transform 1 0 14112 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1470_
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1471_
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1472_
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1473_
timestamp 1698431365
transform 1 0 9744 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1474_
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1475_
timestamp 1698431365
transform -1 0 15680 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1476_
timestamp 1698431365
transform 1 0 13328 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1477_
timestamp 1698431365
transform -1 0 9520 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1478_
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1479_
timestamp 1698431365
transform 1 0 8512 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1480_
timestamp 1698431365
transform -1 0 9184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1481_
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1482_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1483_
timestamp 1698431365
transform 1 0 14336 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1484_
timestamp 1698431365
transform -1 0 17024 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1485_
timestamp 1698431365
transform 1 0 24864 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1486_
timestamp 1698431365
transform -1 0 26432 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1487_
timestamp 1698431365
transform -1 0 23856 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1488_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1489_
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1490_
timestamp 1698431365
transform -1 0 27888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1491_
timestamp 1698431365
transform 1 0 17808 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1492_
timestamp 1698431365
transform -1 0 28112 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1493_
timestamp 1698431365
transform 1 0 23744 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1494_
timestamp 1698431365
transform -1 0 27776 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1495_
timestamp 1698431365
transform -1 0 27664 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1496_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1497_
timestamp 1698431365
transform 1 0 26096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1498_
timestamp 1698431365
transform -1 0 28448 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1499_
timestamp 1698431365
transform 1 0 26656 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1500_
timestamp 1698431365
transform -1 0 26992 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1501_
timestamp 1698431365
transform -1 0 26544 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1502_
timestamp 1698431365
transform 1 0 31024 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1503_
timestamp 1698431365
transform -1 0 26656 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1504_
timestamp 1698431365
transform 1 0 20720 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1505_
timestamp 1698431365
transform -1 0 25536 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1506_
timestamp 1698431365
transform -1 0 26208 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1507_
timestamp 1698431365
transform 1 0 22960 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1508_
timestamp 1698431365
transform 1 0 21392 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1509_
timestamp 1698431365
transform 1 0 20384 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1510_
timestamp 1698431365
transform 1 0 21504 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1511_
timestamp 1698431365
transform -1 0 23744 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1512_
timestamp 1698431365
transform 1 0 23968 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1513_
timestamp 1698431365
transform 1 0 25536 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1514_
timestamp 1698431365
transform 1 0 11424 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1515_
timestamp 1698431365
transform 1 0 11088 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1516_
timestamp 1698431365
transform -1 0 15120 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1517_
timestamp 1698431365
transform 1 0 11424 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1518_
timestamp 1698431365
transform 1 0 10976 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1519_
timestamp 1698431365
transform 1 0 11984 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1520_
timestamp 1698431365
transform -1 0 15456 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1521_
timestamp 1698431365
transform 1 0 6160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1522_
timestamp 1698431365
transform 1 0 7280 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1523_
timestamp 1698431365
transform 1 0 7728 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1524_
timestamp 1698431365
transform -1 0 15008 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1525_
timestamp 1698431365
transform 1 0 15008 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1526_
timestamp 1698431365
transform 1 0 14672 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1527_
timestamp 1698431365
transform 1 0 8512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1528_
timestamp 1698431365
transform 1 0 7504 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1529_
timestamp 1698431365
transform -1 0 9296 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1530_
timestamp 1698431365
transform -1 0 15344 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1531_
timestamp 1698431365
transform 1 0 14336 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1532_
timestamp 1698431365
transform 1 0 7392 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1533_
timestamp 1698431365
transform 1 0 7392 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1534_
timestamp 1698431365
transform 1 0 8064 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1535_
timestamp 1698431365
transform -1 0 15120 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1536_
timestamp 1698431365
transform 1 0 15344 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1537_
timestamp 1698431365
transform -1 0 17024 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1538_
timestamp 1698431365
transform 1 0 24416 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1539_
timestamp 1698431365
transform -1 0 25536 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1540_
timestamp 1698431365
transform 1 0 24192 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1541_
timestamp 1698431365
transform -1 0 21616 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1542_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11984 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1543_
timestamp 1698431365
transform 1 0 12208 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1544_
timestamp 1698431365
transform -1 0 14224 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1545_
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1546_
timestamp 1698431365
transform 1 0 18368 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1547_
timestamp 1698431365
transform -1 0 19488 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1548_
timestamp 1698431365
transform 1 0 13552 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1549_
timestamp 1698431365
transform 1 0 15680 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1550_
timestamp 1698431365
transform 1 0 30576 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1551_
timestamp 1698431365
transform -1 0 30576 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1552_
timestamp 1698431365
transform 1 0 16128 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1553_
timestamp 1698431365
transform 1 0 21616 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1554_
timestamp 1698431365
transform 1 0 21280 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1555_
timestamp 1698431365
transform 1 0 44240 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1556_
timestamp 1698431365
transform 1 0 18368 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1557_
timestamp 1698431365
transform 1 0 22288 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1558_
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1559_
timestamp 1698431365
transform -1 0 23296 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1560_
timestamp 1698431365
transform -1 0 19264 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1561_
timestamp 1698431365
transform 1 0 19264 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1562_
timestamp 1698431365
transform 1 0 20048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1563_
timestamp 1698431365
transform -1 0 31584 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1564_
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1565_
timestamp 1698431365
transform 1 0 14448 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1566_
timestamp 1698431365
transform 1 0 11984 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1567_
timestamp 1698431365
transform 1 0 12880 0 -1 48608
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1568_
timestamp 1698431365
transform -1 0 15120 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1569_
timestamp 1698431365
transform 1 0 14896 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1570_
timestamp 1698431365
transform 1 0 15680 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1571_
timestamp 1698431365
transform 1 0 16016 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1572_
timestamp 1698431365
transform -1 0 31360 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1573_
timestamp 1698431365
transform -1 0 25088 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1574_
timestamp 1698431365
transform -1 0 25760 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1575_
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1576_
timestamp 1698431365
transform 1 0 19264 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1577_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1578_
timestamp 1698431365
transform 1 0 17024 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1579_
timestamp 1698431365
transform 1 0 16128 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1580_
timestamp 1698431365
transform 1 0 16352 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1581_
timestamp 1698431365
transform -1 0 19936 0 -1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1582_
timestamp 1698431365
transform -1 0 18144 0 1 54880
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1583_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18368 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1584_
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1585_
timestamp 1698431365
transform 1 0 18144 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1586_
timestamp 1698431365
transform -1 0 24192 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1587_
timestamp 1698431365
transform 1 0 15904 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1588_
timestamp 1698431365
transform 1 0 19712 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1589_
timestamp 1698431365
transform -1 0 20832 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1590_
timestamp 1698431365
transform -1 0 28112 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1591_
timestamp 1698431365
transform -1 0 16352 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1592_
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1593_
timestamp 1698431365
transform 1 0 15232 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1594_
timestamp 1698431365
transform 1 0 14896 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1595_
timestamp 1698431365
transform -1 0 14672 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1596_
timestamp 1698431365
transform 1 0 14336 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1597_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14784 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1598_
timestamp 1698431365
transform -1 0 15120 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1599_
timestamp 1698431365
transform -1 0 28784 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1600_
timestamp 1698431365
transform -1 0 15456 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1601_
timestamp 1698431365
transform -1 0 18592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1602_
timestamp 1698431365
transform -1 0 16352 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1603_
timestamp 1698431365
transform -1 0 14784 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1604_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14112 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1605_
timestamp 1698431365
transform -1 0 14000 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1606_
timestamp 1698431365
transform -1 0 44240 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1607_
timestamp 1698431365
transform 1 0 43232 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1608_
timestamp 1698431365
transform -1 0 43232 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1609_
timestamp 1698431365
transform -1 0 38640 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1610_
timestamp 1698431365
transform -1 0 36624 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1611_
timestamp 1698431365
transform 1 0 34048 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1612_
timestamp 1698431365
transform -1 0 36400 0 1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1613_
timestamp 1698431365
transform -1 0 35168 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1614_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34832 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1615_
timestamp 1698431365
transform -1 0 39760 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1616_
timestamp 1698431365
transform -1 0 41104 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1617_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 -1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1618_
timestamp 1698431365
transform 1 0 39312 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1619_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39312 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1620_
timestamp 1698431365
transform -1 0 35840 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1621_
timestamp 1698431365
transform -1 0 30576 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1622_
timestamp 1698431365
transform -1 0 35840 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1623_
timestamp 1698431365
transform 1 0 29008 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1624_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18032 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1625_
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1626_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19488 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1627_
timestamp 1698431365
transform 1 0 18592 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1628_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1629_
timestamp 1698431365
transform -1 0 20608 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1630_
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1631_
timestamp 1698431365
transform 1 0 16352 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1632_
timestamp 1698431365
transform -1 0 19264 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1633_
timestamp 1698431365
transform 1 0 19488 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1634_
timestamp 1698431365
transform 1 0 28112 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1635_
timestamp 1698431365
transform 1 0 28560 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1636_
timestamp 1698431365
transform -1 0 16016 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1637_
timestamp 1698431365
transform -1 0 24192 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1638_
timestamp 1698431365
transform 1 0 23296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1639_
timestamp 1698431365
transform -1 0 24864 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1640_
timestamp 1698431365
transform 1 0 22624 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1641_
timestamp 1698431365
transform 1 0 23408 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1642_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25424 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1643_
timestamp 1698431365
transform 1 0 19488 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1644_
timestamp 1698431365
transform -1 0 21952 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1645_
timestamp 1698431365
transform -1 0 19600 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1646_
timestamp 1698431365
transform 1 0 17360 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1647_
timestamp 1698431365
transform -1 0 19488 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1648_
timestamp 1698431365
transform 1 0 6384 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1649_
timestamp 1698431365
transform -1 0 6160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1650_
timestamp 1698431365
transform -1 0 30912 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1651_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1652_
timestamp 1698431365
transform -1 0 29568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1653_
timestamp 1698431365
transform -1 0 12432 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1654_
timestamp 1698431365
transform 1 0 10080 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1655_
timestamp 1698431365
transform -1 0 8288 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1656_
timestamp 1698431365
transform -1 0 28672 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1657_
timestamp 1698431365
transform 1 0 17808 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1658_
timestamp 1698431365
transform -1 0 23296 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1659_
timestamp 1698431365
transform 1 0 23072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1660_
timestamp 1698431365
transform -1 0 19376 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1661_
timestamp 1698431365
transform 1 0 3584 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1662_
timestamp 1698431365
transform -1 0 2912 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1663_
timestamp 1698431365
transform 1 0 29232 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1664_
timestamp 1698431365
transform 1 0 17136 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1665_
timestamp 1698431365
transform 1 0 6272 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1666_
timestamp 1698431365
transform -1 0 6160 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1667_
timestamp 1698431365
transform 1 0 18592 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1668_
timestamp 1698431365
transform -1 0 22288 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1669_
timestamp 1698431365
transform -1 0 18256 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1670_
timestamp 1698431365
transform 1 0 18032 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1671_
timestamp 1698431365
transform 1 0 20048 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1672_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1673_
timestamp 1698431365
transform 1 0 23408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1674_
timestamp 1698431365
transform -1 0 13664 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1675_
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1676_
timestamp 1698431365
transform -1 0 14000 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1677_
timestamp 1698431365
transform 1 0 10976 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1678_
timestamp 1698431365
transform -1 0 11088 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1679_
timestamp 1698431365
transform 1 0 26208 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1680_
timestamp 1698431365
transform 1 0 24192 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1681_
timestamp 1698431365
transform -1 0 25424 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1682_
timestamp 1698431365
transform -1 0 13888 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1683_
timestamp 1698431365
transform 1 0 14560 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1684_
timestamp 1698431365
transform 1 0 13888 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1685_
timestamp 1698431365
transform 1 0 11648 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1686_
timestamp 1698431365
transform -1 0 11424 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1687_
timestamp 1698431365
transform 1 0 21840 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1688_
timestamp 1698431365
transform -1 0 21616 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1689_
timestamp 1698431365
transform 1 0 17696 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1690_
timestamp 1698431365
transform 1 0 10528 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1691_
timestamp 1698431365
transform 1 0 9856 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1692_
timestamp 1698431365
transform 1 0 10304 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1693_
timestamp 1698431365
transform -1 0 10304 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1694_
timestamp 1698431365
transform 1 0 22736 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1695_
timestamp 1698431365
transform 1 0 18816 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1696_
timestamp 1698431365
transform 1 0 19712 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1697_
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1698_
timestamp 1698431365
transform -1 0 22512 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1699_
timestamp 1698431365
transform 1 0 18816 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1700_
timestamp 1698431365
transform -1 0 18816 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1701_
timestamp 1698431365
transform -1 0 22288 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1702_
timestamp 1698431365
transform -1 0 22960 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1703_
timestamp 1698431365
transform -1 0 16800 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1704_
timestamp 1698431365
transform -1 0 18704 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1705_
timestamp 1698431365
transform 1 0 13776 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1706_
timestamp 1698431365
transform -1 0 14000 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1707_
timestamp 1698431365
transform 1 0 12656 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1708_
timestamp 1698431365
transform 1 0 11984 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1709_
timestamp 1698431365
transform -1 0 11760 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1710_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1711_
timestamp 1698431365
transform -1 0 19824 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1712_
timestamp 1698431365
transform 1 0 17360 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1713_
timestamp 1698431365
transform 1 0 16352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1714_
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1715_
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1716_
timestamp 1698431365
transform -1 0 8176 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1717_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1718_
timestamp 1698431365
transform -1 0 2912 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1719_
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1720_
timestamp 1698431365
transform -1 0 4816 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1721_
timestamp 1698431365
transform 1 0 30800 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1722_
timestamp 1698431365
transform 1 0 49616 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1723_
timestamp 1698431365
transform -1 0 46480 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1724_
timestamp 1698431365
transform -1 0 26880 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1725_
timestamp 1698431365
transform -1 0 25088 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1726_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18032 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1727_
timestamp 1698431365
transform -1 0 15568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1728_
timestamp 1698431365
transform 1 0 14112 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1729_
timestamp 1698431365
transform -1 0 14560 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1730_
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1731_
timestamp 1698431365
transform -1 0 10864 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1732_
timestamp 1698431365
transform -1 0 8624 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1733_
timestamp 1698431365
transform -1 0 10640 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1734_
timestamp 1698431365
transform 1 0 6832 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1735_
timestamp 1698431365
transform -1 0 6832 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1736_
timestamp 1698431365
transform -1 0 10080 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1737_
timestamp 1698431365
transform 1 0 7056 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1738_
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1739_
timestamp 1698431365
transform -1 0 26208 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1740_
timestamp 1698431365
transform -1 0 7952 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1741_
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1742_
timestamp 1698431365
transform -1 0 2912 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1743_
timestamp 1698431365
transform 1 0 5936 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1744_
timestamp 1698431365
transform -1 0 4368 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1745_
timestamp 1698431365
transform -1 0 8512 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1746_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1747_
timestamp 1698431365
transform -1 0 3808 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1748_
timestamp 1698431365
transform 1 0 5376 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1749_
timestamp 1698431365
transform -1 0 3024 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1750_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 -1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1751_
timestamp 1698431365
transform -1 0 14336 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1752_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1753_
timestamp 1698431365
transform -1 0 3584 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1754_
timestamp 1698431365
transform 1 0 4816 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1755_
timestamp 1698431365
transform -1 0 4256 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1756_
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1757_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20272 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1758_
timestamp 1698431365
transform 1 0 18704 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1759_
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1760_
timestamp 1698431365
transform -1 0 18704 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1761_
timestamp 1698431365
transform 1 0 19264 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1762_
timestamp 1698431365
transform 1 0 20272 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1763_
timestamp 1698431365
transform -1 0 21952 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1764_
timestamp 1698431365
transform 1 0 17248 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1765_
timestamp 1698431365
transform -1 0 22624 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1766_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20608 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1767_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1768_
timestamp 1698431365
transform 1 0 24752 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1769_
timestamp 1698431365
transform -1 0 18816 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1770_
timestamp 1698431365
transform 1 0 18816 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1771_
timestamp 1698431365
transform 1 0 25200 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1772_
timestamp 1698431365
transform 1 0 30576 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1773_
timestamp 1698431365
transform 1 0 25872 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1774_
timestamp 1698431365
transform -1 0 20720 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1775_
timestamp 1698431365
transform -1 0 21056 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1776_
timestamp 1698431365
transform -1 0 23072 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1777_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22960 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1778_
timestamp 1698431365
transform -1 0 15008 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1779_
timestamp 1698431365
transform -1 0 20944 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1780_
timestamp 1698431365
transform -1 0 13664 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1781_
timestamp 1698431365
transform -1 0 16352 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1782_
timestamp 1698431365
transform 1 0 13664 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1783_
timestamp 1698431365
transform 1 0 27216 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1784_
timestamp 1698431365
transform -1 0 18144 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1785_
timestamp 1698431365
transform 1 0 24192 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1786_
timestamp 1698431365
transform 1 0 26880 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1787_
timestamp 1698431365
transform 1 0 50400 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1788_
timestamp 1698431365
transform -1 0 44912 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1789_
timestamp 1698431365
transform 1 0 44352 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1790_
timestamp 1698431365
transform -1 0 46144 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1791_
timestamp 1698431365
transform -1 0 45584 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1792_
timestamp 1698431365
transform 1 0 43568 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1793_
timestamp 1698431365
transform -1 0 49504 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1794_
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1795_
timestamp 1698431365
transform 1 0 45696 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1796_
timestamp 1698431365
transform 1 0 48384 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1797_
timestamp 1698431365
transform -1 0 47600 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1798_
timestamp 1698431365
transform -1 0 46480 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1799_
timestamp 1698431365
transform -1 0 43568 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1800_
timestamp 1698431365
transform -1 0 48384 0 1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1801_
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1802_
timestamp 1698431365
transform 1 0 49952 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1803_
timestamp 1698431365
transform 1 0 51072 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1804_
timestamp 1698431365
transform 1 0 49504 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1805_
timestamp 1698431365
transform -1 0 50288 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1806_
timestamp 1698431365
transform 1 0 50288 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1807_
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1808_
timestamp 1698431365
transform 1 0 49168 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1809_
timestamp 1698431365
transform -1 0 50176 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1810_
timestamp 1698431365
transform -1 0 51296 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1811_
timestamp 1698431365
transform 1 0 49616 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1812_
timestamp 1698431365
transform -1 0 50736 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1813_
timestamp 1698431365
transform -1 0 49392 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1814_
timestamp 1698431365
transform 1 0 49728 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1815_
timestamp 1698431365
transform -1 0 52080 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1816_
timestamp 1698431365
transform 1 0 50176 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1817_
timestamp 1698431365
transform 1 0 50400 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1818_
timestamp 1698431365
transform -1 0 34272 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1819_
timestamp 1698431365
transform 1 0 26320 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1820_
timestamp 1698431365
transform -1 0 34272 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1821_
timestamp 1698431365
transform -1 0 34496 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1822_
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1823_
timestamp 1698431365
transform -1 0 38752 0 1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1824_
timestamp 1698431365
transform -1 0 36624 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1825_
timestamp 1698431365
transform -1 0 37632 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1826_
timestamp 1698431365
transform -1 0 36736 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1827_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36736 0 -1 34496
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1828_
timestamp 1698431365
transform -1 0 37856 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1829_
timestamp 1698431365
transform 1 0 37856 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1830_
timestamp 1698431365
transform 1 0 39312 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1831_
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1832_
timestamp 1698431365
transform -1 0 36400 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1833_
timestamp 1698431365
transform -1 0 36736 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1834_
timestamp 1698431365
transform 1 0 37184 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1835_
timestamp 1698431365
transform -1 0 38976 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1836_
timestamp 1698431365
transform 1 0 37744 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1837_
timestamp 1698431365
transform -1 0 38864 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1838_
timestamp 1698431365
transform 1 0 37856 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1839_
timestamp 1698431365
transform 1 0 39200 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1840_
timestamp 1698431365
transform 1 0 29344 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1841_
timestamp 1698431365
transform 1 0 36736 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1842_
timestamp 1698431365
transform -1 0 37520 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1843_
timestamp 1698431365
transform -1 0 38416 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1844_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37856 0 -1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1845_
timestamp 1698431365
transform 1 0 38752 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1846_
timestamp 1698431365
transform -1 0 41440 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1847_
timestamp 1698431365
transform -1 0 40544 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1848_
timestamp 1698431365
transform -1 0 40544 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1849_
timestamp 1698431365
transform 1 0 38080 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1850_
timestamp 1698431365
transform 1 0 39424 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1851_
timestamp 1698431365
transform -1 0 40544 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1852_
timestamp 1698431365
transform -1 0 41664 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1853_
timestamp 1698431365
transform -1 0 41888 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1698431365
transform 1 0 41888 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1855_
timestamp 1698431365
transform 1 0 42336 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1856_
timestamp 1698431365
transform 1 0 43568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1857_
timestamp 1698431365
transform 1 0 34272 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1858_
timestamp 1698431365
transform -1 0 47152 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1859_
timestamp 1698431365
transform -1 0 40320 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1860_
timestamp 1698431365
transform -1 0 39424 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1861_
timestamp 1698431365
transform -1 0 40320 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1862_
timestamp 1698431365
transform -1 0 38976 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1863_
timestamp 1698431365
transform 1 0 38528 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1864_
timestamp 1698431365
transform 1 0 39424 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1865_
timestamp 1698431365
transform -1 0 40320 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1866_
timestamp 1698431365
transform -1 0 39984 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1867_
timestamp 1698431365
transform 1 0 36960 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1868_
timestamp 1698431365
transform 1 0 53200 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1869_
timestamp 1698431365
transform 1 0 48944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1870_
timestamp 1698431365
transform -1 0 49280 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform 1 0 49616 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1872_
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1873_
timestamp 1698431365
transform -1 0 55104 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1874_
timestamp 1698431365
transform 1 0 45136 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1875_
timestamp 1698431365
transform 1 0 43680 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1876_
timestamp 1698431365
transform 1 0 49952 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1877_
timestamp 1698431365
transform 1 0 50512 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1878_
timestamp 1698431365
transform 1 0 51744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1879_
timestamp 1698431365
transform -1 0 56112 0 -1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1880_
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1881_
timestamp 1698431365
transform -1 0 52304 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1882_
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1883_
timestamp 1698431365
transform -1 0 48608 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1884_
timestamp 1698431365
transform -1 0 54208 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1885_
timestamp 1698431365
transform -1 0 55776 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1886_
timestamp 1698431365
transform -1 0 48384 0 -1 26656
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1887_
timestamp 1698431365
transform 1 0 45584 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1888_
timestamp 1698431365
transform 1 0 44912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1889_
timestamp 1698431365
transform 1 0 48496 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1890_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42784 0 -1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1891_
timestamp 1698431365
transform 1 0 46928 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1892_
timestamp 1698431365
transform 1 0 44016 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1893_
timestamp 1698431365
transform -1 0 55104 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1894_
timestamp 1698431365
transform 1 0 45696 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1895_
timestamp 1698431365
transform -1 0 47600 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1896_
timestamp 1698431365
transform -1 0 46928 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1897_
timestamp 1698431365
transform -1 0 38416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1898_
timestamp 1698431365
transform -1 0 36064 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1899_
timestamp 1698431365
transform 1 0 42896 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1900_
timestamp 1698431365
transform 1 0 39088 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1901_
timestamp 1698431365
transform -1 0 40432 0 -1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1902_
timestamp 1698431365
transform 1 0 37296 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1903_
timestamp 1698431365
transform 1 0 46592 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1904_
timestamp 1698431365
transform -1 0 49280 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1905_
timestamp 1698431365
transform 1 0 40768 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1906_
timestamp 1698431365
transform 1 0 39424 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1907_
timestamp 1698431365
transform -1 0 39424 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1908_
timestamp 1698431365
transform 1 0 38304 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1909_
timestamp 1698431365
transform 1 0 40320 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1910_
timestamp 1698431365
transform -1 0 42560 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1911_
timestamp 1698431365
transform 1 0 42112 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1912_
timestamp 1698431365
transform 1 0 45584 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1913_
timestamp 1698431365
transform 1 0 46368 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1914_
timestamp 1698431365
transform -1 0 46592 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1915_
timestamp 1698431365
transform 1 0 43792 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1916_
timestamp 1698431365
transform 1 0 43680 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1917_
timestamp 1698431365
transform 1 0 39872 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1918_
timestamp 1698431365
transform 1 0 41664 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1919_
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1920_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1921_
timestamp 1698431365
transform 1 0 41440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1922_
timestamp 1698431365
transform 1 0 42784 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1923_
timestamp 1698431365
transform 1 0 48384 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1924_
timestamp 1698431365
transform 1 0 40880 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1925_
timestamp 1698431365
transform -1 0 44016 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1926_
timestamp 1698431365
transform 1 0 42224 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1927_
timestamp 1698431365
transform 1 0 42112 0 1 39200
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1928_
timestamp 1698431365
transform 1 0 44352 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1929_
timestamp 1698431365
transform 1 0 43008 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1930_
timestamp 1698431365
transform -1 0 43008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1931_
timestamp 1698431365
transform -1 0 45696 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1932_
timestamp 1698431365
transform 1 0 45696 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1933_
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1934_
timestamp 1698431365
transform -1 0 42112 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1935_
timestamp 1698431365
transform 1 0 42000 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1936_
timestamp 1698431365
transform 1 0 41328 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1937_
timestamp 1698431365
transform -1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1938_
timestamp 1698431365
transform -1 0 44016 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1939_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42000 0 -1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1940_
timestamp 1698431365
transform -1 0 50624 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1941_
timestamp 1698431365
transform 1 0 49056 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1942_
timestamp 1698431365
transform 1 0 46256 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1943_
timestamp 1698431365
transform 1 0 46704 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1944_
timestamp 1698431365
transform 1 0 47264 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1945_
timestamp 1698431365
transform 1 0 45808 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1946_
timestamp 1698431365
transform 1 0 49504 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1947_
timestamp 1698431365
transform 1 0 48608 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1948_
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1949_
timestamp 1698431365
transform 1 0 50400 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1950_
timestamp 1698431365
transform -1 0 52192 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1951_
timestamp 1698431365
transform 1 0 50960 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1698431365
transform -1 0 50288 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1953_
timestamp 1698431365
transform 1 0 51184 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1954_
timestamp 1698431365
transform -1 0 52640 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1955_
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1956_
timestamp 1698431365
transform -1 0 51184 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1698431365
transform 1 0 49392 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1958_
timestamp 1698431365
transform 1 0 46144 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1959_
timestamp 1698431365
transform -1 0 48272 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1960_
timestamp 1698431365
transform 1 0 50288 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1961_
timestamp 1698431365
transform 1 0 51744 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1962_
timestamp 1698431365
transform 1 0 50848 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1963_
timestamp 1698431365
transform 1 0 52640 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1964_
timestamp 1698431365
transform 1 0 54432 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1965_
timestamp 1698431365
transform -1 0 48272 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1966_
timestamp 1698431365
transform 1 0 45360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1967_
timestamp 1698431365
transform -1 0 40432 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1968_
timestamp 1698431365
transform -1 0 45360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1969_
timestamp 1698431365
transform -1 0 44240 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1970_
timestamp 1698431365
transform 1 0 32928 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1971_
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1972_
timestamp 1698431365
transform -1 0 52080 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1973_
timestamp 1698431365
transform 1 0 49840 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1974_
timestamp 1698431365
transform 1 0 45920 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1975_
timestamp 1698431365
transform 1 0 47376 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1976_
timestamp 1698431365
transform -1 0 51184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1977_
timestamp 1698431365
transform -1 0 49056 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1978_
timestamp 1698431365
transform 1 0 47264 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1979_
timestamp 1698431365
transform -1 0 50400 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1980_
timestamp 1698431365
transform -1 0 49280 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1981_
timestamp 1698431365
transform -1 0 47488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1982_
timestamp 1698431365
transform -1 0 49504 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1983_
timestamp 1698431365
transform -1 0 53648 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1984_
timestamp 1698431365
transform 1 0 51520 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1985_
timestamp 1698431365
transform 1 0 53760 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1986_
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1987_
timestamp 1698431365
transform 1 0 54432 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1988_
timestamp 1698431365
transform -1 0 56000 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1989_
timestamp 1698431365
transform 1 0 54320 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1990_
timestamp 1698431365
transform 1 0 49056 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1991_
timestamp 1698431365
transform 1 0 49392 0 -1 36064
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1992_
timestamp 1698431365
transform 1 0 46928 0 1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1993_
timestamp 1698431365
transform 1 0 47488 0 1 34496
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1994_
timestamp 1698431365
transform 1 0 54880 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1995_
timestamp 1698431365
transform 1 0 56896 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1996_
timestamp 1698431365
transform 1 0 56448 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1997_
timestamp 1698431365
transform -1 0 58016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1998_
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1698431365
transform 1 0 56000 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2000_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 53872 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2001_
timestamp 1698431365
transform 1 0 57568 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2002_
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2003_
timestamp 1698431365
transform -1 0 39872 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2004_
timestamp 1698431365
transform 1 0 40432 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2005_
timestamp 1698431365
transform 1 0 52864 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2006_
timestamp 1698431365
transform -1 0 57120 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2007_
timestamp 1698431365
transform -1 0 54656 0 -1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2008_
timestamp 1698431365
transform 1 0 53760 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2009_
timestamp 1698431365
transform 1 0 50288 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2010_
timestamp 1698431365
transform -1 0 54320 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2011_
timestamp 1698431365
transform -1 0 55328 0 -1 34496
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2012_
timestamp 1698431365
transform 1 0 49952 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2013_
timestamp 1698431365
transform -1 0 50400 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2014_
timestamp 1698431365
transform -1 0 50736 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2015_
timestamp 1698431365
transform 1 0 31472 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2016_
timestamp 1698431365
transform -1 0 51744 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2017_
timestamp 1698431365
transform -1 0 42784 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2018_
timestamp 1698431365
transform 1 0 47264 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2019_
timestamp 1698431365
transform -1 0 49840 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2020_
timestamp 1698431365
transform -1 0 52640 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2021_
timestamp 1698431365
transform 1 0 53312 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2022_
timestamp 1698431365
transform -1 0 56784 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2023_
timestamp 1698431365
transform -1 0 55552 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2024_
timestamp 1698431365
transform -1 0 52304 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2025_
timestamp 1698431365
transform -1 0 45808 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2026_
timestamp 1698431365
transform -1 0 45248 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2027_
timestamp 1698431365
transform 1 0 43568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2028_
timestamp 1698431365
transform -1 0 43008 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2029_
timestamp 1698431365
transform -1 0 48048 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2030_
timestamp 1698431365
transform -1 0 54208 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2031_
timestamp 1698431365
transform -1 0 56112 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2032_
timestamp 1698431365
transform -1 0 53200 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2033_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2034_
timestamp 1698431365
transform -1 0 45920 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2035_
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2036_
timestamp 1698431365
transform -1 0 51184 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2037_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 54656 0 1 28224
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2038_
timestamp 1698431365
transform 1 0 49728 0 -1 29792
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2039_
timestamp 1698431365
transform -1 0 51632 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2040_
timestamp 1698431365
transform -1 0 50064 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2041_
timestamp 1698431365
transform -1 0 51744 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2042_
timestamp 1698431365
transform 1 0 51408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2043_
timestamp 1698431365
transform -1 0 53200 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2044_
timestamp 1698431365
transform -1 0 52304 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2045_
timestamp 1698431365
transform -1 0 49280 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2046_
timestamp 1698431365
transform -1 0 50624 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2047_
timestamp 1698431365
transform 1 0 49280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2048_
timestamp 1698431365
transform -1 0 49728 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2049_
timestamp 1698431365
transform -1 0 52640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2050_
timestamp 1698431365
transform -1 0 50400 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2051_
timestamp 1698431365
transform -1 0 51856 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2052_
timestamp 1698431365
transform 1 0 51632 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2053_
timestamp 1698431365
transform -1 0 54432 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2054_
timestamp 1698431365
transform -1 0 50960 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2055_
timestamp 1698431365
transform 1 0 51184 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2056_
timestamp 1698431365
transform 1 0 49840 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2057_
timestamp 1698431365
transform 1 0 51520 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2058_
timestamp 1698431365
transform 1 0 50400 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2059_
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2060_
timestamp 1698431365
transform -1 0 35056 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2061_
timestamp 1698431365
transform 1 0 46928 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2062_
timestamp 1698431365
transform -1 0 53536 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2063_
timestamp 1698431365
transform -1 0 49504 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2064_
timestamp 1698431365
transform 1 0 50064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2065_
timestamp 1698431365
transform -1 0 48272 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2066_
timestamp 1698431365
transform -1 0 46032 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2067_
timestamp 1698431365
transform -1 0 48384 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2068_
timestamp 1698431365
transform -1 0 48160 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2069_
timestamp 1698431365
transform 1 0 49056 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2070_
timestamp 1698431365
transform 1 0 45808 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2071_
timestamp 1698431365
transform 1 0 46032 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2072_
timestamp 1698431365
transform 1 0 47152 0 1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2073_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2074_
timestamp 1698431365
transform 1 0 47488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2075_
timestamp 1698431365
transform -1 0 47936 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2076_
timestamp 1698431365
transform 1 0 48160 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2077_
timestamp 1698431365
transform -1 0 48944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2078_
timestamp 1698431365
transform 1 0 46032 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2079_
timestamp 1698431365
transform -1 0 47488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2080_
timestamp 1698431365
transform 1 0 46816 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2081_
timestamp 1698431365
transform 1 0 45920 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2082_
timestamp 1698431365
transform -1 0 44352 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2083_
timestamp 1698431365
transform -1 0 49840 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2084_
timestamp 1698431365
transform -1 0 44464 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2085_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2086_
timestamp 1698431365
transform 1 0 43568 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2087_
timestamp 1698431365
transform -1 0 44464 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2088_
timestamp 1698431365
transform -1 0 43680 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2089_
timestamp 1698431365
transform 1 0 40992 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2090_
timestamp 1698431365
transform 1 0 42000 0 -1 25088
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2091_
timestamp 1698431365
transform 1 0 42560 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2092_
timestamp 1698431365
transform 1 0 42112 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2093_
timestamp 1698431365
transform -1 0 42560 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2094_
timestamp 1698431365
transform -1 0 41440 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2095_
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2096_
timestamp 1698431365
transform -1 0 45808 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2097_
timestamp 1698431365
transform -1 0 42896 0 -1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2098_
timestamp 1698431365
transform 1 0 45920 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2099_
timestamp 1698431365
transform -1 0 40544 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2100_
timestamp 1698431365
transform -1 0 42560 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2101_
timestamp 1698431365
transform 1 0 40656 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2102_
timestamp 1698431365
transform 1 0 39312 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2103_
timestamp 1698431365
transform -1 0 39312 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2104_
timestamp 1698431365
transform 1 0 39424 0 1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2105_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2106_
timestamp 1698431365
transform -1 0 43344 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2107_
timestamp 1698431365
transform 1 0 41888 0 -1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2108_
timestamp 1698431365
transform -1 0 35280 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2109_
timestamp 1698431365
transform 1 0 37968 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2110_
timestamp 1698431365
transform -1 0 39088 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2111_
timestamp 1698431365
transform 1 0 39088 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2112_
timestamp 1698431365
transform -1 0 37520 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2113_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2114_
timestamp 1698431365
transform -1 0 41888 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2115_
timestamp 1698431365
transform 1 0 34048 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2116_
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2117_
timestamp 1698431365
transform 1 0 35280 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2118_
timestamp 1698431365
transform 1 0 35952 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2119_
timestamp 1698431365
transform 1 0 34832 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2120_
timestamp 1698431365
transform -1 0 37520 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2121_
timestamp 1698431365
transform -1 0 40208 0 -1 25088
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2122_
timestamp 1698431365
transform -1 0 38304 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2123_
timestamp 1698431365
transform -1 0 38192 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2124_
timestamp 1698431365
transform -1 0 36624 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2125_
timestamp 1698431365
transform -1 0 33040 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2126_
timestamp 1698431365
transform -1 0 36624 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2127_
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2128_
timestamp 1698431365
transform -1 0 34944 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2129_
timestamp 1698431365
transform 1 0 31920 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2130_
timestamp 1698431365
transform -1 0 33936 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2131_
timestamp 1698431365
transform 1 0 33936 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2132_
timestamp 1698431365
transform 1 0 31808 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2133_
timestamp 1698431365
transform -1 0 34160 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2134_
timestamp 1698431365
transform 1 0 31360 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2135_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2136_
timestamp 1698431365
transform 1 0 31808 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2137_
timestamp 1698431365
transform 1 0 32816 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2138_
timestamp 1698431365
transform 1 0 31808 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2139_
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2140_
timestamp 1698431365
transform -1 0 34384 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2141_
timestamp 1698431365
transform -1 0 35728 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2142_
timestamp 1698431365
transform -1 0 34272 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2143_
timestamp 1698431365
transform -1 0 32704 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2144_
timestamp 1698431365
transform 1 0 33152 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2145_
timestamp 1698431365
transform 1 0 33040 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2146_
timestamp 1698431365
transform -1 0 35504 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2147_
timestamp 1698431365
transform -1 0 34944 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2148_
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2149_
timestamp 1698431365
transform 1 0 44240 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2150_
timestamp 1698431365
transform -1 0 46480 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2151_
timestamp 1698431365
transform 1 0 18928 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2152_
timestamp 1698431365
transform 1 0 20272 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2153_
timestamp 1698431365
transform 1 0 34272 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2154_
timestamp 1698431365
transform -1 0 34832 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2155_
timestamp 1698431365
transform -1 0 29120 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2156_
timestamp 1698431365
transform 1 0 27776 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2157_
timestamp 1698431365
transform -1 0 23856 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2158_
timestamp 1698431365
transform -1 0 20944 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2159_
timestamp 1698431365
transform 1 0 19040 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2160_
timestamp 1698431365
transform 1 0 26656 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2161_
timestamp 1698431365
transform -1 0 26432 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2162_
timestamp 1698431365
transform 1 0 16912 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2163_
timestamp 1698431365
transform 1 0 17808 0 -1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2164_
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2165_
timestamp 1698431365
transform 1 0 29904 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2166_
timestamp 1698431365
transform 1 0 28224 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2167_
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2168_
timestamp 1698431365
transform -1 0 30912 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2169_
timestamp 1698431365
transform -1 0 32928 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2170_
timestamp 1698431365
transform -1 0 33376 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2171_
timestamp 1698431365
transform -1 0 31696 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2172_
timestamp 1698431365
transform -1 0 26208 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2173_
timestamp 1698431365
transform -1 0 16576 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2174_
timestamp 1698431365
transform -1 0 18816 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2175_
timestamp 1698431365
transform 1 0 18928 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _2176_
timestamp 1698431365
transform 1 0 14224 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2177_
timestamp 1698431365
transform -1 0 24192 0 -1 45472
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2178_
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2179_
timestamp 1698431365
transform -1 0 18256 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2180_
timestamp 1698431365
transform 1 0 21504 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2181_
timestamp 1698431365
transform 1 0 27440 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2182_
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2183_
timestamp 1698431365
transform 1 0 27328 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2184_
timestamp 1698431365
transform -1 0 29904 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2185_
timestamp 1698431365
transform 1 0 30016 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2186_
timestamp 1698431365
transform -1 0 33600 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2187_
timestamp 1698431365
transform -1 0 29456 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2188_
timestamp 1698431365
transform 1 0 26208 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2189_
timestamp 1698431365
transform -1 0 24864 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2190_
timestamp 1698431365
transform 1 0 25200 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2191_
timestamp 1698431365
transform 1 0 27216 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2192_
timestamp 1698431365
transform 1 0 28336 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2193_
timestamp 1698431365
transform 1 0 27888 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2194_
timestamp 1698431365
transform 1 0 27888 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2195_
timestamp 1698431365
transform 1 0 31584 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2196_
timestamp 1698431365
transform 1 0 30688 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2197_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29792 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2198_
timestamp 1698431365
transform 1 0 20048 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2199_
timestamp 1698431365
transform 1 0 21952 0 -1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2200_
timestamp 1698431365
transform -1 0 22064 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2201_
timestamp 1698431365
transform -1 0 23632 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2202_
timestamp 1698431365
transform -1 0 22624 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2203_
timestamp 1698431365
transform 1 0 22624 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2204_
timestamp 1698431365
transform 1 0 28560 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2205_
timestamp 1698431365
transform -1 0 30016 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2206_
timestamp 1698431365
transform 1 0 29904 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2207_
timestamp 1698431365
transform 1 0 32256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2208_
timestamp 1698431365
transform 1 0 32368 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2209_
timestamp 1698431365
transform 1 0 30576 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2210_
timestamp 1698431365
transform 1 0 26096 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2211_
timestamp 1698431365
transform -1 0 27664 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2212_
timestamp 1698431365
transform 1 0 27888 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2213_
timestamp 1698431365
transform 1 0 29904 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2214_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29344 0 -1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2215_
timestamp 1698431365
transform 1 0 30128 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2216_
timestamp 1698431365
transform -1 0 30800 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2217_
timestamp 1698431365
transform 1 0 25536 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2218_
timestamp 1698431365
transform 1 0 27888 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2219_
timestamp 1698431365
transform 1 0 26096 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2220_
timestamp 1698431365
transform -1 0 25760 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2221_
timestamp 1698431365
transform -1 0 28112 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2222_
timestamp 1698431365
transform -1 0 27664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2223_
timestamp 1698431365
transform 1 0 26432 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2224_
timestamp 1698431365
transform 1 0 26656 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2225_
timestamp 1698431365
transform 1 0 23968 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2226_
timestamp 1698431365
transform 1 0 10976 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2227_
timestamp 1698431365
transform 1 0 14224 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2228_
timestamp 1698431365
transform 1 0 15568 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2229_
timestamp 1698431365
transform 1 0 25760 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2230_
timestamp 1698431365
transform 1 0 24416 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2231_
timestamp 1698431365
transform -1 0 20272 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2232_
timestamp 1698431365
transform 1 0 31584 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2233_
timestamp 1698431365
transform -1 0 31584 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2234_
timestamp 1698431365
transform -1 0 28000 0 1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2235_
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2236_
timestamp 1698431365
transform 1 0 29120 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2237_
timestamp 1698431365
transform -1 0 29680 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2238_
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2239_
timestamp 1698431365
transform 1 0 22400 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2240_
timestamp 1698431365
transform 1 0 23296 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2241_
timestamp 1698431365
transform 1 0 29792 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2242_
timestamp 1698431365
transform 1 0 30128 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2243_
timestamp 1698431365
transform -1 0 30128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2244_
timestamp 1698431365
transform 1 0 21840 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2245_
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2246_
timestamp 1698431365
transform -1 0 33600 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2247_
timestamp 1698431365
transform -1 0 33040 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2248_
timestamp 1698431365
transform 1 0 32032 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2249_
timestamp 1698431365
transform 1 0 28112 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2250_
timestamp 1698431365
transform 1 0 28784 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2251_
timestamp 1698431365
transform 1 0 16128 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2252_
timestamp 1698431365
transform -1 0 16128 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2253_
timestamp 1698431365
transform 1 0 24976 0 1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2254_
timestamp 1698431365
transform 1 0 28896 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2255_
timestamp 1698431365
transform 1 0 17472 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2256_
timestamp 1698431365
transform 1 0 19936 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2257_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28224 0 -1 45472
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2258_
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2259_
timestamp 1698431365
transform -1 0 34384 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2260_
timestamp 1698431365
transform 1 0 33600 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2261_
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2262_
timestamp 1698431365
transform -1 0 28000 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2263_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25648 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2264_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2265_
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2266_
timestamp 1698431365
transform -1 0 31248 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2267_
timestamp 1698431365
transform 1 0 34384 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2268_
timestamp 1698431365
transform -1 0 34496 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2269_
timestamp 1698431365
transform 1 0 25200 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2270_
timestamp 1698431365
transform 1 0 26656 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2271_
timestamp 1698431365
transform 1 0 32368 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2272_
timestamp 1698431365
transform 1 0 33376 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2273_
timestamp 1698431365
transform 1 0 34272 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2274_
timestamp 1698431365
transform -1 0 28784 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2275_
timestamp 1698431365
transform 1 0 31248 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2276_
timestamp 1698431365
transform 1 0 30688 0 -1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2277_
timestamp 1698431365
transform 1 0 30800 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2278_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2279_
timestamp 1698431365
transform 1 0 38080 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2280_
timestamp 1698431365
transform 1 0 26992 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2281_
timestamp 1698431365
transform 1 0 26432 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2282_
timestamp 1698431365
transform -1 0 29792 0 1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2283_
timestamp 1698431365
transform -1 0 29008 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2284_
timestamp 1698431365
transform -1 0 29904 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2285_
timestamp 1698431365
transform 1 0 35504 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2286_
timestamp 1698431365
transform -1 0 35728 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2287_
timestamp 1698431365
transform -1 0 35952 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2288_
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2289_
timestamp 1698431365
transform -1 0 24864 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2290_
timestamp 1698431365
transform -1 0 28784 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2291_
timestamp 1698431365
transform 1 0 28112 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2292_
timestamp 1698431365
transform 1 0 34384 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2293_
timestamp 1698431365
transform 1 0 35728 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2294_
timestamp 1698431365
transform -1 0 32704 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2295_
timestamp 1698431365
transform 1 0 26544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2296_
timestamp 1698431365
transform 1 0 27552 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2297_
timestamp 1698431365
transform 1 0 29792 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2298_
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2299_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2300_
timestamp 1698431365
transform 1 0 14336 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2301_
timestamp 1698431365
transform 1 0 18368 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2302_
timestamp 1698431365
transform 1 0 19040 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2303_
timestamp 1698431365
transform 1 0 19152 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2304_
timestamp 1698431365
transform -1 0 19712 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2305_
timestamp 1698431365
transform -1 0 13104 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2306_
timestamp 1698431365
transform -1 0 7728 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2307_
timestamp 1698431365
transform -1 0 7840 0 1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2308_
timestamp 1698431365
transform 1 0 4256 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2309_
timestamp 1698431365
transform -1 0 8512 0 -1 51744
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2310_
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2311_
timestamp 1698431365
transform 1 0 6160 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2312_
timestamp 1698431365
transform 1 0 4816 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2313_
timestamp 1698431365
transform 1 0 3248 0 -1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2314_
timestamp 1698431365
transform -1 0 7280 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2315_
timestamp 1698431365
transform 1 0 8512 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2316_
timestamp 1698431365
transform 1 0 10976 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2317_
timestamp 1698431365
transform 1 0 11312 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2318_
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2319_
timestamp 1698431365
transform -1 0 15232 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2320_
timestamp 1698431365
transform 1 0 12096 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2321_
timestamp 1698431365
transform 1 0 16800 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2322_
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2323_
timestamp 1698431365
transform -1 0 19488 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2324_
timestamp 1698431365
transform -1 0 17024 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2325_
timestamp 1698431365
transform -1 0 13552 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2326_
timestamp 1698431365
transform -1 0 12432 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2327_
timestamp 1698431365
transform 1 0 9968 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2328_
timestamp 1698431365
transform -1 0 14672 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2329_
timestamp 1698431365
transform -1 0 10864 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2330_
timestamp 1698431365
transform -1 0 19040 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2331_
timestamp 1698431365
transform -1 0 17920 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2332_
timestamp 1698431365
transform -1 0 15680 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2333_
timestamp 1698431365
transform -1 0 9184 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2334_
timestamp 1698431365
transform 1 0 9632 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2335_
timestamp 1698431365
transform -1 0 10416 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2336_
timestamp 1698431365
transform -1 0 15008 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2337_
timestamp 1698431365
transform 1 0 13552 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2338_
timestamp 1698431365
transform 1 0 10752 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2339_
timestamp 1698431365
transform 1 0 9856 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2340_
timestamp 1698431365
transform -1 0 10864 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2341_
timestamp 1698431365
transform 1 0 10864 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2342_
timestamp 1698431365
transform 1 0 10192 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2343_
timestamp 1698431365
transform -1 0 12432 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2344_
timestamp 1698431365
transform -1 0 18256 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2345_
timestamp 1698431365
transform 1 0 15344 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2346_
timestamp 1698431365
transform 1 0 11760 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2347_
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2348_
timestamp 1698431365
transform 1 0 13328 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2349_
timestamp 1698431365
transform 1 0 13440 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2350_
timestamp 1698431365
transform -1 0 14224 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2351_
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2352_
timestamp 1698431365
transform -1 0 19040 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2353_
timestamp 1698431365
transform 1 0 15120 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2354_
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2355_
timestamp 1698431365
transform -1 0 17024 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2356_
timestamp 1698431365
transform -1 0 15680 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2357_
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2358_
timestamp 1698431365
transform -1 0 16800 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2359_
timestamp 1698431365
transform -1 0 16912 0 -1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2360_
timestamp 1698431365
transform -1 0 10528 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2361_
timestamp 1698431365
transform -1 0 8400 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2362_
timestamp 1698431365
transform 1 0 2464 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2363_
timestamp 1698431365
transform -1 0 4256 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2364_
timestamp 1698431365
transform -1 0 2800 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2365_
timestamp 1698431365
transform 1 0 3808 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2366_
timestamp 1698431365
transform 1 0 4032 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2367_
timestamp 1698431365
transform 1 0 3136 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2368_
timestamp 1698431365
transform 1 0 4032 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2369_
timestamp 1698431365
transform 1 0 5712 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2370_
timestamp 1698431365
transform 1 0 7168 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2371_
timestamp 1698431365
transform -1 0 6832 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2372_
timestamp 1698431365
transform 1 0 6832 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2373_
timestamp 1698431365
transform -1 0 7280 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2374_
timestamp 1698431365
transform -1 0 6384 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2375_
timestamp 1698431365
transform -1 0 4368 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2376_
timestamp 1698431365
transform 1 0 4368 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2377_
timestamp 1698431365
transform 1 0 7504 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2378_
timestamp 1698431365
transform 1 0 5712 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2379_
timestamp 1698431365
transform -1 0 7504 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2380_
timestamp 1698431365
transform -1 0 6160 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2381_
timestamp 1698431365
transform -1 0 6832 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2382_
timestamp 1698431365
transform 1 0 6832 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2383_
timestamp 1698431365
transform -1 0 6160 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2384_
timestamp 1698431365
transform -1 0 6944 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2385_
timestamp 1698431365
transform 1 0 6272 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2386_
timestamp 1698431365
transform 1 0 4816 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2387_
timestamp 1698431365
transform -1 0 7840 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2388_
timestamp 1698431365
transform -1 0 6944 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2389_
timestamp 1698431365
transform -1 0 5712 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2390_
timestamp 1698431365
transform 1 0 3920 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2391_
timestamp 1698431365
transform 1 0 3248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2392_
timestamp 1698431365
transform 1 0 4928 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2393_
timestamp 1698431365
transform 1 0 4144 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2394_
timestamp 1698431365
transform 1 0 4256 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2395_
timestamp 1698431365
transform 1 0 6720 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2396_
timestamp 1698431365
transform -1 0 6048 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2397_
timestamp 1698431365
transform 1 0 5824 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2398_
timestamp 1698431365
transform -1 0 5152 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2399_
timestamp 1698431365
transform -1 0 4256 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2400_
timestamp 1698431365
transform -1 0 3360 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2401_
timestamp 1698431365
transform -1 0 4704 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2402_
timestamp 1698431365
transform -1 0 4144 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2403_
timestamp 1698431365
transform -1 0 4032 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2404_
timestamp 1698431365
transform 1 0 2352 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2405_
timestamp 1698431365
transform 1 0 2240 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2406_
timestamp 1698431365
transform -1 0 4256 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2407_
timestamp 1698431365
transform -1 0 3696 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2408_
timestamp 1698431365
transform 1 0 2576 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2409_
timestamp 1698431365
transform 1 0 25760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2410_
timestamp 1698431365
transform -1 0 22848 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2411_
timestamp 1698431365
transform 1 0 22064 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2412_
timestamp 1698431365
transform 1 0 24192 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2413_
timestamp 1698431365
transform 1 0 26992 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2414_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2415_
timestamp 1698431365
transform -1 0 24416 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2416_
timestamp 1698431365
transform -1 0 24528 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2417_
timestamp 1698431365
transform 1 0 21504 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2418_
timestamp 1698431365
transform -1 0 23296 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2419_
timestamp 1698431365
transform -1 0 22512 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2420_
timestamp 1698431365
transform -1 0 21840 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2421_
timestamp 1698431365
transform -1 0 23296 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2422_
timestamp 1698431365
transform -1 0 20832 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2423_
timestamp 1698431365
transform -1 0 19488 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2424_
timestamp 1698431365
transform -1 0 22064 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2425_
timestamp 1698431365
transform 1 0 19712 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2426_
timestamp 1698431365
transform -1 0 21056 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2427_
timestamp 1698431365
transform 1 0 25648 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2428_
timestamp 1698431365
transform -1 0 25760 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2429_
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2430_
timestamp 1698431365
transform 1 0 18592 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2431_
timestamp 1698431365
transform 1 0 13664 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2432_
timestamp 1698431365
transform -1 0 15008 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2433_
timestamp 1698431365
transform -1 0 25200 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2434_
timestamp 1698431365
transform -1 0 23184 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2435_
timestamp 1698431365
transform 1 0 22624 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2436_
timestamp 1698431365
transform -1 0 23072 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2437_
timestamp 1698431365
transform 1 0 18928 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2438_
timestamp 1698431365
transform -1 0 21280 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2439_
timestamp 1698431365
transform -1 0 20384 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2440_
timestamp 1698431365
transform -1 0 20832 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2441_
timestamp 1698431365
transform 1 0 19600 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2442_
timestamp 1698431365
transform -1 0 21504 0 -1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2443_
timestamp 1698431365
transform 1 0 21728 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2444_
timestamp 1698431365
transform -1 0 26656 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2445_
timestamp 1698431365
transform -1 0 23968 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2446_
timestamp 1698431365
transform 1 0 22624 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2447_
timestamp 1698431365
transform 1 0 23520 0 1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2448_
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2449_
timestamp 1698431365
transform 1 0 21952 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2450_
timestamp 1698431365
transform -1 0 25648 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2451_
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2452_
timestamp 1698431365
transform -1 0 25536 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2453_
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2454_
timestamp 1698431365
transform -1 0 23408 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2455_
timestamp 1698431365
transform 1 0 19376 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2456_
timestamp 1698431365
transform 1 0 22400 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2457_
timestamp 1698431365
transform -1 0 24080 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2458_
timestamp 1698431365
transform 1 0 24080 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2459_
timestamp 1698431365
transform 1 0 23520 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2460_
timestamp 1698431365
transform -1 0 24304 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2461_
timestamp 1698431365
transform 1 0 18256 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2462_
timestamp 1698431365
transform 1 0 19824 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2463_
timestamp 1698431365
transform 1 0 21952 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2464_
timestamp 1698431365
transform 1 0 23408 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2465_
timestamp 1698431365
transform 1 0 24080 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2466_
timestamp 1698431365
transform -1 0 24528 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2467_
timestamp 1698431365
transform 1 0 19712 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2468_
timestamp 1698431365
transform 1 0 23296 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2469_
timestamp 1698431365
transform 1 0 23856 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2470_
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2471_
timestamp 1698431365
transform 1 0 29792 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2472_
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2473_
timestamp 1698431365
transform 1 0 33936 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2474_
timestamp 1698431365
transform 1 0 33600 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2475_
timestamp 1698431365
transform 1 0 29456 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2476_
timestamp 1698431365
transform -1 0 36512 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2477_
timestamp 1698431365
transform 1 0 35616 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2478_
timestamp 1698431365
transform -1 0 16352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2479_
timestamp 1698431365
transform -1 0 20496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2480_
timestamp 1698431365
transform 1 0 17808 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2481_
timestamp 1698431365
transform -1 0 17920 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2482_
timestamp 1698431365
transform -1 0 19264 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2483_
timestamp 1698431365
transform 1 0 18032 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2484_
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2485_
timestamp 1698431365
transform -1 0 13104 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2486_
timestamp 1698431365
transform 1 0 12096 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2487_
timestamp 1698431365
transform -1 0 10416 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2488_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2489_
timestamp 1698431365
transform -1 0 11088 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2490_
timestamp 1698431365
transform -1 0 24192 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2491_
timestamp 1698431365
transform 1 0 23632 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2492_
timestamp 1698431365
transform -1 0 32144 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2493_
timestamp 1698431365
transform 1 0 30800 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2494_
timestamp 1698431365
transform 1 0 29792 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2495_
timestamp 1698431365
transform 1 0 29680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2496_
timestamp 1698431365
transform -1 0 21952 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2497_
timestamp 1698431365
transform 1 0 21952 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2498_
timestamp 1698431365
transform -1 0 21952 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2499_
timestamp 1698431365
transform 1 0 19264 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2500_
timestamp 1698431365
transform -1 0 19712 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2501_
timestamp 1698431365
transform -1 0 21952 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2502_
timestamp 1698431365
transform 1 0 19600 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2503_
timestamp 1698431365
transform 1 0 21840 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2504_
timestamp 1698431365
transform 1 0 25984 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2505_
timestamp 1698431365
transform 1 0 30688 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2506_
timestamp 1698431365
transform 1 0 30352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2507_
timestamp 1698431365
transform 1 0 30128 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2508_
timestamp 1698431365
transform 1 0 30128 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2509_
timestamp 1698431365
transform 1 0 26544 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2510_
timestamp 1698431365
transform 1 0 33040 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2511_
timestamp 1698431365
transform 1 0 32928 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2512_
timestamp 1698431365
transform 1 0 34944 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2513_
timestamp 1698431365
transform 1 0 35504 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2514_
timestamp 1698431365
transform -1 0 13104 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2515_
timestamp 1698431365
transform 1 0 10864 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2516_
timestamp 1698431365
transform -1 0 10752 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2517_
timestamp 1698431365
transform 1 0 11312 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2518_
timestamp 1698431365
transform -1 0 8512 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2519_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2520_
timestamp 1698431365
transform 1 0 22960 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2521_
timestamp 1698431365
transform 1 0 28672 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2522_
timestamp 1698431365
transform -1 0 27216 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2523_
timestamp 1698431365
transform 1 0 29568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2524_
timestamp 1698431365
transform -1 0 31024 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2525_
timestamp 1698431365
transform 1 0 30352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2526_
timestamp 1698431365
transform 1 0 23856 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2527_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2528_
timestamp 1698431365
transform -1 0 32480 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2529_
timestamp 1698431365
transform 1 0 34832 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2530_
timestamp 1698431365
transform -1 0 35280 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2531_
timestamp 1698431365
transform -1 0 24864 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2532_
timestamp 1698431365
transform -1 0 24416 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2533_
timestamp 1698431365
transform 1 0 21280 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2534_
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2535_
timestamp 1698431365
transform -1 0 26320 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2536_
timestamp 1698431365
transform 1 0 22960 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2537_
timestamp 1698431365
transform 1 0 21280 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2538_
timestamp 1698431365
transform 1 0 26320 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2539_
timestamp 1698431365
transform 1 0 25984 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2540_
timestamp 1698431365
transform -1 0 26544 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2541_
timestamp 1698431365
transform 1 0 26544 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2542_
timestamp 1698431365
transform 1 0 26768 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2543_
timestamp 1698431365
transform 1 0 21504 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2544_
timestamp 1698431365
transform 1 0 21728 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2545_
timestamp 1698431365
transform 1 0 20272 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2546_
timestamp 1698431365
transform -1 0 24304 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2547_
timestamp 1698431365
transform -1 0 24976 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2548_
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2549_
timestamp 1698431365
transform 1 0 26208 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2550_
timestamp 1698431365
transform 1 0 25648 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2551_
timestamp 1698431365
transform 1 0 26544 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2552_
timestamp 1698431365
transform -1 0 28112 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2553_
timestamp 1698431365
transform 1 0 26544 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2554_
timestamp 1698431365
transform 1 0 27104 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2555_
timestamp 1698431365
transform 1 0 26656 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2556_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2557_
timestamp 1698431365
transform 1 0 28896 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2558_
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2559_
timestamp 1698431365
transform 1 0 26320 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2560_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2561_
timestamp 1698431365
transform -1 0 33600 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2562_
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2563_
timestamp 1698431365
transform 1 0 35616 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2564_
timestamp 1698431365
transform 1 0 7504 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2565_
timestamp 1698431365
transform 1 0 7056 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2566_
timestamp 1698431365
transform -1 0 6160 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2567_
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2568_
timestamp 1698431365
transform -1 0 7280 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2569_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4032 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2570_
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2571_
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2572_
timestamp 1698431365
transform 1 0 4592 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2573_
timestamp 1698431365
transform 1 0 12208 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2574_
timestamp 1698431365
transform 1 0 9520 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2575_
timestamp 1698431365
transform 1 0 13664 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2576_
timestamp 1698431365
transform 1 0 9520 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2577_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2578_
timestamp 1698431365
transform 1 0 8736 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2579_
timestamp 1698431365
transform 1 0 17360 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2580_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2581_
timestamp 1698431365
transform 1 0 12432 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2582_
timestamp 1698431365
transform 1 0 9856 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2583_
timestamp 1698431365
transform 1 0 16352 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2584_
timestamp 1698431365
transform 1 0 15456 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2585_
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2586_
timestamp 1698431365
transform 1 0 3024 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2587_
timestamp 1698431365
transform 1 0 44800 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2588_
timestamp 1698431365
transform 1 0 21616 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2589_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11760 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2590_
timestamp 1698431365
transform -1 0 12768 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2591_
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2592_
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2593_
timestamp 1698431365
transform 1 0 22960 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2594_
timestamp 1698431365
transform 1 0 10864 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2595_
timestamp 1698431365
transform -1 0 22512 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2596_
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2597_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2598_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2599_
timestamp 1698431365
transform 1 0 5936 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2600_
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2601_
timestamp 1698431365
transform 1 0 2688 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2602_
timestamp 1698431365
transform 1 0 2128 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2603_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2604_
timestamp 1698431365
transform 1 0 1904 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2605_
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2606_
timestamp 1698431365
transform 1 0 17024 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2607_
timestamp 1698431365
transform 1 0 19824 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2608_
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2609_
timestamp 1698431365
transform 1 0 13552 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2610_
timestamp 1698431365
transform 1 0 11984 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2611_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2612_
timestamp 1698431365
transform 1 0 23520 0 1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2613_
timestamp 1698431365
transform 1 0 25536 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2614_
timestamp 1698431365
transform 1 0 27328 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2615_
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2616_
timestamp 1698431365
transform 1 0 30240 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2617_
timestamp 1698431365
transform 1 0 30688 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2618_
timestamp 1698431365
transform 1 0 32256 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2619_
timestamp 1698431365
transform 1 0 34720 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2620_
timestamp 1698431365
transform -1 0 42784 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2621_
timestamp 1698431365
transform -1 0 45808 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2622_
timestamp 1698431365
transform 1 0 26992 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2623_
timestamp 1698431365
transform 1 0 41216 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2624_
timestamp 1698431365
transform -1 0 47936 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2625_
timestamp 1698431365
transform 1 0 46368 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2626_
timestamp 1698431365
transform 1 0 49280 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2627_
timestamp 1698431365
transform 1 0 50288 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2628_
timestamp 1698431365
transform 1 0 51520 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2629_
timestamp 1698431365
transform 1 0 48496 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2630_
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2631_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2632_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2633_
timestamp 1698431365
transform 1 0 39088 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2634_
timestamp 1698431365
transform 1 0 39424 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2635_
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2636_
timestamp 1698431365
transform 1 0 40992 0 1 43904
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2637_
timestamp 1698431365
transform -1 0 44016 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2638_
timestamp 1698431365
transform -1 0 47936 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2639_
timestamp 1698431365
transform 1 0 47152 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2640_
timestamp 1698431365
transform 1 0 50288 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2641_
timestamp 1698431365
transform 1 0 42896 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2642_
timestamp 1698431365
transform -1 0 54432 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2643_
timestamp 1698431365
transform -1 0 58352 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2644_
timestamp 1698431365
transform 1 0 54880 0 1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2645_
timestamp 1698431365
transform -1 0 57680 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2646_
timestamp 1698431365
transform 1 0 41216 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2647_
timestamp 1698431365
transform 1 0 54656 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2648_
timestamp 1698431365
transform 1 0 51744 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2649_
timestamp 1698431365
transform 1 0 48384 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2650_
timestamp 1698431365
transform 1 0 50064 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2651_
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2652_
timestamp 1698431365
transform -1 0 47040 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2653_
timestamp 1698431365
transform 1 0 41440 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2654_
timestamp 1698431365
transform -1 0 41664 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2655_
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2656_
timestamp 1698431365
transform -1 0 40320 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2657_
timestamp 1698431365
transform 1 0 35728 0 -1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2658_
timestamp 1698431365
transform 1 0 33040 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2659_
timestamp 1698431365
transform 1 0 29568 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2660_
timestamp 1698431365
transform 1 0 28672 0 -1 28224
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2661_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2662_
timestamp 1698431365
transform 1 0 36176 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2663_
timestamp 1698431365
transform -1 0 47936 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2664_
timestamp 1698431365
transform 1 0 33376 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2665_
timestamp 1698431365
transform 1 0 36176 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2666_
timestamp 1698431365
transform 1 0 19936 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2667_
timestamp 1698431365
transform 1 0 17696 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2668_
timestamp 1698431365
transform -1 0 30352 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2669_
timestamp 1698431365
transform 1 0 27888 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2670_
timestamp 1698431365
transform 1 0 28336 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2671_
timestamp 1698431365
transform 1 0 27440 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2672_
timestamp 1698431365
transform 1 0 31024 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2673_
timestamp 1698431365
transform 1 0 29456 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2674_
timestamp 1698431365
transform 1 0 26208 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2675_
timestamp 1698431365
transform 1 0 31584 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2676_
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2677_
timestamp 1698431365
transform 1 0 34496 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2678_
timestamp 1698431365
transform 1 0 34944 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2679_
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2680_
timestamp 1698431365
transform 1 0 34832 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2681_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2682_
timestamp 1698431365
transform 1 0 31808 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2683_
timestamp 1698431365
transform 1 0 7952 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2684_
timestamp 1698431365
transform 1 0 7728 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2685_
timestamp 1698431365
transform 1 0 7840 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2686_
timestamp 1698431365
transform 1 0 7952 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2687_
timestamp 1698431365
transform 1 0 7840 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2688_
timestamp 1698431365
transform 1 0 8288 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2689_
timestamp 1698431365
transform 1 0 9744 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2690_
timestamp 1698431365
transform 1 0 12320 0 -1 54880
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2691_
timestamp 1698431365
transform 1 0 16912 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2692_
timestamp 1698431365
transform 1 0 15232 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2693_
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2694_
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2695_
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2696_
timestamp 1698431365
transform -1 0 8960 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2697_
timestamp 1698431365
transform 1 0 5264 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2698_
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2699_
timestamp 1698431365
transform -1 0 7728 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2700_
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2701_
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2702_
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2703_
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2704_
timestamp 1698431365
transform -1 0 8736 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2705_
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2706_
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2707_
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2708_
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2709_
timestamp 1698431365
transform -1 0 28672 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2710_
timestamp 1698431365
transform 1 0 23296 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2711_
timestamp 1698431365
transform 1 0 19488 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2712_
timestamp 1698431365
transform 1 0 16240 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2713_
timestamp 1698431365
transform 1 0 15344 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2714_
timestamp 1698431365
transform -1 0 28336 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2715_
timestamp 1698431365
transform -1 0 24640 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2716_
timestamp 1698431365
transform 1 0 18032 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2717_
timestamp 1698431365
transform 1 0 12208 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2718_
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2719_
timestamp 1698431365
transform -1 0 28336 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2720_
timestamp 1698431365
transform -1 0 24080 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2721_
timestamp 1698431365
transform -1 0 25536 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2722_
timestamp 1698431365
transform -1 0 28112 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2723_
timestamp 1698431365
transform 1 0 33376 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2724_
timestamp 1698431365
transform -1 0 38528 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2725_
timestamp 1698431365
transform 1 0 15456 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2726_
timestamp 1698431365
transform 1 0 16352 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2727_
timestamp 1698431365
transform 1 0 8624 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2728_
timestamp 1698431365
transform 1 0 9408 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2729_
timestamp 1698431365
transform -1 0 33824 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2730_
timestamp 1698431365
transform -1 0 32368 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2731_
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2732_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2733_
timestamp 1698431365
transform -1 0 33936 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2734_
timestamp 1698431365
transform -1 0 32704 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2735_
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2736_
timestamp 1698431365
transform -1 0 39424 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2737_
timestamp 1698431365
transform 1 0 8064 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2738_
timestamp 1698431365
transform 1 0 6832 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2739_
timestamp 1698431365
transform 1 0 25424 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2740_
timestamp 1698431365
transform -1 0 32032 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2741_
timestamp 1698431365
transform 1 0 30912 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2742_
timestamp 1698431365
transform 1 0 34048 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2743_
timestamp 1698431365
transform 1 0 20720 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2744_
timestamp 1698431365
transform 1 0 21952 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2745_
timestamp 1698431365
transform 1 0 25200 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2746_
timestamp 1698431365
transform 1 0 26544 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2747_
timestamp 1698431365
transform 1 0 20048 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2748_
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2749_
timestamp 1698431365
transform 1 0 25536 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2750_
timestamp 1698431365
transform 1 0 25536 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2751_
timestamp 1698431365
transform -1 0 28784 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2752_
timestamp 1698431365
transform -1 0 32256 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2753_
timestamp 1698431365
transform 1 0 31584 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2754_
timestamp 1698431365
transform -1 0 38416 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2755_
timestamp 1698431365
transform 1 0 3808 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2756_
timestamp 1698431365
transform 1 0 5488 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__I asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11872 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__I
timestamp 1698431365
transform 1 0 30240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A3
timestamp 1698431365
transform -1 0 13776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1374__A1
timestamp 1698431365
transform 1 0 17024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A1
timestamp 1698431365
transform 1 0 16576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A2
timestamp 1698431365
transform -1 0 16128 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A1
timestamp 1698431365
transform 1 0 13888 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A1
timestamp 1698431365
transform 1 0 11760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__I
timestamp 1698431365
transform -1 0 17920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__I
timestamp 1698431365
transform 1 0 16576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A1
timestamp 1698431365
transform -1 0 11312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1464__I
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1476__S
timestamp 1698431365
transform 1 0 15232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A1
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__A1
timestamp 1698431365
transform 1 0 26320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__A1
timestamp 1698431365
transform 1 0 23968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__A2
timestamp 1698431365
transform 1 0 26656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__S
timestamp 1698431365
transform 1 0 15456 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__S
timestamp 1698431365
transform -1 0 16352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__A1
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__A1
timestamp 1698431365
transform 1 0 27440 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__A2
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__B
timestamp 1698431365
transform 1 0 17248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__I
timestamp 1698431365
transform 1 0 22960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__I
timestamp 1698431365
transform -1 0 46928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A1
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A1
timestamp 1698431365
transform 1 0 23072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A1
timestamp 1698431365
transform -1 0 21952 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__B
timestamp 1698431365
transform 1 0 22512 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__A1
timestamp 1698431365
transform 1 0 17472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__B
timestamp 1698431365
transform 1 0 22960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A1
timestamp 1698431365
transform -1 0 13888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__B
timestamp 1698431365
transform -1 0 14336 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__I
timestamp 1698431365
transform 1 0 27888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__I
timestamp 1698431365
transform -1 0 15680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A1
timestamp 1698431365
transform -1 0 11536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__I
timestamp 1698431365
transform 1 0 16240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__A1
timestamp 1698431365
transform -1 0 19936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__I
timestamp 1698431365
transform -1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1698431365
transform 1 0 18480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I
timestamp 1698431365
transform 1 0 17808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__I
timestamp 1698431365
transform 1 0 23744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A2
timestamp 1698431365
transform -1 0 13888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A2
timestamp 1698431365
transform -1 0 14336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A1
timestamp 1698431365
transform 1 0 19376 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__A1
timestamp 1698431365
transform 1 0 22736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__I
timestamp 1698431365
transform -1 0 17024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__A2
timestamp 1698431365
transform 1 0 19152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__I
timestamp 1698431365
transform -1 0 13776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A2
timestamp 1698431365
transform 1 0 20048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__A1
timestamp 1698431365
transform -1 0 7616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__I
timestamp 1698431365
transform 1 0 48160 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A1
timestamp 1698431365
transform 1 0 15568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A2
timestamp 1698431365
transform -1 0 16016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__I
timestamp 1698431365
transform -1 0 9072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A1
timestamp 1698431365
transform 1 0 11088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A2
timestamp 1698431365
transform 1 0 10864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__I
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1698431365
transform -1 0 7728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A2
timestamp 1698431365
transform -1 0 6160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__A1
timestamp 1698431365
transform -1 0 8512 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__A2
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__A1
timestamp 1698431365
transform 1 0 14896 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A1
timestamp 1698431365
transform 1 0 19040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A2
timestamp 1698431365
transform 1 0 20048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__C
timestamp 1698431365
transform -1 0 27440 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__I
timestamp 1698431365
transform 1 0 28112 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A1
timestamp 1698431365
transform -1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__A1
timestamp 1698431365
transform -1 0 27776 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__I
timestamp 1698431365
transform 1 0 51072 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A1
timestamp 1698431365
transform -1 0 51072 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__I
timestamp 1698431365
transform 1 0 26096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__B
timestamp 1698431365
transform 1 0 33152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__B
timestamp 1698431365
transform -1 0 35728 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__A1
timestamp 1698431365
transform 1 0 40208 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__A1
timestamp 1698431365
transform -1 0 39312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__I
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__A1
timestamp 1698431365
transform 1 0 39648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__B
timestamp 1698431365
transform 1 0 40768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__A1
timestamp 1698431365
transform 1 0 38304 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__I
timestamp 1698431365
transform 1 0 38080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A1
timestamp 1698431365
transform 1 0 46368 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__I
timestamp 1698431365
transform 1 0 43792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__B
timestamp 1698431365
transform -1 0 43568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A2
timestamp 1698431365
transform 1 0 43568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__C
timestamp 1698431365
transform -1 0 43568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__I
timestamp 1698431365
transform 1 0 43232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A2
timestamp 1698431365
transform 1 0 45920 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__B
timestamp 1698431365
transform 1 0 44240 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__A1
timestamp 1698431365
transform -1 0 47824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__I
timestamp 1698431365
transform 1 0 47152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A2
timestamp 1698431365
transform -1 0 49504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A1
timestamp 1698431365
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A1
timestamp 1698431365
transform -1 0 50960 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A1
timestamp 1698431365
transform 1 0 48832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1956__A2
timestamp 1698431365
transform 1 0 52528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__A1
timestamp 1698431365
transform 1 0 43344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A2
timestamp 1698431365
transform 1 0 43456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__C
timestamp 1698431365
transform -1 0 44464 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__I
timestamp 1698431365
transform 1 0 46816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__B
timestamp 1698431365
transform 1 0 48160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__B
timestamp 1698431365
transform -1 0 46704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A2
timestamp 1698431365
transform 1 0 51632 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__C
timestamp 1698431365
transform 1 0 52080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__A1
timestamp 1698431365
transform -1 0 57344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A2
timestamp 1698431365
transform 1 0 56672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__C
timestamp 1698431365
transform 1 0 56000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A1
timestamp 1698431365
transform 1 0 57792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A2
timestamp 1698431365
transform 1 0 56672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__C
timestamp 1698431365
transform -1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1698431365
transform 1 0 50736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__B
timestamp 1698431365
transform 1 0 48832 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__A2
timestamp 1698431365
transform -1 0 51408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__C
timestamp 1698431365
transform 1 0 50960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2027__A2
timestamp 1698431365
transform 1 0 42896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__A1
timestamp 1698431365
transform 1 0 41664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2034__B
timestamp 1698431365
transform 1 0 44800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__A2
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__C
timestamp 1698431365
transform 1 0 43792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__B2
timestamp 1698431365
transform 1 0 53200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__C
timestamp 1698431365
transform 1 0 52752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A2
timestamp 1698431365
transform 1 0 54432 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__C
timestamp 1698431365
transform 1 0 52752 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A1
timestamp 1698431365
transform 1 0 49504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2057__A1
timestamp 1698431365
transform -1 0 53088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__A2
timestamp 1698431365
transform 1 0 52080 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__C
timestamp 1698431365
transform 1 0 51632 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__B
timestamp 1698431365
transform 1 0 51184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__B
timestamp 1698431365
transform 1 0 46928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2066__C
timestamp 1698431365
transform -1 0 41888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__A2
timestamp 1698431365
transform -1 0 48384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__B
timestamp 1698431365
transform 1 0 48832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__A1
timestamp 1698431365
transform -1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__A1
timestamp 1698431365
transform 1 0 45696 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__B
timestamp 1698431365
transform -1 0 43680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2093__A2
timestamp 1698431365
transform -1 0 42784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2094__A1
timestamp 1698431365
transform 1 0 40992 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__B
timestamp 1698431365
transform -1 0 45920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__A2
timestamp 1698431365
transform 1 0 42784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__C
timestamp 1698431365
transform -1 0 41216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2109__A1
timestamp 1698431365
transform 1 0 39088 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A2
timestamp 1698431365
transform 1 0 39984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__B
timestamp 1698431365
transform 1 0 40432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__A1
timestamp 1698431365
transform -1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__C
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__C
timestamp 1698431365
transform -1 0 35392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A2
timestamp 1698431365
transform -1 0 37072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__A1
timestamp 1698431365
transform -1 0 34048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2133__C
timestamp 1698431365
transform 1 0 31584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__C
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__A2
timestamp 1698431365
transform 1 0 34496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__C
timestamp 1698431365
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2148__A1
timestamp 1698431365
transform 1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__A1
timestamp 1698431365
transform -1 0 46928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__A2
timestamp 1698431365
transform 1 0 45808 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A1
timestamp 1698431365
transform 1 0 45360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A2
timestamp 1698431365
transform -1 0 47376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A1
timestamp 1698431365
transform 1 0 35392 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__A1
timestamp 1698431365
transform 1 0 33936 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__A2
timestamp 1698431365
transform 1 0 20160 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2159__A2
timestamp 1698431365
transform -1 0 17808 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2160__I
timestamp 1698431365
transform 1 0 25312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A3
timestamp 1698431365
transform 1 0 19152 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2167__B
timestamp 1698431365
transform -1 0 30128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A1
timestamp 1698431365
transform 1 0 27216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A2
timestamp 1698431365
transform -1 0 27328 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__B2
timestamp 1698431365
transform -1 0 26880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2211__A1
timestamp 1698431365
transform -1 0 25200 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__B2
timestamp 1698431365
transform 1 0 28000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__I
timestamp 1698431365
transform -1 0 26096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__I
timestamp 1698431365
transform 1 0 26432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__B
timestamp 1698431365
transform 1 0 31920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__A1
timestamp 1698431365
transform 1 0 24528 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A1
timestamp 1698431365
transform 1 0 28672 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2268__B
timestamp 1698431365
transform 1 0 33376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__A1
timestamp 1698431365
transform 1 0 24080 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2278__B
timestamp 1698431365
transform -1 0 38192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2285__I
timestamp 1698431365
transform 1 0 34160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2286__B
timestamp 1698431365
transform 1 0 36624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1698431365
transform 1 0 27552 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__B2
timestamp 1698431365
transform 1 0 31360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A1
timestamp 1698431365
transform 1 0 32592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2316__A1
timestamp 1698431365
transform -1 0 10976 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__A1
timestamp 1698431365
transform 1 0 12208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__C
timestamp 1698431365
transform -1 0 14896 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__A1
timestamp 1698431365
transform 1 0 15456 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A1
timestamp 1698431365
transform -1 0 16240 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A2
timestamp 1698431365
transform 1 0 17472 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__A1
timestamp 1698431365
transform 1 0 11760 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2332__A1
timestamp 1698431365
transform 1 0 15904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2337__B
timestamp 1698431365
transform 1 0 15904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2338__A1
timestamp 1698431365
transform 1 0 11648 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__A2
timestamp 1698431365
transform 1 0 15456 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__B
timestamp 1698431365
transform -1 0 16576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2357__B
timestamp 1698431365
transform 1 0 21392 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A1
timestamp 1698431365
transform -1 0 9968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__B
timestamp 1698431365
transform 1 0 23072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__A1
timestamp 1698431365
transform 1 0 25312 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2429__A1
timestamp 1698431365
transform 1 0 22736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__C
timestamp 1698431365
transform 1 0 25424 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2458__A1
timestamp 1698431365
transform 1 0 25312 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__A1
timestamp 1698431365
transform 1 0 24976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A1
timestamp 1698431365
transform 1 0 25984 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__I
timestamp 1698431365
transform 1 0 29568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2472__A1
timestamp 1698431365
transform 1 0 23744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2475__I
timestamp 1698431365
transform 1 0 29232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2478__I
timestamp 1698431365
transform 1 0 16128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A2
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__I
timestamp 1698431365
transform -1 0 19488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__A1
timestamp 1698431365
transform -1 0 13552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__A2
timestamp 1698431365
transform 1 0 23408 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A1
timestamp 1698431365
transform 1 0 21952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A1
timestamp 1698431365
transform 1 0 24640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2509__A1
timestamp 1698431365
transform 1 0 27888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2509__A2
timestamp 1698431365
transform 1 0 26320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__A1
timestamp 1698431365
transform -1 0 13552 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__I
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A1
timestamp 1698431365
transform 1 0 23744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2523__I
timestamp 1698431365
transform 1 0 30464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__A1
timestamp 1698431365
transform 1 0 24192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__I
timestamp 1698431365
transform -1 0 25088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A1
timestamp 1698431365
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A2
timestamp 1698431365
transform 1 0 24864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__I
timestamp 1698431365
transform -1 0 25648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A1
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A2
timestamp 1698431365
transform 1 0 25984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__A1
timestamp 1698431365
transform -1 0 22848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__A2
timestamp 1698431365
transform 1 0 21280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A1
timestamp 1698431365
transform 1 0 25424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__A1
timestamp 1698431365
transform 1 0 26320 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__I
timestamp 1698431365
transform 1 0 27216 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__A1
timestamp 1698431365
transform 1 0 26768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2564__A1
timestamp 1698431365
transform 1 0 9184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2569__CLK
timestamp 1698431365
transform -1 0 7504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2570__CLK
timestamp 1698431365
transform 1 0 10080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__CLK
timestamp 1698431365
transform 1 0 8064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__CLK
timestamp 1698431365
transform 1 0 15680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2574__CLK
timestamp 1698431365
transform 1 0 12992 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__CLK
timestamp 1698431365
transform 1 0 12544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__CLK
timestamp 1698431365
transform 1 0 12880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__CLK
timestamp 1698431365
transform 1 0 12208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__CLK
timestamp 1698431365
transform 1 0 21616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__CLK
timestamp 1698431365
transform 1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__CLK
timestamp 1698431365
transform 1 0 12208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__CLK
timestamp 1698431365
transform 1 0 13552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__CLK
timestamp 1698431365
transform 1 0 19824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__CLK
timestamp 1698431365
transform 1 0 18928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__CLK
timestamp 1698431365
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__CLK
timestamp 1698431365
transform -1 0 6496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__CLK
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__CLK
timestamp 1698431365
transform -1 0 15120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__CLK
timestamp 1698431365
transform 1 0 12768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__CLK
timestamp 1698431365
transform -1 0 18816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__CLK
timestamp 1698431365
transform 1 0 23184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__CLK
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__CLK
timestamp 1698431365
transform -1 0 15680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__CLK
timestamp 1698431365
transform 1 0 13104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__CLK
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2598__CLK
timestamp 1698431365
transform 1 0 8960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2599__CLK
timestamp 1698431365
transform 1 0 9184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__CLK
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2601__CLK
timestamp 1698431365
transform 1 0 5936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2602__CLK
timestamp 1698431365
transform 1 0 5712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2603__CLK
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__CLK
timestamp 1698431365
transform -1 0 5376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__CLK
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2606__CLK
timestamp 1698431365
transform 1 0 20496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__CLK
timestamp 1698431365
transform 1 0 23296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__CLK
timestamp 1698431365
transform 1 0 23072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__CLK
timestamp 1698431365
transform 1 0 16800 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__CLK
timestamp 1698431365
transform 1 0 23296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__CLK
timestamp 1698431365
transform 1 0 29680 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__CLK
timestamp 1698431365
transform 1 0 30800 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__CLK
timestamp 1698431365
transform 1 0 33712 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__CLK
timestamp 1698431365
transform 1 0 34160 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__CLK
timestamp 1698431365
transform 1 0 32032 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__CLK
timestamp 1698431365
transform 1 0 34496 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__CLK
timestamp 1698431365
transform 1 0 30464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__CLK
timestamp 1698431365
transform 1 0 44912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__CLK
timestamp 1698431365
transform 1 0 49840 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__CLK
timestamp 1698431365
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__CLK
timestamp 1698431365
transform 1 0 51408 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__CLK
timestamp 1698431365
transform -1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__CLK
timestamp 1698431365
transform 1 0 40320 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__CLK
timestamp 1698431365
transform 1 0 42560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__CLK
timestamp 1698431365
transform 1 0 42896 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__CLK
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2636__CLK
timestamp 1698431365
transform 1 0 44464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__CLK
timestamp 1698431365
transform -1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__CLK
timestamp 1698431365
transform 1 0 48160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__CLK
timestamp 1698431365
transform 1 0 46256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__CLK
timestamp 1698431365
transform -1 0 50288 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__CLK
timestamp 1698431365
transform 1 0 46368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__CLK
timestamp 1698431365
transform -1 0 51184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2643__CLK
timestamp 1698431365
transform 1 0 54880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__CLK
timestamp 1698431365
transform 1 0 55552 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__CLK
timestamp 1698431365
transform 1 0 55328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__CLK
timestamp 1698431365
transform 1 0 44912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__CLK
timestamp 1698431365
transform 1 0 54432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__CLK
timestamp 1698431365
transform 1 0 53648 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__CLK
timestamp 1698431365
transform 1 0 48160 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2650__CLK
timestamp 1698431365
transform 1 0 49840 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__CLK
timestamp 1698431365
transform 1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__CLK
timestamp 1698431365
transform -1 0 47264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2653__CLK
timestamp 1698431365
transform -1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2654__CLK
timestamp 1698431365
transform 1 0 41888 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__CLK
timestamp 1698431365
transform 1 0 42112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2656__CLK
timestamp 1698431365
transform 1 0 41888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2657__CLK
timestamp 1698431365
transform 1 0 35504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2658__CLK
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2659__CLK
timestamp 1698431365
transform 1 0 29344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__CLK
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__CLK
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__CLK
timestamp 1698431365
transform 1 0 40208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__CLK
timestamp 1698431365
transform 1 0 48160 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2664__CLK
timestamp 1698431365
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2665__CLK
timestamp 1698431365
transform 1 0 35728 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2665__D
timestamp 1698431365
transform -1 0 35504 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2666__CLK
timestamp 1698431365
transform 1 0 19712 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__CLK
timestamp 1698431365
transform 1 0 16800 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__CLK
timestamp 1698431365
transform 1 0 30352 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__CLK
timestamp 1698431365
transform 1 0 27664 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2670__CLK
timestamp 1698431365
transform 1 0 31808 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__CLK
timestamp 1698431365
transform 1 0 30688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__CLK
timestamp 1698431365
transform -1 0 34048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__CLK
timestamp 1698431365
transform 1 0 32704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2674__CLK
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2675__CLK
timestamp 1698431365
transform 1 0 35056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__CLK
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2677__CLK
timestamp 1698431365
transform 1 0 37744 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__CLK
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__CLK
timestamp 1698431365
transform 1 0 38976 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__CLK
timestamp 1698431365
transform 1 0 37072 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__CLK
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__CLK
timestamp 1698431365
transform 1 0 7728 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__CLK
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__CLK
timestamp 1698431365
transform 1 0 7616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2686__CLK
timestamp 1698431365
transform 1 0 7728 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__CLK
timestamp 1698431365
transform 1 0 7952 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__CLK
timestamp 1698431365
transform 1 0 8064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__CLK
timestamp 1698431365
transform 1 0 9520 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__CLK
timestamp 1698431365
transform 1 0 12096 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__CLK
timestamp 1698431365
transform 1 0 20944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__CLK
timestamp 1698431365
transform 1 0 18704 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__CLK
timestamp 1698431365
transform 1 0 5040 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__CLK
timestamp 1698431365
transform 1 0 5040 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__CLK
timestamp 1698431365
transform 1 0 5040 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__CLK
timestamp 1698431365
transform 1 0 9184 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__CLK
timestamp 1698431365
transform 1 0 8736 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__CLK
timestamp 1698431365
transform 1 0 8400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__CLK
timestamp 1698431365
transform 1 0 9520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__CLK
timestamp 1698431365
transform 1 0 9184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__CLK
timestamp 1698431365
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__CLK
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__CLK
timestamp 1698431365
transform 1 0 8736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__CLK
timestamp 1698431365
transform 1 0 5040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__CLK
timestamp 1698431365
transform -1 0 4816 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__CLK
timestamp 1698431365
transform 1 0 5040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__CLK
timestamp 1698431365
transform 1 0 5040 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__CLK
timestamp 1698431365
transform 1 0 22960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__CLK
timestamp 1698431365
transform 1 0 22624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__CLK
timestamp 1698431365
transform -1 0 22960 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__CLK
timestamp 1698431365
transform -1 0 19712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__CLK
timestamp 1698431365
transform 1 0 18592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2715__CLK
timestamp 1698431365
transform 1 0 21840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__CLK
timestamp 1698431365
transform 1 0 21392 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2718__CLK
timestamp 1698431365
transform 1 0 16800 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2719__CLK
timestamp 1698431365
transform 1 0 28336 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2720__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2721__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2722__CLK
timestamp 1698431365
transform 1 0 28336 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2723__CLK
timestamp 1698431365
transform 1 0 36848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__CLK
timestamp 1698431365
transform 1 0 38752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__CLK
timestamp 1698431365
transform 1 0 17808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__CLK
timestamp 1698431365
transform 1 0 19712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__CLK
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2728__CLK
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2729__CLK
timestamp 1698431365
transform -1 0 34272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__CLK
timestamp 1698431365
transform -1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__CLK
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__CLK
timestamp 1698431365
transform 1 0 33376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__CLK
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__CLK
timestamp 1698431365
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__CLK
timestamp 1698431365
transform 1 0 39648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__CLK
timestamp 1698431365
transform 1 0 11760 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2738__CLK
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2739__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2740__CLK
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__CLK
timestamp 1698431365
transform 1 0 30688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2742__CLK
timestamp 1698431365
transform 1 0 37520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__CLK
timestamp 1698431365
transform 1 0 24192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__CLK
timestamp 1698431365
transform 1 0 25648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2747__CLK
timestamp 1698431365
transform 1 0 22176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2748__CLK
timestamp 1698431365
transform 1 0 25200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2749__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2750__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2751__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2752__CLK
timestamp 1698431365
transform 1 0 32480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2753__CLK
timestamp 1698431365
transform 1 0 34832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2754__CLK
timestamp 1698431365
transform 1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2755__CLK
timestamp 1698431365
transform 1 0 7056 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2756__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 29680 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 12544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 8624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 26432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 9632 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 9072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 21280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 20160 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 44016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 43344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 36176 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 31808 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 45024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 44576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 20160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 20048 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 40208 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 14896 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 15344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 4704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output11_I
timestamp 1698431365
transform 1 0 29904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30016 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_wb_clk_i asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1698431365
transform 1 0 6272 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1698431365
transform 1 0 21056 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1698431365
transform 1 0 21952 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1698431365
transform -1 0 8960 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1698431365
transform 1 0 6160 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1698431365
transform 1 0 15120 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1698431365
transform 1 0 37296 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1698431365
transform 1 0 32928 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1698431365
transform 1 0 45584 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1698431365
transform 1 0 44688 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1698431365
transform 1 0 33040 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1698431365
transform -1 0 32704 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1698431365
transform 1 0 45024 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1698431365
transform 1 0 45248 0 -1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_206 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_214 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25312 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_218 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_235
timestamp 1698431365
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698431365
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_88
timestamp 1698431365
transform 1 0 11200 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_96
timestamp 1698431365
transform 1 0 12096 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_128
timestamp 1698431365
transform 1 0 15680 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_158
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_166
timestamp 1698431365
transform 1 0 19936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_170
timestamp 1698431365
transform 1 0 20384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_172
timestamp 1698431365
transform 1 0 20608 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_202
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_254
timestamp 1698431365
transform 1 0 29792 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698431365
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698431365
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_123
timestamp 1698431365
transform 1 0 15120 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_131
timestamp 1698431365
transform 1 0 16016 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_163
timestamp 1698431365
transform 1 0 19600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_167
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_80
timestamp 1698431365
transform 1 0 10304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_84
timestamp 1698431365
transform 1 0 10752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_86
timestamp 1698431365
transform 1 0 10976 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_93
timestamp 1698431365
transform 1 0 11760 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_101
timestamp 1698431365
transform 1 0 12656 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_105
timestamp 1698431365
transform 1 0 13104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_113
timestamp 1698431365
transform 1 0 14000 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_117
timestamp 1698431365
transform 1 0 14448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_158
timestamp 1698431365
transform 1 0 19040 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_174
timestamp 1698431365
transform 1 0 20832 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_208
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_216
timestamp 1698431365
transform 1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_220
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_240
timestamp 1698431365
transform 1 0 28224 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_272
timestamp 1698431365
transform 1 0 31808 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_73
timestamp 1698431365
transform 1 0 9520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_75
timestamp 1698431365
transform 1 0 9744 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_155
timestamp 1698431365
transform 1 0 18704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_159
timestamp 1698431365
transform 1 0 19152 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_188
timestamp 1698431365
transform 1 0 22400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_192
timestamp 1698431365
transform 1 0 22848 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_208
timestamp 1698431365
transform 1 0 24640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_212
timestamp 1698431365
transform 1 0 25088 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_220
timestamp 1698431365
transform 1 0 25984 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_224
timestamp 1698431365
transform 1 0 26432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_226
timestamp 1698431365
transform 1 0 26656 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_233
timestamp 1698431365
transform 1 0 27440 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_88
timestamp 1698431365
transform 1 0 11200 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_92
timestamp 1698431365
transform 1 0 11648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_94
timestamp 1698431365
transform 1 0 11872 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_110
timestamp 1698431365
transform 1 0 13664 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_126
timestamp 1698431365
transform 1 0 15456 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_157
timestamp 1698431365
transform 1 0 18928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_161
timestamp 1698431365
transform 1 0 19376 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_165
timestamp 1698431365
transform 1 0 19824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_224
timestamp 1698431365
transform 1 0 26432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_240
timestamp 1698431365
transform 1 0 28224 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_272
timestamp 1698431365
transform 1 0 31808 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_72
timestamp 1698431365
transform 1 0 9408 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_76
timestamp 1698431365
transform 1 0 9856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_78
timestamp 1698431365
transform 1 0 10080 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_85
timestamp 1698431365
transform 1 0 10864 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_122
timestamp 1698431365
transform 1 0 15008 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_138
timestamp 1698431365
transform 1 0 16800 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_142
timestamp 1698431365
transform 1 0 17248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_144
timestamp 1698431365
transform 1 0 17472 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_165
timestamp 1698431365
transform 1 0 19824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_179
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_211
timestamp 1698431365
transform 1 0 24976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_215
timestamp 1698431365
transform 1 0 25424 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_259
timestamp 1698431365
transform 1 0 30352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_290
timestamp 1698431365
transform 1 0 33824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_294
timestamp 1698431365
transform 1 0 34272 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_310
timestamp 1698431365
transform 1 0 36064 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_489
timestamp 1698431365
transform 1 0 56112 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_505
timestamp 1698431365
transform 1 0 57904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_38
timestamp 1698431365
transform 1 0 5600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_40
timestamp 1698431365
transform 1 0 5824 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_107
timestamp 1698431365
transform 1 0 13328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_111
timestamp 1698431365
transform 1 0 13776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_113
timestamp 1698431365
transform 1 0 14000 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_129
timestamp 1698431365
transform 1 0 15792 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_165
timestamp 1698431365
transform 1 0 19824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_169
timestamp 1698431365
transform 1 0 20272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_173
timestamp 1698431365
transform 1 0 20720 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_177
timestamp 1698431365
transform 1 0 21168 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_180
timestamp 1698431365
transform 1 0 21504 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_214
timestamp 1698431365
transform 1 0 25312 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_239
timestamp 1698431365
transform 1 0 28112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_245
timestamp 1698431365
transform 1 0 28784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_247
timestamp 1698431365
transform 1 0 29008 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_277
timestamp 1698431365
transform 1 0 32368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_286
timestamp 1698431365
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_66
timestamp 1698431365
transform 1 0 8736 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_82
timestamp 1698431365
transform 1 0 10528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_136
timestamp 1698431365
transform 1 0 16576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_181
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_197
timestamp 1698431365
transform 1 0 23408 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_205
timestamp 1698431365
transform 1 0 24304 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_209
timestamp 1698431365
transform 1 0 24752 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_212
timestamp 1698431365
transform 1 0 25088 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_218
timestamp 1698431365
transform 1 0 25760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_237
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_251
timestamp 1698431365
transform 1 0 29456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_259
timestamp 1698431365
transform 1 0 30352 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_269
timestamp 1698431365
transform 1 0 31472 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_301
timestamp 1698431365
transform 1 0 35056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_309
timestamp 1698431365
transform 1 0 35952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698431365
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698431365
transform 1 0 56112 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_505
timestamp 1698431365
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_42
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_64
timestamp 1698431365
transform 1 0 8512 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_103
timestamp 1698431365
transform 1 0 12880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_107
timestamp 1698431365
transform 1 0 13328 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_111
timestamp 1698431365
transform 1 0 13776 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_118
timestamp 1698431365
transform 1 0 14560 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_128
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_194
timestamp 1698431365
transform 1 0 23072 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_198
timestamp 1698431365
transform 1 0 23520 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_202
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_245
timestamp 1698431365
transform 1 0 28784 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_249
timestamp 1698431365
transform 1 0 29232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_251
timestamp 1698431365
transform 1 0 29456 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_275
timestamp 1698431365
transform 1 0 32144 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_298
timestamp 1698431365
transform 1 0 34720 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_302
timestamp 1698431365
transform 1 0 35168 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_304
timestamp 1698431365
transform 1 0 35392 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_311
timestamp 1698431365
transform 1 0 36176 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_343
timestamp 1698431365
transform 1 0 39760 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_347
timestamp 1698431365
transform 1 0 40208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698431365
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_18
timestamp 1698431365
transform 1 0 3360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_26
timestamp 1698431365
transform 1 0 4256 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_30
timestamp 1698431365
transform 1 0 4704 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_33
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_66
timestamp 1698431365
transform 1 0 8736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_70
timestamp 1698431365
transform 1 0 9184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_155
timestamp 1698431365
transform 1 0 18704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_157
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_193
timestamp 1698431365
transform 1 0 22960 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_209
timestamp 1698431365
transform 1 0 24752 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_213
timestamp 1698431365
transform 1 0 25200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_237
timestamp 1698431365
transform 1 0 27888 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_269
timestamp 1698431365
transform 1 0 31472 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_277
timestamp 1698431365
transform 1 0 32368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_281
timestamp 1698431365
transform 1 0 32816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_298
timestamp 1698431365
transform 1 0 34720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_321
timestamp 1698431365
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_489
timestamp 1698431365
transform 1 0 56112 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698431365
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_46
timestamp 1698431365
transform 1 0 6496 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_62
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_74
timestamp 1698431365
transform 1 0 9632 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_87
timestamp 1698431365
transform 1 0 11088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_95
timestamp 1698431365
transform 1 0 11984 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_111
timestamp 1698431365
transform 1 0 13776 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_127
timestamp 1698431365
transform 1 0 15568 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_131
timestamp 1698431365
transform 1 0 16016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_133
timestamp 1698431365
transform 1 0 16240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_162
timestamp 1698431365
transform 1 0 19488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_166
timestamp 1698431365
transform 1 0 19936 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_174
timestamp 1698431365
transform 1 0 20832 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_178
timestamp 1698431365
transform 1 0 21280 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_183
timestamp 1698431365
transform 1 0 21840 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_222
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_235
timestamp 1698431365
transform 1 0 27664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_239
timestamp 1698431365
transform 1 0 28112 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_247
timestamp 1698431365
transform 1 0 29008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_257
timestamp 1698431365
transform 1 0 30128 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_273
timestamp 1698431365
transform 1 0 31920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_277
timestamp 1698431365
transform 1 0 32368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_340
timestamp 1698431365
transform 1 0 39424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_344
timestamp 1698431365
transform 1 0 39872 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_4
timestamp 1698431365
transform 1 0 1792 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_52
timestamp 1698431365
transform 1 0 7168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_60
timestamp 1698431365
transform 1 0 8064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_62
timestamp 1698431365
transform 1 0 8288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_94
timestamp 1698431365
transform 1 0 11872 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_100
timestamp 1698431365
transform 1 0 12544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_122
timestamp 1698431365
transform 1 0 15008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_130
timestamp 1698431365
transform 1 0 15904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698431365
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_272
timestamp 1698431365
transform 1 0 31808 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_288
timestamp 1698431365
transform 1 0 33600 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_296
timestamp 1698431365
transform 1 0 34496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698431365
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_489
timestamp 1698431365
transform 1 0 56112 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_505
timestamp 1698431365
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_10
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_26
timestamp 1698431365
transform 1 0 4256 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_36
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_40
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_56
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_64
timestamp 1698431365
transform 1 0 8512 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_98
timestamp 1698431365
transform 1 0 12320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_105
timestamp 1698431365
transform 1 0 13104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_124
timestamp 1698431365
transform 1 0 15232 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_128
timestamp 1698431365
transform 1 0 15680 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_131
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_148
timestamp 1698431365
transform 1 0 17920 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_164
timestamp 1698431365
transform 1 0 19712 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_168
timestamp 1698431365
transform 1 0 20160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_202
timestamp 1698431365
transform 1 0 23968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_218
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_239
timestamp 1698431365
transform 1 0 28112 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_247
timestamp 1698431365
transform 1 0 29008 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_297
timestamp 1698431365
transform 1 0 34608 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_329
timestamp 1698431365
transform 1 0 38192 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_345
timestamp 1698431365
transform 1 0 39984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_20
timestamp 1698431365
transform 1 0 3584 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_27
timestamp 1698431365
transform 1 0 4368 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_43
timestamp 1698431365
transform 1 0 6160 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_47
timestamp 1698431365
transform 1 0 6608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_88
timestamp 1698431365
transform 1 0 11200 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_116
timestamp 1698431365
transform 1 0 14336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_118
timestamp 1698431365
transform 1 0 14560 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_127
timestamp 1698431365
transform 1 0 15568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_143
timestamp 1698431365
transform 1 0 17360 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_206
timestamp 1698431365
transform 1 0 24416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_218
timestamp 1698431365
transform 1 0 25760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_263
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_295
timestamp 1698431365
transform 1 0 34384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_489
timestamp 1698431365
transform 1 0 56112 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_505
timestamp 1698431365
transform 1 0 57904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_10
timestamp 1698431365
transform 1 0 2464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_41
timestamp 1698431365
transform 1 0 5936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_43
timestamp 1698431365
transform 1 0 6160 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_83
timestamp 1698431365
transform 1 0 10640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_105
timestamp 1698431365
transform 1 0 13104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_109
timestamp 1698431365
transform 1 0 13552 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_119
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_123
timestamp 1698431365
transform 1 0 15120 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_129
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_148
timestamp 1698431365
transform 1 0 17920 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_156
timestamp 1698431365
transform 1 0 18816 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_162
timestamp 1698431365
transform 1 0 19488 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_184
timestamp 1698431365
transform 1 0 21952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_192
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_194
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_201
timestamp 1698431365
transform 1 0 23856 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_245
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_261
timestamp 1698431365
transform 1 0 30576 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_332
timestamp 1698431365
transform 1 0 38528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_336
timestamp 1698431365
transform 1 0 38976 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_344
timestamp 1698431365
transform 1 0 39872 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_348
timestamp 1698431365
transform 1 0 40320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_52
timestamp 1698431365
transform 1 0 7168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_59
timestamp 1698431365
transform 1 0 7952 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_139
timestamp 1698431365
transform 1 0 16912 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_146
timestamp 1698431365
transform 1 0 17696 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_153
timestamp 1698431365
transform 1 0 18480 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_181
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_183
timestamp 1698431365
transform 1 0 21840 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_186
timestamp 1698431365
transform 1 0 22176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_216
timestamp 1698431365
transform 1 0 25536 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_489
timestamp 1698431365
transform 1 0 56112 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_505
timestamp 1698431365
transform 1 0 57904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_6
timestamp 1698431365
transform 1 0 2016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_30
timestamp 1698431365
transform 1 0 4704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_38
timestamp 1698431365
transform 1 0 5600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_40
timestamp 1698431365
transform 1 0 5824 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_51
timestamp 1698431365
transform 1 0 7056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_65
timestamp 1698431365
transform 1 0 8624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_78
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_82
timestamp 1698431365
transform 1 0 10528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_84
timestamp 1698431365
transform 1 0 10752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_91
timestamp 1698431365
transform 1 0 11536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_95
timestamp 1698431365
transform 1 0 11984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_99
timestamp 1698431365
transform 1 0 12432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_111
timestamp 1698431365
transform 1 0 13776 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_113
timestamp 1698431365
transform 1 0 14000 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_148
timestamp 1698431365
transform 1 0 17920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_222
timestamp 1698431365
transform 1 0 26208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_246
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_254
timestamp 1698431365
transform 1 0 29792 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_258
timestamp 1698431365
transform 1 0 30240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_315
timestamp 1698431365
transform 1 0 36624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_319
timestamp 1698431365
transform 1 0 37072 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_335
timestamp 1698431365
transform 1 0 38864 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_343
timestamp 1698431365
transform 1 0 39760 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_347
timestamp 1698431365
transform 1 0 40208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_52
timestamp 1698431365
transform 1 0 7168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_54
timestamp 1698431365
transform 1 0 7392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_85
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_89
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_93
timestamp 1698431365
transform 1 0 11760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_111
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_130
timestamp 1698431365
transform 1 0 15904 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_134
timestamp 1698431365
transform 1 0 16352 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_150
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_164
timestamp 1698431365
transform 1 0 19712 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698431365
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_193
timestamp 1698431365
transform 1 0 22960 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_221
timestamp 1698431365
transform 1 0 26096 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_239
timestamp 1698431365
transform 1 0 28112 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_259
timestamp 1698431365
transform 1 0 30352 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_275
timestamp 1698431365
transform 1 0 32144 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_283
timestamp 1698431365
transform 1 0 33040 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_287
timestamp 1698431365
transform 1 0 33488 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_294
timestamp 1698431365
transform 1 0 34272 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_302
timestamp 1698431365
transform 1 0 35168 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698431365
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_489
timestamp 1698431365
transform 1 0 56112 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_505
timestamp 1698431365
transform 1 0 57904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_6
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_51
timestamp 1698431365
transform 1 0 7056 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_59
timestamp 1698431365
transform 1 0 7952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_61
timestamp 1698431365
transform 1 0 8176 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_82
timestamp 1698431365
transform 1 0 10528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_84
timestamp 1698431365
transform 1 0 10752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_95
timestamp 1698431365
transform 1 0 11984 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_116
timestamp 1698431365
transform 1 0 14336 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_124
timestamp 1698431365
transform 1 0 15232 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_154
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_170
timestamp 1698431365
transform 1 0 20384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_172
timestamp 1698431365
transform 1 0 20608 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_179
timestamp 1698431365
transform 1 0 21392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_199
timestamp 1698431365
transform 1 0 23632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_218
timestamp 1698431365
transform 1 0 25760 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_222
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_225
timestamp 1698431365
transform 1 0 26544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_229
timestamp 1698431365
transform 1 0 26992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_239
timestamp 1698431365
transform 1 0 28112 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_243
timestamp 1698431365
transform 1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_274
timestamp 1698431365
transform 1 0 32032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698431365
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_297
timestamp 1698431365
transform 1 0 34608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_301
timestamp 1698431365
transform 1 0 35056 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_331
timestamp 1698431365
transform 1 0 38416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_335
timestamp 1698431365
transform 1 0 38864 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_343
timestamp 1698431365
transform 1 0 39760 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_347
timestamp 1698431365
transform 1 0 40208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698431365
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_6
timestamp 1698431365
transform 1 0 2016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_15
timestamp 1698431365
transform 1 0 3024 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_22
timestamp 1698431365
transform 1 0 3808 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_30
timestamp 1698431365
transform 1 0 4704 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_41
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_43
timestamp 1698431365
transform 1 0 6160 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_64
timestamp 1698431365
transform 1 0 8512 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_66
timestamp 1698431365
transform 1 0 8736 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698431365
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_85
timestamp 1698431365
transform 1 0 10864 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_96
timestamp 1698431365
transform 1 0 12096 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_115
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_124
timestamp 1698431365
transform 1 0 15232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_140
timestamp 1698431365
transform 1 0 17024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_142
timestamp 1698431365
transform 1 0 17248 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_206
timestamp 1698431365
transform 1 0 24416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_240
timestamp 1698431365
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_249
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_265
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_269
timestamp 1698431365
transform 1 0 31472 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_299
timestamp 1698431365
transform 1 0 34832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698431365
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_357
timestamp 1698431365
transform 1 0 41328 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_373
timestamp 1698431365
transform 1 0 43120 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_381
timestamp 1698431365
transform 1 0 44016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698431365
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_489
timestamp 1698431365
transform 1 0 56112 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_505
timestamp 1698431365
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_18
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_26
timestamp 1698431365
transform 1 0 4256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_28
timestamp 1698431365
transform 1 0 4480 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_58
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_62
timestamp 1698431365
transform 1 0 8288 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698431365
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_78
timestamp 1698431365
transform 1 0 10080 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_86
timestamp 1698431365
transform 1 0 10976 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_96
timestamp 1698431365
transform 1 0 12096 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_112
timestamp 1698431365
transform 1 0 13888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_114
timestamp 1698431365
transform 1 0 14112 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_146
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_149
timestamp 1698431365
transform 1 0 18032 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_171
timestamp 1698431365
transform 1 0 20496 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_198
timestamp 1698431365
transform 1 0 23520 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_202
timestamp 1698431365
transform 1 0 23968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_265
timestamp 1698431365
transform 1 0 31024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_288
timestamp 1698431365
transform 1 0 33600 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_356
timestamp 1698431365
transform 1 0 41216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_362
timestamp 1698431365
transform 1 0 41888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_366
timestamp 1698431365
transform 1 0 42336 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_382
timestamp 1698431365
transform 1 0 44128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_390
timestamp 1698431365
transform 1 0 45024 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_394
timestamp 1698431365
transform 1 0 45472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_398
timestamp 1698431365
transform 1 0 45920 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_406
timestamp 1698431365
transform 1 0 46816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_410
timestamp 1698431365
transform 1 0 47264 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_418
timestamp 1698431365
transform 1 0 48160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_6
timestamp 1698431365
transform 1 0 2016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_14
timestamp 1698431365
transform 1 0 2912 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_18
timestamp 1698431365
transform 1 0 3360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_43
timestamp 1698431365
transform 1 0 6160 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_51
timestamp 1698431365
transform 1 0 7056 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_71
timestamp 1698431365
transform 1 0 9296 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_129
timestamp 1698431365
transform 1 0 15792 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_137
timestamp 1698431365
transform 1 0 16688 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_161
timestamp 1698431365
transform 1 0 19376 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698431365
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_189
timestamp 1698431365
transform 1 0 22512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_198
timestamp 1698431365
transform 1 0 23520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_202
timestamp 1698431365
transform 1 0 23968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_219
timestamp 1698431365
transform 1 0 25872 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_231
timestamp 1698431365
transform 1 0 27216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_235
timestamp 1698431365
transform 1 0 27664 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_253
timestamp 1698431365
transform 1 0 29680 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_261
timestamp 1698431365
transform 1 0 30576 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_293
timestamp 1698431365
transform 1 0 34160 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_297
timestamp 1698431365
transform 1 0 34608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_368
timestamp 1698431365
transform 1 0 42560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_372
timestamp 1698431365
transform 1 0 43008 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_376
timestamp 1698431365
transform 1 0 43456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_378
timestamp 1698431365
transform 1 0 43680 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_416
timestamp 1698431365
transform 1 0 47936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_420
timestamp 1698431365
transform 1 0 48384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_424
timestamp 1698431365
transform 1 0 48832 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_432
timestamp 1698431365
transform 1 0 49728 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_435
timestamp 1698431365
transform 1 0 50064 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_489
timestamp 1698431365
transform 1 0 56112 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_505
timestamp 1698431365
transform 1 0 57904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_31
timestamp 1698431365
transform 1 0 4816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_35
timestamp 1698431365
transform 1 0 5264 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_51
timestamp 1698431365
transform 1 0 7056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_53
timestamp 1698431365
transform 1 0 7280 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_82
timestamp 1698431365
transform 1 0 10528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_90
timestamp 1698431365
transform 1 0 11424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_122
timestamp 1698431365
transform 1 0 15008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_126
timestamp 1698431365
transform 1 0 15456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_130
timestamp 1698431365
transform 1 0 15904 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_146
timestamp 1698431365
transform 1 0 17696 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_152
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_155
timestamp 1698431365
transform 1 0 18704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_163
timestamp 1698431365
transform 1 0 19600 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_181
timestamp 1698431365
transform 1 0 21616 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_232
timestamp 1698431365
transform 1 0 27328 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_240
timestamp 1698431365
transform 1 0 28224 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_244
timestamp 1698431365
transform 1 0 28672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_250
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_258
timestamp 1698431365
transform 1 0 30240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_262
timestamp 1698431365
transform 1 0 30688 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_270
timestamp 1698431365
transform 1 0 31584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_303
timestamp 1698431365
transform 1 0 35280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_338
timestamp 1698431365
transform 1 0 39200 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_416
timestamp 1698431365
transform 1 0 47936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_433
timestamp 1698431365
transform 1 0 49840 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_464
timestamp 1698431365
transform 1 0 53312 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_480
timestamp 1698431365
transform 1 0 55104 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_488
timestamp 1698431365
transform 1 0 56000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_31
timestamp 1698431365
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_52
timestamp 1698431365
transform 1 0 7168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_61
timestamp 1698431365
transform 1 0 8176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_63
timestamp 1698431365
transform 1 0 8400 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_70
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_72
timestamp 1698431365
transform 1 0 9408 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_102
timestamp 1698431365
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698431365
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_133
timestamp 1698431365
transform 1 0 16240 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_141
timestamp 1698431365
transform 1 0 17136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_203
timestamp 1698431365
transform 1 0 24080 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_262
timestamp 1698431365
transform 1 0 30688 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_278
timestamp 1698431365
transform 1 0 32480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_308
timestamp 1698431365
transform 1 0 35840 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_323
timestamp 1698431365
transform 1 0 37520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_335
timestamp 1698431365
transform 1 0 38864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_339
timestamp 1698431365
transform 1 0 39312 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_405
timestamp 1698431365
transform 1 0 46704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_443
timestamp 1698431365
transform 1 0 50960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_447
timestamp 1698431365
transform 1 0 51408 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_489
timestamp 1698431365
transform 1 0 56112 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_505
timestamp 1698431365
transform 1 0 57904 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_14
timestamp 1698431365
transform 1 0 2912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_59
timestamp 1698431365
transform 1 0 7952 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_67
timestamp 1698431365
transform 1 0 8848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_76
timestamp 1698431365
transform 1 0 9856 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_92
timestamp 1698431365
transform 1 0 11648 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_170
timestamp 1698431365
transform 1 0 20384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_245
timestamp 1698431365
transform 1 0 28784 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_252
timestamp 1698431365
transform 1 0 29568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_268
timestamp 1698431365
transform 1 0 31360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_303
timestamp 1698431365
transform 1 0 35280 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_329
timestamp 1698431365
transform 1 0 38192 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_406
timestamp 1698431365
transform 1 0 46816 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_458
timestamp 1698431365
transform 1 0 52640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_462
timestamp 1698431365
transform 1 0 53088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_478
timestamp 1698431365
transform 1 0 54880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698431365
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_18
timestamp 1698431365
transform 1 0 3360 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_22
timestamp 1698431365
transform 1 0 3808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_24
timestamp 1698431365
transform 1 0 4032 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_46
timestamp 1698431365
transform 1 0 6496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_50
timestamp 1698431365
transform 1 0 6944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_52
timestamp 1698431365
transform 1 0 7168 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_68
timestamp 1698431365
transform 1 0 8960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_72
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_80
timestamp 1698431365
transform 1 0 10304 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_84
timestamp 1698431365
transform 1 0 10752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_109
timestamp 1698431365
transform 1 0 13552 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_112
timestamp 1698431365
transform 1 0 13888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_131
timestamp 1698431365
transform 1 0 16016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_135
timestamp 1698431365
transform 1 0 16464 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_222
timestamp 1698431365
transform 1 0 26208 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698431365
transform 1 0 28000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_276
timestamp 1698431365
transform 1 0 32256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_280
timestamp 1698431365
transform 1 0 32704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_282
timestamp 1698431365
transform 1 0 32928 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_297
timestamp 1698431365
transform 1 0 34608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_310
timestamp 1698431365
transform 1 0 36064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_375
timestamp 1698431365
transform 1 0 43344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_407
timestamp 1698431365
transform 1 0 46928 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_432
timestamp 1698431365
transform 1 0 49728 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_453
timestamp 1698431365
transform 1 0 52080 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_461
timestamp 1698431365
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_465
timestamp 1698431365
transform 1 0 53424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_469
timestamp 1698431365
transform 1 0 53872 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_501
timestamp 1698431365
transform 1 0 57456 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_18
timestamp 1698431365
transform 1 0 3360 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_22
timestamp 1698431365
transform 1 0 3808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_53
timestamp 1698431365
transform 1 0 7280 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_55
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_62
timestamp 1698431365
transform 1 0 8288 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_102
timestamp 1698431365
transform 1 0 12768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_106
timestamp 1698431365
transform 1 0 13216 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_122
timestamp 1698431365
transform 1 0 15008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_124
timestamp 1698431365
transform 1 0 15232 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_131
timestamp 1698431365
transform 1 0 16016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_196
timestamp 1698431365
transform 1 0 23296 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_228
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_236
timestamp 1698431365
transform 1 0 27776 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_252
timestamp 1698431365
transform 1 0 29568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_268
timestamp 1698431365
transform 1 0 31360 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_272
timestamp 1698431365
transform 1 0 31808 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_300
timestamp 1698431365
transform 1 0 34944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_302
timestamp 1698431365
transform 1 0 35168 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_309
timestamp 1698431365
transform 1 0 35952 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_362
timestamp 1698431365
transform 1 0 41888 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_419
timestamp 1698431365
transform 1 0 48272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_449
timestamp 1698431365
transform 1 0 51632 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_479
timestamp 1698431365
transform 1 0 54992 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_487
timestamp 1698431365
transform 1 0 55888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_489
timestamp 1698431365
transform 1 0 56112 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_43
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_47
timestamp 1698431365
transform 1 0 6608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_99
timestamp 1698431365
transform 1 0 12432 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_103
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_122
timestamp 1698431365
transform 1 0 15008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_124
timestamp 1698431365
transform 1 0 15232 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_162
timestamp 1698431365
transform 1 0 19488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_166
timestamp 1698431365
transform 1 0 19936 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_179
timestamp 1698431365
transform 1 0 21392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_186
timestamp 1698431365
transform 1 0 22176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_192
timestamp 1698431365
transform 1 0 22848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_212
timestamp 1698431365
transform 1 0 25088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_249
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_332
timestamp 1698431365
transform 1 0 38528 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_336
timestamp 1698431365
transform 1 0 38976 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_359
timestamp 1698431365
transform 1 0 41552 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_378
timestamp 1698431365
transform 1 0 43680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_380
timestamp 1698431365
transform 1 0 43904 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_405
timestamp 1698431365
transform 1 0 46704 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_452
timestamp 1698431365
transform 1 0 51968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_466
timestamp 1698431365
transform 1 0 53536 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_472
timestamp 1698431365
transform 1 0 54208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_476
timestamp 1698431365
transform 1 0 54656 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_508
timestamp 1698431365
transform 1 0 58240 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_34
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_42
timestamp 1698431365
transform 1 0 6048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_44
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698431365
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_76
timestamp 1698431365
transform 1 0 9856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_80
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_87
timestamp 1698431365
transform 1 0 11088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_95
timestamp 1698431365
transform 1 0 11984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_126
timestamp 1698431365
transform 1 0 15456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_130
timestamp 1698431365
transform 1 0 15904 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_150
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_196
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_228
timestamp 1698431365
transform 1 0 26880 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_236
timestamp 1698431365
transform 1 0 27776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_240
timestamp 1698431365
transform 1 0 28224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_242
timestamp 1698431365
transform 1 0 28448 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_255
timestamp 1698431365
transform 1 0 29904 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_263
timestamp 1698431365
transform 1 0 30800 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_267
timestamp 1698431365
transform 1 0 31248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_269
timestamp 1698431365
transform 1 0 31472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_272
timestamp 1698431365
transform 1 0 31808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_293
timestamp 1698431365
transform 1 0 34160 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_299
timestamp 1698431365
transform 1 0 34832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_301
timestamp 1698431365
transform 1 0 35056 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_315
timestamp 1698431365
transform 1 0 36624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_364
timestamp 1698431365
transform 1 0 42112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_370
timestamp 1698431365
transform 1 0 42784 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_374
timestamp 1698431365
transform 1 0 43232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_378
timestamp 1698431365
transform 1 0 43680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_380
timestamp 1698431365
transform 1 0 43904 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_426
timestamp 1698431365
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_480
timestamp 1698431365
transform 1 0 55104 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_488
timestamp 1698431365
transform 1 0 56000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_508
timestamp 1698431365
transform 1 0 58240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_43
timestamp 1698431365
transform 1 0 6160 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_58
timestamp 1698431365
transform 1 0 7840 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_74
timestamp 1698431365
transform 1 0 9632 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_97
timestamp 1698431365
transform 1 0 12208 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_113
timestamp 1698431365
transform 1 0 14000 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_129
timestamp 1698431365
transform 1 0 15792 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_225
timestamp 1698431365
transform 1 0 26544 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_263
timestamp 1698431365
transform 1 0 30800 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_267
timestamp 1698431365
transform 1 0 31248 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_301
timestamp 1698431365
transform 1 0 35056 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_323
timestamp 1698431365
transform 1 0 37520 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_327
timestamp 1698431365
transform 1 0 37968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_343
timestamp 1698431365
transform 1 0 39760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_347
timestamp 1698431365
transform 1 0 40208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_351
timestamp 1698431365
transform 1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_353
timestamp 1698431365
transform 1 0 40880 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_461
timestamp 1698431365
transform 1 0 52976 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_472
timestamp 1698431365
transform 1 0 54208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_505
timestamp 1698431365
transform 1 0 57904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_101
timestamp 1698431365
transform 1 0 12656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_105
timestamp 1698431365
transform 1 0 13104 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_154
timestamp 1698431365
transform 1 0 18592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_191
timestamp 1698431365
transform 1 0 22736 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_214
timestamp 1698431365
transform 1 0 25312 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_417
timestamp 1698431365
transform 1 0 48048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_419
timestamp 1698431365
transform 1 0 48272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_428
timestamp 1698431365
transform 1 0 49280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_432
timestamp 1698431365
transform 1 0 49728 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_445
timestamp 1698431365
transform 1 0 51184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_474
timestamp 1698431365
transform 1 0 54432 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_498
timestamp 1698431365
transform 1 0 57120 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_506
timestamp 1698431365
transform 1 0 58016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_68
timestamp 1698431365
transform 1 0 8960 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_76
timestamp 1698431365
transform 1 0 9856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_95
timestamp 1698431365
transform 1 0 11984 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_136
timestamp 1698431365
transform 1 0 16576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_140
timestamp 1698431365
transform 1 0 17024 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_148
timestamp 1698431365
transform 1 0 17920 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_154
timestamp 1698431365
transform 1 0 18592 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_164
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_183
timestamp 1698431365
transform 1 0 21840 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_253
timestamp 1698431365
transform 1 0 29680 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_257
timestamp 1698431365
transform 1 0 30128 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_265
timestamp 1698431365
transform 1 0 31024 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_269
timestamp 1698431365
transform 1 0 31472 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_271
timestamp 1698431365
transform 1 0 31696 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_307
timestamp 1698431365
transform 1 0 35728 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_326
timestamp 1698431365
transform 1 0 37856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_330
timestamp 1698431365
transform 1 0 38304 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_360
timestamp 1698431365
transform 1 0 41664 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_372
timestamp 1698431365
transform 1 0 43008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_374
timestamp 1698431365
transform 1 0 43232 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_377
timestamp 1698431365
transform 1 0 43568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_416
timestamp 1698431365
transform 1 0 47936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_495
timestamp 1698431365
transform 1 0 56784 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_503
timestamp 1698431365
transform 1 0 57680 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_507
timestamp 1698431365
transform 1 0 58128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_34
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_36
timestamp 1698431365
transform 1 0 5376 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_80
timestamp 1698431365
transform 1 0 10304 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_92
timestamp 1698431365
transform 1 0 11648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_94
timestamp 1698431365
transform 1 0 11872 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_124
timestamp 1698431365
transform 1 0 15232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_128
timestamp 1698431365
transform 1 0 15680 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_163
timestamp 1698431365
transform 1 0 19600 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_179
timestamp 1698431365
transform 1 0 21392 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_193
timestamp 1698431365
transform 1 0 22960 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_197
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_224
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_232
timestamp 1698431365
transform 1 0 27328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_234
timestamp 1698431365
transform 1 0 27552 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_266
timestamp 1698431365
transform 1 0 31136 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_270
timestamp 1698431365
transform 1 0 31584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_305
timestamp 1698431365
transform 1 0 35504 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_337
timestamp 1698431365
transform 1 0 39088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_341
timestamp 1698431365
transform 1 0 39536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_356
timestamp 1698431365
transform 1 0 41216 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_372
timestamp 1698431365
transform 1 0 43008 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_380
timestamp 1698431365
transform 1 0 43904 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_386
timestamp 1698431365
transform 1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_414
timestamp 1698431365
transform 1 0 47712 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_418
timestamp 1698431365
transform 1 0 48160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_484
timestamp 1698431365
transform 1 0 55552 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_488
timestamp 1698431365
transform 1 0 56000 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_53
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_61
timestamp 1698431365
transform 1 0 8176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_65
timestamp 1698431365
transform 1 0 8624 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_95
timestamp 1698431365
transform 1 0 11984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_99
timestamp 1698431365
transform 1 0 12432 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_123
timestamp 1698431365
transform 1 0 15120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_125
timestamp 1698431365
transform 1 0 15344 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_194
timestamp 1698431365
transform 1 0 23072 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_210
timestamp 1698431365
transform 1 0 24864 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_214
timestamp 1698431365
transform 1 0 25312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_216
timestamp 1698431365
transform 1 0 25536 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_233
timestamp 1698431365
transform 1 0 27440 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_237
timestamp 1698431365
transform 1 0 27888 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_239
timestamp 1698431365
transform 1 0 28112 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_310
timestamp 1698431365
transform 1 0 36064 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_345
timestamp 1698431365
transform 1 0 39984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_357
timestamp 1698431365
transform 1 0 41328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_359
timestamp 1698431365
transform 1 0 41552 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_376
timestamp 1698431365
transform 1 0 43456 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_395
timestamp 1698431365
transform 1 0 45584 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_426
timestamp 1698431365
transform 1 0 49056 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_436
timestamp 1698431365
transform 1 0 50176 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_444
timestamp 1698431365
transform 1 0 51072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_446
timestamp 1698431365
transform 1 0 51296 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_463
timestamp 1698431365
transform 1 0 53200 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_472
timestamp 1698431365
transform 1 0 54208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_503
timestamp 1698431365
transform 1 0 57680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_507
timestamp 1698431365
transform 1 0 58128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_116
timestamp 1698431365
transform 1 0 14336 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_120
timestamp 1698431365
transform 1 0 14784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_160
timestamp 1698431365
transform 1 0 19264 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_241
timestamp 1698431365
transform 1 0 28336 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_245
timestamp 1698431365
transform 1 0 28784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_251
timestamp 1698431365
transform 1 0 29456 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_264
timestamp 1698431365
transform 1 0 30912 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_340
timestamp 1698431365
transform 1 0 39424 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_348
timestamp 1698431365
transform 1 0 40320 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_378
timestamp 1698431365
transform 1 0 43680 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_397
timestamp 1698431365
transform 1 0 45808 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_401
timestamp 1698431365
transform 1 0 46256 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_418
timestamp 1698431365
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_424
timestamp 1698431365
transform 1 0 48832 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_441
timestamp 1698431365
transform 1 0 50736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_445
timestamp 1698431365
transform 1 0 51184 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_449
timestamp 1698431365
transform 1 0 51632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_476
timestamp 1698431365
transform 1 0 54656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_480
timestamp 1698431365
transform 1 0 55104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_484
timestamp 1698431365
transform 1 0 55552 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_488
timestamp 1698431365
transform 1 0 56000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_109
timestamp 1698431365
transform 1 0 13552 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_122
timestamp 1698431365
transform 1 0 15008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_124
timestamp 1698431365
transform 1 0 15232 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_150
timestamp 1698431365
transform 1 0 18144 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_160
timestamp 1698431365
transform 1 0 19264 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_164
timestamp 1698431365
transform 1 0 19712 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_229
timestamp 1698431365
transform 1 0 26992 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_233
timestamp 1698431365
transform 1 0 27440 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_261
timestamp 1698431365
transform 1 0 30576 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_294
timestamp 1698431365
transform 1 0 34272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_298
timestamp 1698431365
transform 1 0 34720 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_306
timestamp 1698431365
transform 1 0 35616 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_310
timestamp 1698431365
transform 1 0 36064 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_331
timestamp 1698431365
transform 1 0 38416 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_335
timestamp 1698431365
transform 1 0 38864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_337
timestamp 1698431365
transform 1 0 39088 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_350
timestamp 1698431365
transform 1 0 40544 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_354
timestamp 1698431365
transform 1 0 40992 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_391
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_399
timestamp 1698431365
transform 1 0 46032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_403
timestamp 1698431365
transform 1 0 46480 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_428
timestamp 1698431365
transform 1 0 49280 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_438
timestamp 1698431365
transform 1 0 50400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_454
timestamp 1698431365
transform 1 0 52192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_465
timestamp 1698431365
transform 1 0 53424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_467
timestamp 1698431365
transform 1 0 53648 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_96
timestamp 1698431365
transform 1 0 12096 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_126
timestamp 1698431365
transform 1 0 15456 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_132
timestamp 1698431365
transform 1 0 16128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_146
timestamp 1698431365
transform 1 0 17696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_148
timestamp 1698431365
transform 1 0 17920 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_178
timestamp 1698431365
transform 1 0 21280 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_208
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_228
timestamp 1698431365
transform 1 0 26880 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_259
timestamp 1698431365
transform 1 0 30352 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_269
timestamp 1698431365
transform 1 0 31472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_271
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_286
timestamp 1698431365
transform 1 0 33376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_296
timestamp 1698431365
transform 1 0 34496 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_304
timestamp 1698431365
transform 1 0 35392 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_307
timestamp 1698431365
transform 1 0 35728 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_315
timestamp 1698431365
transform 1 0 36624 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_324
timestamp 1698431365
transform 1 0 37632 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_340
timestamp 1698431365
transform 1 0 39424 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_348
timestamp 1698431365
transform 1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_356
timestamp 1698431365
transform 1 0 41216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_366
timestamp 1698431365
transform 1 0 42336 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_370
timestamp 1698431365
transform 1 0 42784 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_373
timestamp 1698431365
transform 1 0 43120 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_385
timestamp 1698431365
transform 1 0 44464 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_393
timestamp 1698431365
transform 1 0 45360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_395
timestamp 1698431365
transform 1 0 45584 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_413
timestamp 1698431365
transform 1 0 47600 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_417
timestamp 1698431365
transform 1 0 48048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698431365
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_439
timestamp 1698431365
transform 1 0 50512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_443
timestamp 1698431365
transform 1 0 50960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_447
timestamp 1698431365
transform 1 0 51408 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_489
timestamp 1698431365
transform 1 0 56112 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_496
timestamp 1698431365
transform 1 0 56896 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_504
timestamp 1698431365
transform 1 0 57792 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_508
timestamp 1698431365
transform 1 0 58240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_136
timestamp 1698431365
transform 1 0 16576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_140
timestamp 1698431365
transform 1 0 17024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_144
timestamp 1698431365
transform 1 0 17472 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_159
timestamp 1698431365
transform 1 0 19152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_163
timestamp 1698431365
transform 1 0 19600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_173
timestamp 1698431365
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_181
timestamp 1698431365
transform 1 0 21616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_191
timestamp 1698431365
transform 1 0 22736 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_195
timestamp 1698431365
transform 1 0 23184 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_229
timestamp 1698431365
transform 1 0 26992 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_253
timestamp 1698431365
transform 1 0 29680 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_257
timestamp 1698431365
transform 1 0 30128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_261
timestamp 1698431365
transform 1 0 30576 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_277
timestamp 1698431365
transform 1 0 32368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_279
timestamp 1698431365
transform 1 0 32592 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_290
timestamp 1698431365
transform 1 0 33824 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_294
timestamp 1698431365
transform 1 0 34272 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_296
timestamp 1698431365
transform 1 0 34496 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_306
timestamp 1698431365
transform 1 0 35616 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_346
timestamp 1698431365
transform 1 0 40096 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_350
timestamp 1698431365
transform 1 0 40544 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_358
timestamp 1698431365
transform 1 0 41440 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_362
timestamp 1698431365
transform 1 0 41888 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_372
timestamp 1698431365
transform 1 0 43008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_376
timestamp 1698431365
transform 1 0 43456 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_383
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_395
timestamp 1698431365
transform 1 0 45584 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_399
timestamp 1698431365
transform 1 0 46032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_412
timestamp 1698431365
transform 1 0 47488 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_428
timestamp 1698431365
transform 1 0 49280 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_432
timestamp 1698431365
transform 1 0 49728 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_459
timestamp 1698431365
transform 1 0 52752 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_104
timestamp 1698431365
transform 1 0 12992 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_112
timestamp 1698431365
transform 1 0 13888 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_122
timestamp 1698431365
transform 1 0 15008 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_128
timestamp 1698431365
transform 1 0 15680 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_176
timestamp 1698431365
transform 1 0 21056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_180
timestamp 1698431365
transform 1 0 21504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_184
timestamp 1698431365
transform 1 0 21952 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_188
timestamp 1698431365
transform 1 0 22400 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_190
timestamp 1698431365
transform 1 0 22624 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_193
timestamp 1698431365
transform 1 0 22960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_197
timestamp 1698431365
transform 1 0 23408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_201
timestamp 1698431365
transform 1 0 23856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_203
timestamp 1698431365
transform 1 0 24080 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_216
timestamp 1698431365
transform 1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_343
timestamp 1698431365
transform 1 0 39760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_347
timestamp 1698431365
transform 1 0 40208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_370
timestamp 1698431365
transform 1 0 42784 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_400
timestamp 1698431365
transform 1 0 46144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_404
timestamp 1698431365
transform 1 0 46592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_408
timestamp 1698431365
transform 1 0 47040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_438
timestamp 1698431365
transform 1 0 50400 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_482
timestamp 1698431365
transform 1 0 55328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_506
timestamp 1698431365
transform 1 0 58016 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_113
timestamp 1698431365
transform 1 0 14000 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_152
timestamp 1698431365
transform 1 0 18368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_181
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_191
timestamp 1698431365
transform 1 0 22736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_222
timestamp 1698431365
transform 1 0 26208 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_231
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_239
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_253
timestamp 1698431365
transform 1 0 29680 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_263
timestamp 1698431365
transform 1 0 30800 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_279
timestamp 1698431365
transform 1 0 32592 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_283
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_306
timestamp 1698431365
transform 1 0 35616 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_310
timestamp 1698431365
transform 1 0 36064 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_334
timestamp 1698431365
transform 1 0 38752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_336
timestamp 1698431365
transform 1 0 38976 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_366
timestamp 1698431365
transform 1 0 42336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_370
timestamp 1698431365
transform 1 0 42784 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_374
timestamp 1698431365
transform 1 0 43232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_398
timestamp 1698431365
transform 1 0 45920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_467
timestamp 1698431365
transform 1 0 53648 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_506
timestamp 1698431365
transform 1 0 58016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_508
timestamp 1698431365
transform 1 0 58240 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_88
timestamp 1698431365
transform 1 0 11200 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_92
timestamp 1698431365
transform 1 0 11648 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_124
timestamp 1698431365
transform 1 0 15232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_189
timestamp 1698431365
transform 1 0 22512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_218
timestamp 1698431365
transform 1 0 25760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_220
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_223
timestamp 1698431365
transform 1 0 26320 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_231
timestamp 1698431365
transform 1 0 27216 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_235
timestamp 1698431365
transform 1 0 27664 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_256
timestamp 1698431365
transform 1 0 30016 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_265
timestamp 1698431365
transform 1 0 31024 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_273
timestamp 1698431365
transform 1 0 31920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_294
timestamp 1698431365
transform 1 0 34272 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_310
timestamp 1698431365
transform 1 0 36064 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_345
timestamp 1698431365
transform 1 0 39984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_368
timestamp 1698431365
transform 1 0 42560 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_372
timestamp 1698431365
transform 1 0 43008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_374
timestamp 1698431365
transform 1 0 43232 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_377
timestamp 1698431365
transform 1 0 43568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_381
timestamp 1698431365
transform 1 0 44016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_401
timestamp 1698431365
transform 1 0 46256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_405
timestamp 1698431365
transform 1 0 46704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_428
timestamp 1698431365
transform 1 0 49280 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_472
timestamp 1698431365
transform 1 0 54208 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_165
timestamp 1698431365
transform 1 0 19824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_192
timestamp 1698431365
transform 1 0 22848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_204
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_218
timestamp 1698431365
transform 1 0 25760 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_226
timestamp 1698431365
transform 1 0 26656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_230
timestamp 1698431365
transform 1 0 27104 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_237
timestamp 1698431365
transform 1 0 27888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_249
timestamp 1698431365
transform 1 0 29232 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_258
timestamp 1698431365
transform 1 0 30240 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_280
timestamp 1698431365
transform 1 0 32704 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_294
timestamp 1698431365
transform 1 0 34272 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_302
timestamp 1698431365
transform 1 0 35168 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_306
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_338
timestamp 1698431365
transform 1 0 39200 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_369
timestamp 1698431365
transform 1 0 42672 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_373
timestamp 1698431365
transform 1 0 43120 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_404
timestamp 1698431365
transform 1 0 46592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_408
timestamp 1698431365
transform 1 0 47040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_410
timestamp 1698431365
transform 1 0 47264 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_419
timestamp 1698431365
transform 1 0 48272 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_444
timestamp 1698431365
transform 1 0 51072 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_448
timestamp 1698431365
transform 1 0 51520 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_451
timestamp 1698431365
transform 1 0 51856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_502
timestamp 1698431365
transform 1 0 57568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_506
timestamp 1698431365
transform 1 0 58016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_508
timestamp 1698431365
transform 1 0 58240 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_10
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_14
timestamp 1698431365
transform 1 0 2912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_16
timestamp 1698431365
transform 1 0 3136 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_39
timestamp 1698431365
transform 1 0 5712 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_43
timestamp 1698431365
transform 1 0 6160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_50
timestamp 1698431365
transform 1 0 6944 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_80
timestamp 1698431365
transform 1 0 10304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_84
timestamp 1698431365
transform 1 0 10752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_190
timestamp 1698431365
transform 1 0 22624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_192
timestamp 1698431365
transform 1 0 22848 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_203
timestamp 1698431365
transform 1 0 24080 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_224
timestamp 1698431365
transform 1 0 26432 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_228
timestamp 1698431365
transform 1 0 26880 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_258
timestamp 1698431365
transform 1 0 30240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_262
timestamp 1698431365
transform 1 0 30688 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_271
timestamp 1698431365
transform 1 0 31696 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_399
timestamp 1698431365
transform 1 0 46032 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_415
timestamp 1698431365
transform 1 0 47824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_417
timestamp 1698431365
transform 1 0 48048 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_430
timestamp 1698431365
transform 1 0 49504 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_434
timestamp 1698431365
transform 1 0 49952 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_484
timestamp 1698431365
transform 1 0 55552 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_496
timestamp 1698431365
transform 1 0 56896 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_500
timestamp 1698431365
transform 1 0 57344 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_31
timestamp 1698431365
transform 1 0 4816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_68
timestamp 1698431365
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_72
timestamp 1698431365
transform 1 0 9408 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_102
timestamp 1698431365
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_187
timestamp 1698431365
transform 1 0 22288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_191
timestamp 1698431365
transform 1 0 22736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_195
timestamp 1698431365
transform 1 0 23184 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_199
timestamp 1698431365
transform 1 0 23632 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_201
timestamp 1698431365
transform 1 0 23856 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_216
timestamp 1698431365
transform 1 0 25536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_218
timestamp 1698431365
transform 1 0 25760 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_227
timestamp 1698431365
transform 1 0 26768 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_234
timestamp 1698431365
transform 1 0 27552 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_236
timestamp 1698431365
transform 1 0 27776 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_249
timestamp 1698431365
transform 1 0 29232 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_256
timestamp 1698431365
transform 1 0 30016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_260
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_267
timestamp 1698431365
transform 1 0 31248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_269
timestamp 1698431365
transform 1 0 31472 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_299
timestamp 1698431365
transform 1 0 34832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_303
timestamp 1698431365
transform 1 0 35280 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_336
timestamp 1698431365
transform 1 0 38976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_344
timestamp 1698431365
transform 1 0 39872 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_360
timestamp 1698431365
transform 1 0 41664 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_364
timestamp 1698431365
transform 1 0 42112 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_372
timestamp 1698431365
transform 1 0 43008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_374
timestamp 1698431365
transform 1 0 43232 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_381
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_400
timestamp 1698431365
transform 1 0 46144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_404
timestamp 1698431365
transform 1 0 46592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_406
timestamp 1698431365
transform 1 0 46816 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_440
timestamp 1698431365
transform 1 0 50624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_442
timestamp 1698431365
transform 1 0 50848 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_453
timestamp 1698431365
transform 1 0 52080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_466
timestamp 1698431365
transform 1 0 53536 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_482
timestamp 1698431365
transform 1 0 55328 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_498
timestamp 1698431365
transform 1 0 57120 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_506
timestamp 1698431365
transform 1 0 58016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_508
timestamp 1698431365
transform 1 0 58240 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_31
timestamp 1698431365
transform 1 0 4816 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_58
timestamp 1698431365
transform 1 0 7840 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_88
timestamp 1698431365
transform 1 0 11200 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_96
timestamp 1698431365
transform 1 0 12096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_100
timestamp 1698431365
transform 1 0 12544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_104
timestamp 1698431365
transform 1 0 12992 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_108
timestamp 1698431365
transform 1 0 13440 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_112
timestamp 1698431365
transform 1 0 13888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_129
timestamp 1698431365
transform 1 0 15792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_137
timestamp 1698431365
transform 1 0 16688 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_139
timestamp 1698431365
transform 1 0 16912 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_180
timestamp 1698431365
transform 1 0 21504 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_218
timestamp 1698431365
transform 1 0 25760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_222
timestamp 1698431365
transform 1 0 26208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_226
timestamp 1698431365
transform 1 0 26656 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_236
timestamp 1698431365
transform 1 0 27776 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_244
timestamp 1698431365
transform 1 0 28672 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_250
timestamp 1698431365
transform 1 0 29344 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_258
timestamp 1698431365
transform 1 0 30240 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_270
timestamp 1698431365
transform 1 0 31584 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_278
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_286
timestamp 1698431365
transform 1 0 33376 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_295
timestamp 1698431365
transform 1 0 34384 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_311
timestamp 1698431365
transform 1 0 36176 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_319
timestamp 1698431365
transform 1 0 37072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_335
timestamp 1698431365
transform 1 0 38864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_339
timestamp 1698431365
transform 1 0 39312 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_347
timestamp 1698431365
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_349
timestamp 1698431365
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_354
timestamp 1698431365
transform 1 0 40992 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_377
timestamp 1698431365
transform 1 0 43568 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_396
timestamp 1698431365
transform 1 0 45696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_400
timestamp 1698431365
transform 1 0 46144 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_419
timestamp 1698431365
transform 1 0 48272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_434
timestamp 1698431365
transform 1 0 49952 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_436
timestamp 1698431365
transform 1 0 50176 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_466
timestamp 1698431365
transform 1 0 53536 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_482
timestamp 1698431365
transform 1 0 55328 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_508
timestamp 1698431365
transform 1 0 58240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_18
timestamp 1698431365
transform 1 0 3360 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_22
timestamp 1698431365
transform 1 0 3808 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_50
timestamp 1698431365
transform 1 0 6944 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_68
timestamp 1698431365
transform 1 0 8960 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_84
timestamp 1698431365
transform 1 0 10752 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_88
timestamp 1698431365
transform 1 0 11200 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_166
timestamp 1698431365
transform 1 0 19936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_170
timestamp 1698431365
transform 1 0 20384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_172
timestamp 1698431365
transform 1 0 20608 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_185
timestamp 1698431365
transform 1 0 22064 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_192
timestamp 1698431365
transform 1 0 22848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_204
timestamp 1698431365
transform 1 0 24192 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_208
timestamp 1698431365
transform 1 0 24640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_222
timestamp 1698431365
transform 1 0 26208 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_260
timestamp 1698431365
transform 1 0 30464 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_268
timestamp 1698431365
transform 1 0 31360 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_272
timestamp 1698431365
transform 1 0 31808 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_288
timestamp 1698431365
transform 1 0 33600 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_304
timestamp 1698431365
transform 1 0 35392 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_312
timestamp 1698431365
transform 1 0 36288 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_346
timestamp 1698431365
transform 1 0 40096 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_350
timestamp 1698431365
transform 1 0 40544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_381
timestamp 1698431365
transform 1 0 44016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_404
timestamp 1698431365
transform 1 0 46592 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_438
timestamp 1698431365
transform 1 0 50400 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_452
timestamp 1698431365
transform 1 0 51968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_454
timestamp 1698431365
transform 1 0 52192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_489
timestamp 1698431365
transform 1 0 56112 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_505
timestamp 1698431365
transform 1 0 57904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_18
timestamp 1698431365
transform 1 0 3360 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_34
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_36
timestamp 1698431365
transform 1 0 5376 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_107
timestamp 1698431365
transform 1 0 13328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_109
timestamp 1698431365
transform 1 0 13552 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_146
timestamp 1698431365
transform 1 0 17696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_160
timestamp 1698431365
transform 1 0 19264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_172
timestamp 1698431365
transform 1 0 20608 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_176
timestamp 1698431365
transform 1 0 21056 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_190
timestamp 1698431365
transform 1 0 22624 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_225
timestamp 1698431365
transform 1 0 26544 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_235
timestamp 1698431365
transform 1 0 27664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_257
timestamp 1698431365
transform 1 0 30128 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_261
timestamp 1698431365
transform 1 0 30576 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_298
timestamp 1698431365
transform 1 0 34720 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_334
timestamp 1698431365
transform 1 0 38752 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_338
timestamp 1698431365
transform 1 0 39200 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_348
timestamp 1698431365
transform 1 0 40320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_381
timestamp 1698431365
transform 1 0 44016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_403
timestamp 1698431365
transform 1 0 46480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_407
timestamp 1698431365
transform 1 0 46928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_411
timestamp 1698431365
transform 1 0 47376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_415
timestamp 1698431365
transform 1 0 47824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_417
timestamp 1698431365
transform 1 0 48048 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_455
timestamp 1698431365
transform 1 0 52304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_459
timestamp 1698431365
transform 1 0 52752 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_475
timestamp 1698431365
transform 1 0 54544 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_483
timestamp 1698431365
transform 1 0 55440 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_487
timestamp 1698431365
transform 1 0 55888 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_489
timestamp 1698431365
transform 1 0 56112 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_31
timestamp 1698431365
transform 1 0 4816 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_39
timestamp 1698431365
transform 1 0 5712 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_54
timestamp 1698431365
transform 1 0 7392 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_56
timestamp 1698431365
transform 1 0 7616 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_88
timestamp 1698431365
transform 1 0 11200 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_92
timestamp 1698431365
transform 1 0 11648 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_102
timestamp 1698431365
transform 1 0 12768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_118
timestamp 1698431365
transform 1 0 14560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_120
timestamp 1698431365
transform 1 0 14784 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_129
timestamp 1698431365
transform 1 0 15792 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_134
timestamp 1698431365
transform 1 0 16352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_138
timestamp 1698431365
transform 1 0 16800 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_199
timestamp 1698431365
transform 1 0 23632 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_207
timestamp 1698431365
transform 1 0 24528 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_211
timestamp 1698431365
transform 1 0 24976 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_240
timestamp 1698431365
transform 1 0 28224 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_244
timestamp 1698431365
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_263
timestamp 1698431365
transform 1 0 30800 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_271
timestamp 1698431365
transform 1 0 31696 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_309
timestamp 1698431365
transform 1 0 35952 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_313
timestamp 1698431365
transform 1 0 36400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_329
timestamp 1698431365
transform 1 0 38192 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_333
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_345
timestamp 1698431365
transform 1 0 39984 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_353
timestamp 1698431365
transform 1 0 40880 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_416
timestamp 1698431365
transform 1 0 47936 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_420
timestamp 1698431365
transform 1 0 48384 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_426
timestamp 1698431365
transform 1 0 49056 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_430
timestamp 1698431365
transform 1 0 49504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_452
timestamp 1698431365
transform 1 0 51968 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_454
timestamp 1698431365
transform 1 0 52192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_489
timestamp 1698431365
transform 1 0 56112 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_505
timestamp 1698431365
transform 1 0 57904 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_10
timestamp 1698431365
transform 1 0 2464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_76
timestamp 1698431365
transform 1 0 9856 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_84
timestamp 1698431365
transform 1 0 10752 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_92
timestamp 1698431365
transform 1 0 11648 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_96
timestamp 1698431365
transform 1 0 12096 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_99
timestamp 1698431365
transform 1 0 12432 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_107
timestamp 1698431365
transform 1 0 13328 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_111
timestamp 1698431365
transform 1 0 13776 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_123
timestamp 1698431365
transform 1 0 15120 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_125
timestamp 1698431365
transform 1 0 15344 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_128
timestamp 1698431365
transform 1 0 15680 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_170
timestamp 1698431365
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_186
timestamp 1698431365
transform 1 0 22176 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_200
timestamp 1698431365
transform 1 0 23744 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_208
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_227
timestamp 1698431365
transform 1 0 26768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_261
timestamp 1698431365
transform 1 0 30576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_288
timestamp 1698431365
transform 1 0 33600 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_296
timestamp 1698431365
transform 1 0 34496 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_298
timestamp 1698431365
transform 1 0 34720 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_313
timestamp 1698431365
transform 1 0 36400 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_317
timestamp 1698431365
transform 1 0 36848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_321
timestamp 1698431365
transform 1 0 37296 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_329
timestamp 1698431365
transform 1 0 38192 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_360
timestamp 1698431365
transform 1 0 41664 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_362
timestamp 1698431365
transform 1 0 41888 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_406
timestamp 1698431365
transform 1 0 46816 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_414
timestamp 1698431365
transform 1 0 47712 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_418
timestamp 1698431365
transform 1 0 48160 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_474
timestamp 1698431365
transform 1 0 54432 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_10
timestamp 1698431365
transform 1 0 2464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_14
timestamp 1698431365
transform 1 0 2912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_16
timestamp 1698431365
transform 1 0 3136 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_25
timestamp 1698431365
transform 1 0 4144 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_31
timestamp 1698431365
transform 1 0 4816 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_86
timestamp 1698431365
transform 1 0 10976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_88
timestamp 1698431365
transform 1 0 11200 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_97
timestamp 1698431365
transform 1 0 12208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_122
timestamp 1698431365
transform 1 0 15008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_124
timestamp 1698431365
transform 1 0 15232 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_136
timestamp 1698431365
transform 1 0 16576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_151
timestamp 1698431365
transform 1 0 18256 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_158
timestamp 1698431365
transform 1 0 19040 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_169
timestamp 1698431365
transform 1 0 20272 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_173
timestamp 1698431365
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_181
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_183
timestamp 1698431365
transform 1 0 21840 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_201
timestamp 1698431365
transform 1 0 23856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_205
timestamp 1698431365
transform 1 0 24304 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_232
timestamp 1698431365
transform 1 0 27328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_236
timestamp 1698431365
transform 1 0 27776 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_253
timestamp 1698431365
transform 1 0 29680 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_266
timestamp 1698431365
transform 1 0 31136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_270
timestamp 1698431365
transform 1 0 31584 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_278
timestamp 1698431365
transform 1 0 32480 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_281
timestamp 1698431365
transform 1 0 32816 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_289
timestamp 1698431365
transform 1 0 33712 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_313
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_346
timestamp 1698431365
transform 1 0 40096 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_371
timestamp 1698431365
transform 1 0 42896 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_379
timestamp 1698431365
transform 1 0 43792 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_383
timestamp 1698431365
transform 1 0 44240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_391
timestamp 1698431365
transform 1 0 45136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_395
timestamp 1698431365
transform 1 0 45584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_399
timestamp 1698431365
transform 1 0 46032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_454
timestamp 1698431365
transform 1 0 52192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_489
timestamp 1698431365
transform 1 0 56112 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_505
timestamp 1698431365
transform 1 0 57904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_74
timestamp 1698431365
transform 1 0 9632 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_82
timestamp 1698431365
transform 1 0 10528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_117
timestamp 1698431365
transform 1 0 14448 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_127
timestamp 1698431365
transform 1 0 15568 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_164
timestamp 1698431365
transform 1 0 19712 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_192
timestamp 1698431365
transform 1 0 22848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_248
timestamp 1698431365
transform 1 0 29120 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_273
timestamp 1698431365
transform 1 0 31920 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_277
timestamp 1698431365
transform 1 0 32368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_288
timestamp 1698431365
transform 1 0 33600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_292
timestamp 1698431365
transform 1 0 34048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_329
timestamp 1698431365
transform 1 0 38192 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_346
timestamp 1698431365
transform 1 0 40096 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_368
timestamp 1698431365
transform 1 0 42560 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_376
timestamp 1698431365
transform 1 0 43456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_380
timestamp 1698431365
transform 1 0 43904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_382
timestamp 1698431365
transform 1 0 44128 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_403
timestamp 1698431365
transform 1 0 46480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_407
timestamp 1698431365
transform 1 0 46928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_411
timestamp 1698431365
transform 1 0 47376 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_419
timestamp 1698431365
transform 1 0 48272 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_440
timestamp 1698431365
transform 1 0 50624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_442
timestamp 1698431365
transform 1 0 50848 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_451
timestamp 1698431365
transform 1 0 51856 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_483
timestamp 1698431365
transform 1 0 55440 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_487
timestamp 1698431365
transform 1 0 55888 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_489
timestamp 1698431365
transform 1 0 56112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_6
timestamp 1698431365
transform 1 0 2016 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_30
timestamp 1698431365
transform 1 0 4704 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_66
timestamp 1698431365
transform 1 0 8736 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_68
timestamp 1698431365
transform 1 0 8960 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_71
timestamp 1698431365
transform 1 0 9296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_75
timestamp 1698431365
transform 1 0 9744 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_85
timestamp 1698431365
transform 1 0 10864 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_91
timestamp 1698431365
transform 1 0 11536 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_95
timestamp 1698431365
transform 1 0 11984 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_102
timestamp 1698431365
transform 1 0 12768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_124
timestamp 1698431365
transform 1 0 15232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_128
timestamp 1698431365
transform 1 0 15680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_132
timestamp 1698431365
transform 1 0 16128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_170
timestamp 1698431365
transform 1 0 20384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_179
timestamp 1698431365
transform 1 0 21392 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_212
timestamp 1698431365
transform 1 0 25088 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_214
timestamp 1698431365
transform 1 0 25312 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_238
timestamp 1698431365
transform 1 0 28000 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_275
timestamp 1698431365
transform 1 0 32144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_283
timestamp 1698431365
transform 1 0 33040 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_285
timestamp 1698431365
transform 1 0 33264 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_300
timestamp 1698431365
transform 1 0 34944 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_308
timestamp 1698431365
transform 1 0 35840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1698431365
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_327
timestamp 1698431365
transform 1 0 37968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_329
timestamp 1698431365
transform 1 0 38192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_336
timestamp 1698431365
transform 1 0 38976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_350
timestamp 1698431365
transform 1 0 40544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_416
timestamp 1698431365
transform 1 0 47936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_420
timestamp 1698431365
transform 1 0 48384 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_436
timestamp 1698431365
transform 1 0 50176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_440
timestamp 1698431365
transform 1 0 50624 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_443
timestamp 1698431365
transform 1 0 50960 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_451
timestamp 1698431365
transform 1 0 51856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_489
timestamp 1698431365
transform 1 0 56112 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_505
timestamp 1698431365
transform 1 0 57904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_6
timestamp 1698431365
transform 1 0 2016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_8
timestamp 1698431365
transform 1 0 2240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_54
timestamp 1698431365
transform 1 0 7392 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_62
timestamp 1698431365
transform 1 0 8288 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_91
timestamp 1698431365
transform 1 0 11536 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_100
timestamp 1698431365
transform 1 0 12544 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_108
timestamp 1698431365
transform 1 0 13440 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_112
timestamp 1698431365
transform 1 0 13888 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_114
timestamp 1698431365
transform 1 0 14112 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_120
timestamp 1698431365
transform 1 0 14784 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_122
timestamp 1698431365
transform 1 0 15008 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_128
timestamp 1698431365
transform 1 0 15680 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_132
timestamp 1698431365
transform 1 0 16128 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_158
timestamp 1698431365
transform 1 0 19040 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_160
timestamp 1698431365
transform 1 0 19264 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_204
timestamp 1698431365
transform 1 0 24192 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_208
timestamp 1698431365
transform 1 0 24640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_214
timestamp 1698431365
transform 1 0 25312 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_240
timestamp 1698431365
transform 1 0 28224 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_325
timestamp 1698431365
transform 1 0 37744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_327
timestamp 1698431365
transform 1 0 37968 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_334
timestamp 1698431365
transform 1 0 38752 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_338
timestamp 1698431365
transform 1 0 39200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_370
timestamp 1698431365
transform 1 0 42784 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_378
timestamp 1698431365
transform 1 0 43680 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_382
timestamp 1698431365
transform 1 0 44128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_384
timestamp 1698431365
transform 1 0 44352 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_387
timestamp 1698431365
transform 1 0 44688 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698431365
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_457
timestamp 1698431365
transform 1 0 52528 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_489
timestamp 1698431365
transform 1 0 56112 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_31
timestamp 1698431365
transform 1 0 4816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_53
timestamp 1698431365
transform 1 0 7280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_55
timestamp 1698431365
transform 1 0 7504 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_87
timestamp 1698431365
transform 1 0 11088 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_91
timestamp 1698431365
transform 1 0 11536 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_95
timestamp 1698431365
transform 1 0 11984 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_111
timestamp 1698431365
transform 1 0 13776 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_124
timestamp 1698431365
transform 1 0 15232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_126
timestamp 1698431365
transform 1 0 15456 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_132
timestamp 1698431365
transform 1 0 16128 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_136
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_138
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_158
timestamp 1698431365
transform 1 0 19040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_174
timestamp 1698431365
transform 1 0 20832 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_187
timestamp 1698431365
transform 1 0 22288 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_208
timestamp 1698431365
transform 1 0 24640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_210
timestamp 1698431365
transform 1 0 24864 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_223
timestamp 1698431365
transform 1 0 26320 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_225
timestamp 1698431365
transform 1 0 26544 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_242
timestamp 1698431365
transform 1 0 28448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_244
timestamp 1698431365
transform 1 0 28672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_254
timestamp 1698431365
transform 1 0 29792 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_276
timestamp 1698431365
transform 1 0 32256 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_285
timestamp 1698431365
transform 1 0 33264 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_301
timestamp 1698431365
transform 1 0 35056 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_309
timestamp 1698431365
transform 1 0 35952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_313
timestamp 1698431365
transform 1 0 36400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_333
timestamp 1698431365
transform 1 0 38640 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_358
timestamp 1698431365
transform 1 0 41440 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_374
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_378
timestamp 1698431365
transform 1 0 43680 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_380
timestamp 1698431365
transform 1 0 43904 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_383
timestamp 1698431365
transform 1 0 44240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_391
timestamp 1698431365
transform 1 0 45136 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_393
timestamp 1698431365
transform 1 0 45360 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_400
timestamp 1698431365
transform 1 0 46144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_431
timestamp 1698431365
transform 1 0 49616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_435
timestamp 1698431365
transform 1 0 50064 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_443
timestamp 1698431365
transform 1 0 50960 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698431365
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_489
timestamp 1698431365
transform 1 0 56112 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_505
timestamp 1698431365
transform 1 0 57904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_6
timestamp 1698431365
transform 1 0 2016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_8
timestamp 1698431365
transform 1 0 2240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_26
timestamp 1698431365
transform 1 0 4256 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_42
timestamp 1698431365
transform 1 0 6048 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_49
timestamp 1698431365
transform 1 0 6832 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_59
timestamp 1698431365
transform 1 0 7952 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_67
timestamp 1698431365
transform 1 0 8848 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_69
timestamp 1698431365
transform 1 0 9072 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_80
timestamp 1698431365
transform 1 0 10304 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_137
timestamp 1698431365
transform 1 0 16688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_139
timestamp 1698431365
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_150
timestamp 1698431365
transform 1 0 18144 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_175
timestamp 1698431365
transform 1 0 20944 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_224
timestamp 1698431365
transform 1 0 26432 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_235
timestamp 1698431365
transform 1 0 27664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_288
timestamp 1698431365
transform 1 0 33600 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_290
timestamp 1698431365
transform 1 0 33824 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_299
timestamp 1698431365
transform 1 0 34832 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_305
timestamp 1698431365
transform 1 0 35504 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_309
timestamp 1698431365
transform 1 0 35952 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_340
timestamp 1698431365
transform 1 0 39424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_381
timestamp 1698431365
transform 1 0 44016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_383
timestamp 1698431365
transform 1 0 44240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_392
timestamp 1698431365
transform 1 0 45248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_394
timestamp 1698431365
transform 1 0 45472 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_413
timestamp 1698431365
transform 1 0 47600 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_417
timestamp 1698431365
transform 1 0 48048 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_419
timestamp 1698431365
transform 1 0 48272 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_442
timestamp 1698431365
transform 1 0 50848 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_446
timestamp 1698431365
transform 1 0 51296 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_478
timestamp 1698431365
transform 1 0 54880 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698431365
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698431365
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_31
timestamp 1698431365
transform 1 0 4816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_39
timestamp 1698431365
transform 1 0 5712 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_58
timestamp 1698431365
transform 1 0 7840 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_88
timestamp 1698431365
transform 1 0 11200 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_96
timestamp 1698431365
transform 1 0 12096 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_100
timestamp 1698431365
transform 1 0 12544 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_149
timestamp 1698431365
transform 1 0 18032 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_151
timestamp 1698431365
transform 1 0 18256 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_166
timestamp 1698431365
transform 1 0 19936 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_168
timestamp 1698431365
transform 1 0 20160 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_182
timestamp 1698431365
transform 1 0 21728 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_186
timestamp 1698431365
transform 1 0 22176 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_196
timestamp 1698431365
transform 1 0 23296 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_200
timestamp 1698431365
transform 1 0 23744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_202
timestamp 1698431365
transform 1 0 23968 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_205
timestamp 1698431365
transform 1 0 24304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_209
timestamp 1698431365
transform 1 0 24752 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_219
timestamp 1698431365
transform 1 0 25872 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_227
timestamp 1698431365
transform 1 0 26768 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_262
timestamp 1698431365
transform 1 0 30688 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_270
timestamp 1698431365
transform 1 0 31584 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_321
timestamp 1698431365
transform 1 0 37296 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_353
timestamp 1698431365
transform 1 0 40880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_355
timestamp 1698431365
transform 1 0 41104 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_395
timestamp 1698431365
transform 1 0 45584 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_428
timestamp 1698431365
transform 1 0 49280 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_450
timestamp 1698431365
transform 1 0 51744 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1698431365
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_489
timestamp 1698431365
transform 1 0 56112 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_505
timestamp 1698431365
transform 1 0 57904 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_10
timestamp 1698431365
transform 1 0 2464 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_17
timestamp 1698431365
transform 1 0 3248 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_21
timestamp 1698431365
transform 1 0 3696 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_63
timestamp 1698431365
transform 1 0 8400 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_82
timestamp 1698431365
transform 1 0 10528 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_86
timestamp 1698431365
transform 1 0 10976 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_156
timestamp 1698431365
transform 1 0 18816 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_168
timestamp 1698431365
transform 1 0 20160 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_173
timestamp 1698431365
transform 1 0 20720 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_177
timestamp 1698431365
transform 1 0 21168 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_181
timestamp 1698431365
transform 1 0 21616 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_189
timestamp 1698431365
transform 1 0 22512 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_203
timestamp 1698431365
transform 1 0 24080 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_228
timestamp 1698431365
transform 1 0 26880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_230
timestamp 1698431365
transform 1 0 27104 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_240
timestamp 1698431365
transform 1 0 28224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_309
timestamp 1698431365
transform 1 0 35952 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_313
timestamp 1698431365
transform 1 0 36400 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_345
timestamp 1698431365
transform 1 0 39984 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_349
timestamp 1698431365
transform 1 0 40432 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_368
timestamp 1698431365
transform 1 0 42560 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_389
timestamp 1698431365
transform 1 0 44912 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_416
timestamp 1698431365
transform 1 0 47936 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_430
timestamp 1698431365
transform 1 0 49504 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_466
timestamp 1698431365
transform 1 0 53536 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_482
timestamp 1698431365
transform 1 0 55328 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_18
timestamp 1698431365
transform 1 0 3360 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_20
timestamp 1698431365
transform 1 0 3584 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_61
timestamp 1698431365
transform 1 0 8176 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_65
timestamp 1698431365
transform 1 0 8624 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_81
timestamp 1698431365
transform 1 0 10416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_91
timestamp 1698431365
transform 1 0 11536 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_99
timestamp 1698431365
transform 1 0 12432 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_103
timestamp 1698431365
transform 1 0 12880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_174
timestamp 1698431365
transform 1 0 20832 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_185
timestamp 1698431365
transform 1 0 22064 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_189
timestamp 1698431365
transform 1 0 22512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_205
timestamp 1698431365
transform 1 0 24304 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_219
timestamp 1698431365
transform 1 0 25872 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_223
timestamp 1698431365
transform 1 0 26320 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_225
timestamp 1698431365
transform 1 0 26544 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_228
timestamp 1698431365
transform 1 0 26880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_255
timestamp 1698431365
transform 1 0 29904 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_257
timestamp 1698431365
transform 1 0 30128 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_264
timestamp 1698431365
transform 1 0 30912 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_302
timestamp 1698431365
transform 1 0 35168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_306
timestamp 1698431365
transform 1 0 35616 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_313
timestamp 1698431365
transform 1 0 36400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_332
timestamp 1698431365
transform 1 0 38528 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_334
timestamp 1698431365
transform 1 0 38752 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_353
timestamp 1698431365
transform 1 0 40880 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_367
timestamp 1698431365
transform 1 0 42448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_369
timestamp 1698431365
transform 1 0 42672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_416
timestamp 1698431365
transform 1 0 47936 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_420
timestamp 1698431365
transform 1 0 48384 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_430
timestamp 1698431365
transform 1 0 49504 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_445
timestamp 1698431365
transform 1 0 51184 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_449
timestamp 1698431365
transform 1 0 51632 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_453
timestamp 1698431365
transform 1 0 52080 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_489
timestamp 1698431365
transform 1 0 56112 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_505
timestamp 1698431365
transform 1 0 57904 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_31
timestamp 1698431365
transform 1 0 4816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_64
timestamp 1698431365
transform 1 0 8512 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_68
timestamp 1698431365
transform 1 0 8960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_90
timestamp 1698431365
transform 1 0 11424 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_94
timestamp 1698431365
transform 1 0 11872 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_149
timestamp 1698431365
transform 1 0 18032 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_159
timestamp 1698431365
transform 1 0 19152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_180
timestamp 1698431365
transform 1 0 21504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_198
timestamp 1698431365
transform 1 0 23520 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_207
timestamp 1698431365
transform 1 0 24528 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_209
timestamp 1698431365
transform 1 0 24752 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_228
timestamp 1698431365
transform 1 0 26880 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_232
timestamp 1698431365
transform 1 0 27328 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_262
timestamp 1698431365
transform 1 0 30688 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_277
timestamp 1698431365
transform 1 0 32368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_279
timestamp 1698431365
transform 1 0 32592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_347
timestamp 1698431365
transform 1 0 40208 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698431365
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_358
timestamp 1698431365
transform 1 0 41440 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_366
timestamp 1698431365
transform 1 0 42336 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_382
timestamp 1698431365
transform 1 0 44128 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_386
timestamp 1698431365
transform 1 0 44576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_390
timestamp 1698431365
transform 1 0 45024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_418
timestamp 1698431365
transform 1 0 48160 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_440
timestamp 1698431365
transform 1 0 50624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_444
timestamp 1698431365
transform 1 0 51072 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_476
timestamp 1698431365
transform 1 0 54656 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_484
timestamp 1698431365
transform 1 0 55552 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_488
timestamp 1698431365
transform 1 0 56000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1698431365
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_31
timestamp 1698431365
transform 1 0 4816 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_57
timestamp 1698431365
transform 1 0 7728 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_95
timestamp 1698431365
transform 1 0 11984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_139
timestamp 1698431365
transform 1 0 16912 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_162
timestamp 1698431365
transform 1 0 19488 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_172
timestamp 1698431365
transform 1 0 20608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_174
timestamp 1698431365
transform 1 0 20832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_185
timestamp 1698431365
transform 1 0 22064 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_187
timestamp 1698431365
transform 1 0 22288 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_194
timestamp 1698431365
transform 1 0 23072 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_213
timestamp 1698431365
transform 1 0 25200 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_217
timestamp 1698431365
transform 1 0 25648 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_233
timestamp 1698431365
transform 1 0 27440 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_243
timestamp 1698431365
transform 1 0 28560 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_255
timestamp 1698431365
transform 1 0 29904 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_259
timestamp 1698431365
transform 1 0 30352 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_261
timestamp 1698431365
transform 1 0 30576 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_264
timestamp 1698431365
transform 1 0 30912 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_313
timestamp 1698431365
transform 1 0 36400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_380
timestamp 1698431365
transform 1 0 43904 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698431365
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_424
timestamp 1698431365
transform 1 0 48832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_426
timestamp 1698431365
transform 1 0 49056 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_448
timestamp 1698431365
transform 1 0 51520 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_452
timestamp 1698431365
transform 1 0 51968 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_454
timestamp 1698431365
transform 1 0 52192 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_486
timestamp 1698431365
transform 1 0 55776 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_502
timestamp 1698431365
transform 1 0 57568 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_506
timestamp 1698431365
transform 1 0 58016 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_508
timestamp 1698431365
transform 1 0 58240 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_18
timestamp 1698431365
transform 1 0 3360 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_26
timestamp 1698431365
transform 1 0 4256 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_64
timestamp 1698431365
transform 1 0 8512 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_68
timestamp 1698431365
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_76
timestamp 1698431365
transform 1 0 9856 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_99
timestamp 1698431365
transform 1 0 12432 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_119
timestamp 1698431365
transform 1 0 14672 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_139
timestamp 1698431365
transform 1 0 16912 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_160
timestamp 1698431365
transform 1 0 19264 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_164
timestamp 1698431365
transform 1 0 19712 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_173
timestamp 1698431365
transform 1 0 20720 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_181
timestamp 1698431365
transform 1 0 21616 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_183
timestamp 1698431365
transform 1 0 21840 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_202
timestamp 1698431365
transform 1 0 23968 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_270
timestamp 1698431365
transform 1 0 31584 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_274
timestamp 1698431365
transform 1 0 32032 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_278
timestamp 1698431365
transform 1 0 32480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_322
timestamp 1698431365
transform 1 0 37408 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_347
timestamp 1698431365
transform 1 0 40208 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1698431365
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_354
timestamp 1698431365
transform 1 0 40992 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_381
timestamp 1698431365
transform 1 0 44016 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_389
timestamp 1698431365
transform 1 0 44912 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_393
timestamp 1698431365
transform 1 0 45360 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_410
timestamp 1698431365
transform 1 0 47264 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_416
timestamp 1698431365
transform 1 0 47936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_477
timestamp 1698431365
transform 1 0 54768 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_485
timestamp 1698431365
transform 1 0 55664 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_489
timestamp 1698431365
transform 1 0 56112 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698431365
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_18
timestamp 1698431365
transform 1 0 3360 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_22
timestamp 1698431365
transform 1 0 3808 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_32
timestamp 1698431365
transform 1 0 4928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_57
timestamp 1698431365
transform 1 0 7728 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_61
timestamp 1698431365
transform 1 0 8176 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_91
timestamp 1698431365
transform 1 0 11536 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_153
timestamp 1698431365
transform 1 0 18480 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_157
timestamp 1698431365
transform 1 0 18928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_161
timestamp 1698431365
transform 1 0 19376 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_163
timestamp 1698431365
transform 1 0 19600 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_166
timestamp 1698431365
transform 1 0 19936 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_239
timestamp 1698431365
transform 1 0 28112 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_243
timestamp 1698431365
transform 1 0 28560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_255
timestamp 1698431365
transform 1 0 29904 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_257
timestamp 1698431365
transform 1 0 30128 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_287
timestamp 1698431365
transform 1 0 33488 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_291
timestamp 1698431365
transform 1 0 33936 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_299
timestamp 1698431365
transform 1 0 34832 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_303
timestamp 1698431365
transform 1 0 35280 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_313
timestamp 1698431365
transform 1 0 36400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_348
timestamp 1698431365
transform 1 0 40320 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_374
timestamp 1698431365
transform 1 0 43232 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_382
timestamp 1698431365
transform 1 0 44128 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_384
timestamp 1698431365
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_395
timestamp 1698431365
transform 1 0 45584 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_417
timestamp 1698431365
transform 1 0 48048 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_425
timestamp 1698431365
transform 1 0 48944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_453
timestamp 1698431365
transform 1 0 52080 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_489
timestamp 1698431365
transform 1 0 56112 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_505
timestamp 1698431365
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_34
timestamp 1698431365
transform 1 0 5152 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_50
timestamp 1698431365
transform 1 0 6944 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_58
timestamp 1698431365
transform 1 0 7840 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_62
timestamp 1698431365
transform 1 0 8288 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_76
timestamp 1698431365
transform 1 0 9856 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_78
timestamp 1698431365
transform 1 0 10080 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_87
timestamp 1698431365
transform 1 0 11088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_105
timestamp 1698431365
transform 1 0 13104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_115
timestamp 1698431365
transform 1 0 14224 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_131
timestamp 1698431365
transform 1 0 16016 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_133
timestamp 1698431365
transform 1 0 16240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_138
timestamp 1698431365
transform 1 0 16800 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_144
timestamp 1698431365
transform 1 0 17472 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_195
timestamp 1698431365
transform 1 0 23184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_218
timestamp 1698431365
transform 1 0 25760 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_222
timestamp 1698431365
transform 1 0 26208 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_230
timestamp 1698431365
transform 1 0 27104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_261
timestamp 1698431365
transform 1 0 30576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_265
timestamp 1698431365
transform 1 0 31024 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_269
timestamp 1698431365
transform 1 0 31472 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_271
timestamp 1698431365
transform 1 0 31696 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_278
timestamp 1698431365
transform 1 0 32480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_290
timestamp 1698431365
transform 1 0 33824 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_318
timestamp 1698431365
transform 1 0 36960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_349
timestamp 1698431365
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_357
timestamp 1698431365
transform 1 0 41328 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_359
timestamp 1698431365
transform 1 0 41552 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_383
timestamp 1698431365
transform 1 0 44240 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_387
timestamp 1698431365
transform 1 0 44688 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_417
timestamp 1698431365
transform 1 0 48048 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_419
timestamp 1698431365
transform 1 0 48272 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_441
timestamp 1698431365
transform 1 0 50736 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_473
timestamp 1698431365
transform 1 0 54320 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_489
timestamp 1698431365
transform 1 0 56112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698431365
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_31
timestamp 1698431365
transform 1 0 4816 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_69
timestamp 1698431365
transform 1 0 9072 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_104
timestamp 1698431365
transform 1 0 12992 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_113
timestamp 1698431365
transform 1 0 14000 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_129
timestamp 1698431365
transform 1 0 15792 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_137
timestamp 1698431365
transform 1 0 16688 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_209
timestamp 1698431365
transform 1 0 24752 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_213
timestamp 1698431365
transform 1 0 25200 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_255
timestamp 1698431365
transform 1 0 29904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_259
timestamp 1698431365
transform 1 0 30352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_261
timestamp 1698431365
transform 1 0 30576 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_291
timestamp 1698431365
transform 1 0 33936 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_295
timestamp 1698431365
transform 1 0 34384 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_299
timestamp 1698431365
transform 1 0 34832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_312
timestamp 1698431365
transform 1 0 36288 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_314
timestamp 1698431365
transform 1 0 36512 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_321
timestamp 1698431365
transform 1 0 37296 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_323
timestamp 1698431365
transform 1 0 37520 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_349
timestamp 1698431365
transform 1 0 40432 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_357
timestamp 1698431365
transform 1 0 41328 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_361
timestamp 1698431365
transform 1 0 41776 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_363
timestamp 1698431365
transform 1 0 42000 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_372
timestamp 1698431365
transform 1 0 43008 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_380
timestamp 1698431365
transform 1 0 43904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_384
timestamp 1698431365
transform 1 0 44352 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_395
timestamp 1698431365
transform 1 0 45584 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_403
timestamp 1698431365
transform 1 0 46480 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_419
timestamp 1698431365
transform 1 0 48272 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_450
timestamp 1698431365
transform 1 0 51744 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_454
timestamp 1698431365
transform 1 0 52192 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_489
timestamp 1698431365
transform 1 0 56112 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_505
timestamp 1698431365
transform 1 0 57904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_6
timestamp 1698431365
transform 1 0 2016 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_34
timestamp 1698431365
transform 1 0 5152 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_38
timestamp 1698431365
transform 1 0 5600 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_58
timestamp 1698431365
transform 1 0 7840 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_88
timestamp 1698431365
transform 1 0 11200 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_129
timestamp 1698431365
transform 1 0 15792 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_131
timestamp 1698431365
transform 1 0 16016 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_144
timestamp 1698431365
transform 1 0 17472 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_166
timestamp 1698431365
transform 1 0 19936 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_170
timestamp 1698431365
transform 1 0 20384 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_209
timestamp 1698431365
transform 1 0 24752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_216
timestamp 1698431365
transform 1 0 25536 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_220
timestamp 1698431365
transform 1 0 25984 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_225
timestamp 1698431365
transform 1 0 26544 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_251
timestamp 1698431365
transform 1 0 29456 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_261
timestamp 1698431365
transform 1 0 30576 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_269
timestamp 1698431365
transform 1 0 31472 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_273
timestamp 1698431365
transform 1 0 31920 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_276
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_286
timestamp 1698431365
transform 1 0 33376 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_294
timestamp 1698431365
transform 1 0 34272 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_327
timestamp 1698431365
transform 1 0 37968 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_335
timestamp 1698431365
transform 1 0 38864 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_340
timestamp 1698431365
transform 1 0 39424 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_345
timestamp 1698431365
transform 1 0 39984 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_349
timestamp 1698431365
transform 1 0 40432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_356
timestamp 1698431365
transform 1 0 41216 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_364
timestamp 1698431365
transform 1 0 42112 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_397
timestamp 1698431365
transform 1 0 45808 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_413
timestamp 1698431365
transform 1 0 47600 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_417
timestamp 1698431365
transform 1 0 48048 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_419
timestamp 1698431365
transform 1 0 48272 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_31
timestamp 1698431365
transform 1 0 4816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_68
timestamp 1698431365
transform 1 0 8960 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_72
timestamp 1698431365
transform 1 0 9408 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_104
timestamp 1698431365
transform 1 0 12992 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_115
timestamp 1698431365
transform 1 0 14224 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_121
timestamp 1698431365
transform 1 0 14896 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_129
timestamp 1698431365
transform 1 0 15792 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_162
timestamp 1698431365
transform 1 0 19488 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_166
timestamp 1698431365
transform 1 0 19936 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_173
timestamp 1698431365
transform 1 0 20720 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_378
timestamp 1698431365
transform 1 0 43680 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_382
timestamp 1698431365
transform 1 0 44128 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_384
timestamp 1698431365
transform 1 0 44352 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_451
timestamp 1698431365
transform 1 0 51856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_489
timestamp 1698431365
transform 1 0 56112 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_505
timestamp 1698431365
transform 1 0 57904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_18
timestamp 1698431365
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_26
timestamp 1698431365
transform 1 0 4256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_46
timestamp 1698431365
transform 1 0 6496 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_48
timestamp 1698431365
transform 1 0 6720 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_57
timestamp 1698431365
transform 1 0 7728 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_59
timestamp 1698431365
transform 1 0 7952 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_81
timestamp 1698431365
transform 1 0 10416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_93
timestamp 1698431365
transform 1 0 11760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_101
timestamp 1698431365
transform 1 0 12656 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_108
timestamp 1698431365
transform 1 0 13440 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_135
timestamp 1698431365
transform 1 0 16464 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_140
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_147
timestamp 1698431365
transform 1 0 17808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_159
timestamp 1698431365
transform 1 0 19152 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_210
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_224
timestamp 1698431365
transform 1 0 26432 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_244
timestamp 1698431365
transform 1 0 28672 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_253
timestamp 1698431365
transform 1 0 29680 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_267
timestamp 1698431365
transform 1 0 31248 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_284
timestamp 1698431365
transform 1 0 33152 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_298
timestamp 1698431365
transform 1 0 34720 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_318
timestamp 1698431365
transform 1 0 36960 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_332
timestamp 1698431365
transform 1 0 38528 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_396
timestamp 1698431365
transform 1 0 45696 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_405
timestamp 1698431365
transform 1 0 46704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_407
timestamp 1698431365
transform 1 0 46928 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_418
timestamp 1698431365
transform 1 0 48160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_420
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_429
timestamp 1698431365
transform 1 0 49392 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_441
timestamp 1698431365
transform 1 0 50736 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_444
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_453
timestamp 1698431365
transform 1 0 52080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_465
timestamp 1698431365
transform 1 0 53424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_473
timestamp 1698431365
transform 1 0 54320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_475
timestamp 1698431365
transform 1 0 54544 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_490
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_506
timestamp 1698431365
transform 1 0 58016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 19152 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 20384 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 38864 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform 1 0 15792 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 17136 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output7 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23184 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output8 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21056 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output9
timestamp 1698431365
transform 1 0 22624 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output10
timestamp 1698431365
transform -1 0 26432 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output11
timestamp 1698431365
transform -1 0 28000 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output12
timestamp 1698431365
transform 1 0 28336 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output13
timestamp 1698431365
transform 1 0 30128 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output14
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output15
timestamp 1698431365
transform 1 0 33600 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output16
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output17
timestamp 1698431365
transform 1 0 37408 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output18
timestamp 1698431365
transform -1 0 38416 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output19
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output20
timestamp 1698431365
transform -1 0 42784 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_21 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_22
timestamp 1698431365
transform 1 0 21840 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_23
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_24
timestamp 1698431365
transform -1 0 26544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_25
timestamp 1698431365
transform -1 0 28672 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_26
timestamp 1698431365
transform -1 0 29232 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_27
timestamp 1698431365
transform 1 0 29232 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_28
timestamp 1698431365
transform -1 0 31808 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_29
timestamp 1698431365
transform -1 0 33376 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_30
timestamp 1698431365
transform -1 0 35616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_31
timestamp 1698431365
transform -1 0 36624 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_32
timestamp 1698431365
transform -1 0 39424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_33
timestamp 1698431365
transform -1 0 38864 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_34
timestamp 1698431365
transform -1 0 39984 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_35
timestamp 1698431365
transform 1 0 4704 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_36
timestamp 1698431365
transform -1 0 7280 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_37
timestamp 1698431365
transform -1 0 8512 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_38
timestamp 1698431365
transform -1 0 9968 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_39
timestamp 1698431365
transform -1 0 11312 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_40
timestamp 1698431365
transform -1 0 12656 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_41
timestamp 1698431365
transform -1 0 14000 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_42
timestamp 1698431365
transform 1 0 14448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_43
timestamp 1698431365
transform 1 0 14896 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_44
timestamp 1698431365
transform 1 0 15344 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_45
timestamp 1698431365
transform 1 0 18032 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_46
timestamp 1698431365
transform -1 0 20720 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_47
timestamp 1698431365
transform -1 0 41216 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_48
timestamp 1698431365
transform -1 0 43904 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_49
timestamp 1698431365
transform -1 0 43680 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_50
timestamp 1698431365
transform -1 0 45248 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_51
timestamp 1698431365
transform -1 0 46256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_52
timestamp 1698431365
transform -1 0 47712 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_53
timestamp 1698431365
transform -1 0 48944 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_54
timestamp 1698431365
transform -1 0 50288 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_55
timestamp 1698431365
transform -1 0 51632 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_56
timestamp 1698431365
transform -1 0 52976 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_57
timestamp 1698431365
transform -1 0 54320 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  urish_simon_says_58
timestamp 1698431365
transform -1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_59 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_60
timestamp 1698431365
transform -1 0 7728 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_61
timestamp 1698431365
transform -1 0 8960 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_62
timestamp 1698431365
transform -1 0 10416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_63
timestamp 1698431365
transform -1 0 11760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_64
timestamp 1698431365
transform -1 0 13440 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_65
timestamp 1698431365
transform -1 0 14448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_66
timestamp 1698431365
transform -1 0 15792 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_67
timestamp 1698431365
transform 1 0 15904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_68
timestamp 1698431365
transform -1 0 19488 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_69
timestamp 1698431365
transform -1 0 19712 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_70
timestamp 1698431365
transform -1 0 21056 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_71
timestamp 1698431365
transform -1 0 43232 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_72
timestamp 1698431365
transform -1 0 44352 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_73
timestamp 1698431365
transform -1 0 44800 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_74
timestamp 1698431365
transform -1 0 45696 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_75
timestamp 1698431365
transform -1 0 46704 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_76
timestamp 1698431365
transform -1 0 48160 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_77
timestamp 1698431365
transform -1 0 49392 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_78
timestamp 1698431365
transform -1 0 50736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_79
timestamp 1698431365
transform -1 0 52080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_80
timestamp 1698431365
transform -1 0 53424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_81
timestamp 1698431365
transform -1 0 55328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  urish_simon_says_82
timestamp 1698431365
transform -1 0 56224 0 -1 56448
box -86 -86 534 870
<< labels >>
flabel metal2 s 4928 59200 5040 60000 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 18368 59200 18480 60000 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 19712 59200 19824 60000 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 21056 59200 21168 60000 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 22400 59200 22512 60000 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 23744 59200 23856 60000 0 FreeSans 448 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 25088 59200 25200 60000 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 26432 59200 26544 60000 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 27776 59200 27888 60000 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 29120 59200 29232 60000 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 30464 59200 30576 60000 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 6272 59200 6384 60000 0 FreeSans 448 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 31808 59200 31920 60000 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 33152 59200 33264 60000 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 34496 59200 34608 60000 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 35840 59200 35952 60000 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 37184 59200 37296 60000 0 FreeSans 448 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 38528 59200 38640 60000 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 39872 59200 39984 60000 0 FreeSans 448 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 41216 59200 41328 60000 0 FreeSans 448 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 42560 59200 42672 60000 0 FreeSans 448 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 43904 59200 44016 60000 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 7616 59200 7728 60000 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 45248 59200 45360 60000 0 FreeSans 448 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 46592 59200 46704 60000 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 47936 59200 48048 60000 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 49280 59200 49392 60000 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 50624 59200 50736 60000 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 51968 59200 52080 60000 0 FreeSans 448 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 53312 59200 53424 60000 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 54656 59200 54768 60000 0 FreeSans 448 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 8960 59200 9072 60000 0 FreeSans 448 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 10304 59200 10416 60000 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 11648 59200 11760 60000 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 12992 59200 13104 60000 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 14336 59200 14448 60000 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 15680 59200 15792 60000 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 17024 59200 17136 60000 0 FreeSans 448 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 5824 59200 5936 60000 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 19264 59200 19376 60000 0 FreeSans 448 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 20608 59200 20720 60000 0 FreeSans 448 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 21952 59200 22064 60000 0 FreeSans 448 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 23296 59200 23408 60000 0 FreeSans 448 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 24640 59200 24752 60000 0 FreeSans 448 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 25984 59200 26096 60000 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 27328 59200 27440 60000 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 28672 59200 28784 60000 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 30016 59200 30128 60000 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 31360 59200 31472 60000 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 7168 59200 7280 60000 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 32704 59200 32816 60000 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 34048 59200 34160 60000 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 35392 59200 35504 60000 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 36736 59200 36848 60000 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 38080 59200 38192 60000 0 FreeSans 448 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 39424 59200 39536 60000 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 40768 59200 40880 60000 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 42112 59200 42224 60000 0 FreeSans 448 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 43456 59200 43568 60000 0 FreeSans 448 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 44800 59200 44912 60000 0 FreeSans 448 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 8512 59200 8624 60000 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 46144 59200 46256 60000 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 47488 59200 47600 60000 0 FreeSans 448 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 48832 59200 48944 60000 0 FreeSans 448 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 50176 59200 50288 60000 0 FreeSans 448 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 51520 59200 51632 60000 0 FreeSans 448 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 52864 59200 52976 60000 0 FreeSans 448 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 54208 59200 54320 60000 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 55552 59200 55664 60000 0 FreeSans 448 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 9856 59200 9968 60000 0 FreeSans 448 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 11200 59200 11312 60000 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 12544 59200 12656 60000 0 FreeSans 448 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 13888 59200 14000 60000 0 FreeSans 448 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 15232 59200 15344 60000 0 FreeSans 448 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 16576 59200 16688 60000 0 FreeSans 448 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 17920 59200 18032 60000 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 5376 59200 5488 60000 0 FreeSans 448 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 18816 59200 18928 60000 0 FreeSans 448 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 20160 59200 20272 60000 0 FreeSans 448 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 21504 59200 21616 60000 0 FreeSans 448 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 22848 59200 22960 60000 0 FreeSans 448 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 24192 59200 24304 60000 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 25536 59200 25648 60000 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 26880 59200 26992 60000 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 28224 59200 28336 60000 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 29568 59200 29680 60000 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 30912 59200 31024 60000 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 6720 59200 6832 60000 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 32256 59200 32368 60000 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 33600 59200 33712 60000 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 34944 59200 35056 60000 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 36288 59200 36400 60000 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 37632 59200 37744 60000 0 FreeSans 448 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 38976 59200 39088 60000 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 40320 59200 40432 60000 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 41664 59200 41776 60000 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 43008 59200 43120 60000 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 44352 59200 44464 60000 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 8064 59200 8176 60000 0 FreeSans 448 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 45696 59200 45808 60000 0 FreeSans 448 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 47040 59200 47152 60000 0 FreeSans 448 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 48384 59200 48496 60000 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 49728 59200 49840 60000 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 51072 59200 51184 60000 0 FreeSans 448 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 52416 59200 52528 60000 0 FreeSans 448 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 53760 59200 53872 60000 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 55104 59200 55216 60000 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 9408 59200 9520 60000 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 10752 59200 10864 60000 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 12096 59200 12208 60000 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 13440 59200 13552 60000 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 14784 59200 14896 60000 0 FreeSans 448 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 16128 59200 16240 60000 0 FreeSans 448 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 17472 59200 17584 60000 0 FreeSans 448 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 114 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 114 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 115 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 115 nsew ground bidirectional
flabel metal2 s 4032 59200 4144 60000 0 FreeSans 448 90 0 0 wb_clk_i
port 116 nsew signal input
flabel metal2 s 4480 59200 4592 60000 0 FreeSans 448 90 0 0 wb_rst_i
port 117 nsew signal input
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal3 21336 21448 21336 21448 0 _0000_
rlabel metal2 17416 17640 17416 17640 0 _0001_
rlabel metal2 15512 24024 15512 24024 0 _0002_
rlabel metal2 17416 19208 17416 19208 0 _0003_
rlabel metal2 25480 21000 25480 21000 0 _0004_
rlabel metal2 22624 38920 22624 38920 0 _0005_
rlabel metal2 13608 35056 13608 35056 0 _0006_
rlabel metal3 13328 37912 13328 37912 0 _0007_
rlabel metal2 16408 34552 16408 34552 0 _0008_
rlabel metal2 13608 40936 13608 40936 0 _0009_
rlabel metal2 23968 35000 23968 35000 0 _0010_
rlabel metal3 14112 39032 14112 39032 0 _0011_
rlabel metal2 21560 35952 21560 35952 0 _0012_
rlabel metal3 42392 55160 42392 55160 0 _0013_
rlabel metal2 43736 53928 43736 53928 0 _0014_
rlabel metal2 4984 25032 4984 25032 0 _0015_
rlabel metal2 7784 25144 7784 25144 0 _0016_
rlabel metal2 2464 20664 2464 20664 0 _0017_
rlabel metal2 5544 20328 5544 20328 0 _0018_
rlabel metal2 13160 26628 13160 26628 0 _0019_
rlabel metal2 10528 24808 10528 24808 0 _0020_
rlabel metal2 14392 22624 14392 22624 0 _0021_
rlabel metal2 10920 22008 10920 22008 0 _0022_
rlabel metal2 10360 27328 10360 27328 0 _0023_
rlabel metal2 9744 29624 9744 29624 0 _0024_
rlabel metal2 18312 19712 18312 19712 0 _0025_
rlabel metal3 22288 19096 22288 19096 0 _0026_
rlabel metal2 13384 5208 13384 5208 0 _0027_
rlabel metal2 11256 6328 11256 6328 0 _0028_
rlabel metal2 17304 5600 17304 5600 0 _0029_
rlabel metal2 16464 6776 16464 6776 0 _0030_
rlabel metal2 2464 22456 2464 22456 0 _0031_
rlabel metal2 3976 23464 3976 23464 0 _0032_
rlabel metal2 45752 53424 45752 53424 0 _0033_
rlabel metal2 14280 10304 14280 10304 0 _0034_
rlabel metal2 10360 8512 10360 8512 0 _0035_
rlabel metal2 6384 10808 6384 10808 0 _0036_
rlabel metal2 6888 9352 6888 9352 0 _0037_
rlabel metal2 2464 16184 2464 16184 0 _0038_
rlabel metal2 3864 14756 3864 14756 0 _0039_
rlabel metal2 3080 18760 3080 18760 0 _0040_
rlabel metal2 2520 18368 2520 18368 0 _0041_
rlabel metal2 2856 13440 2856 13440 0 _0042_
rlabel metal2 2520 13048 2520 13048 0 _0043_
rlabel metal2 17976 10304 17976 10304 0 _0044_
rlabel metal2 20776 10080 20776 10080 0 _0045_
rlabel metal2 26488 30184 26488 30184 0 _0046_
rlabel metal2 14504 29904 14504 29904 0 _0047_
rlabel metal2 12936 30128 12936 30128 0 _0048_
rlabel metal2 14280 29736 14280 29736 0 _0049_
rlabel metal2 24472 33712 24472 33712 0 _0050_
rlabel metal2 27888 37352 27888 37352 0 _0051_
rlabel metal3 43512 47320 43512 47320 0 _0052_
rlabel metal2 46648 48048 46648 48048 0 _0053_
rlabel metal2 47320 46200 47320 46200 0 _0054_
rlabel metal2 50232 45416 50232 45416 0 _0055_
rlabel metal2 51240 48608 51240 48608 0 _0056_
rlabel metal2 52472 51688 52472 51688 0 _0057_
rlabel metal2 49112 53368 49112 53368 0 _0058_
rlabel metal3 52416 50456 52416 50456 0 _0059_
rlabel metal2 34104 33208 34104 33208 0 _0060_
rlabel metal2 37352 32984 37352 32984 0 _0061_
rlabel metal2 40040 35224 40040 35224 0 _0062_
rlabel metal3 39928 36568 39928 36568 0 _0063_
rlabel metal3 40992 46536 40992 46536 0 _0064_
rlabel metal2 41944 44464 41944 44464 0 _0065_
rlabel metal2 43064 36904 43064 36904 0 _0066_
rlabel metal2 46088 40208 46088 40208 0 _0067_
rlabel metal2 48888 40208 48888 40208 0 _0068_
rlabel metal3 49672 40152 49672 40152 0 _0069_
rlabel metal3 44520 34216 44520 34216 0 _0070_
rlabel metal2 53480 36064 53480 36064 0 _0071_
rlabel metal2 57400 31892 57400 31892 0 _0072_
rlabel metal2 55832 34496 55832 34496 0 _0073_
rlabel metal2 56728 30856 56728 30856 0 _0074_
rlabel metal2 42504 31248 42504 31248 0 _0075_
rlabel metal2 55552 27160 55552 27160 0 _0076_
rlabel metal2 51464 25704 51464 25704 0 _0077_
rlabel metal2 49336 29176 49336 29176 0 _0078_
rlabel metal2 50960 21672 50960 21672 0 _0079_
rlabel metal2 45640 21672 45640 21672 0 _0080_
rlabel metal2 46088 21896 46088 21896 0 _0081_
rlabel metal2 42392 28056 42392 28056 0 _0082_
rlabel metal2 40936 28112 40936 28112 0 _0083_
rlabel metal2 39144 20608 39144 20608 0 _0084_
rlabel metal2 39368 26600 39368 26600 0 _0085_
rlabel metal2 36680 21784 36680 21784 0 _0086_
rlabel metal3 34888 26824 34888 26824 0 _0087_
rlabel metal2 30520 25872 30520 25872 0 _0088_
rlabel metal3 31416 26824 31416 26824 0 _0089_
rlabel metal2 33880 31304 33880 31304 0 _0090_
rlabel metal2 37128 31304 37128 31304 0 _0091_
rlabel metal2 46200 43960 46200 43960 0 _0092_
rlabel metal2 34328 46928 34328 46928 0 _0093_
rlabel metal2 35448 46480 35448 46480 0 _0094_
rlabel metal3 20104 52808 20104 52808 0 _0095_
rlabel metal2 18872 53368 18872 53368 0 _0096_
rlabel metal2 29344 32648 29344 32648 0 _0097_
rlabel metal2 28840 29736 28840 29736 0 _0098_
rlabel metal2 29624 49756 29624 49756 0 _0099_
rlabel metal2 28168 49392 28168 49392 0 _0100_
rlabel metal2 28840 48664 28840 48664 0 _0101_
rlabel metal2 30464 34216 30464 34216 0 _0102_
rlabel metal2 27160 34440 27160 34440 0 _0103_
rlabel metal2 32648 39004 32648 39004 0 _0104_
rlabel metal2 33880 36848 33880 36848 0 _0105_
rlabel metal3 34832 44968 34832 44968 0 _0106_
rlabel metal3 35336 43400 35336 43400 0 _0107_
rlabel metal2 37800 39816 37800 39816 0 _0108_
rlabel metal2 35728 40488 35728 40488 0 _0109_
rlabel metal2 36232 42000 36232 42000 0 _0110_
rlabel metal2 32760 41328 32760 41328 0 _0111_
rlabel metal2 8904 41664 8904 41664 0 _0112_
rlabel metal2 8680 43064 8680 43064 0 _0113_
rlabel metal2 8792 45136 8792 45136 0 _0114_
rlabel metal3 9296 47544 9296 47544 0 _0115_
rlabel metal2 8792 50904 8792 50904 0 _0116_
rlabel metal2 11704 51744 11704 51744 0 _0117_
rlabel metal2 10696 53760 10696 53760 0 _0118_
rlabel metal2 13496 51800 13496 51800 0 _0119_
rlabel metal3 17696 48440 17696 48440 0 _0120_
rlabel metal2 16296 51800 16296 51800 0 _0121_
rlabel metal2 2744 53368 2744 53368 0 _0122_
rlabel metal2 2520 54936 2520 54936 0 _0123_
rlabel metal2 2520 51296 2520 51296 0 _0124_
rlabel metal2 7672 54768 7672 54768 0 _0125_
rlabel metal2 6440 50456 6440 50456 0 _0126_
rlabel metal2 2520 49224 2520 49224 0 _0127_
rlabel metal2 6776 48608 6776 48608 0 _0128_
rlabel metal2 5880 43792 5880 43792 0 _0129_
rlabel metal2 6664 37688 6664 37688 0 _0130_
rlabel metal2 3528 37688 3528 37688 0 _0131_
rlabel metal2 2520 39760 2520 39760 0 _0132_
rlabel metal2 6552 40768 6552 40768 0 _0133_
rlabel metal2 2520 41496 2520 41496 0 _0134_
rlabel metal2 3304 43932 3304 43932 0 _0135_
rlabel metal2 2464 44408 2464 44408 0 _0136_
rlabel metal2 2520 47880 2520 47880 0 _0137_
rlabel metal2 27664 27944 27664 27944 0 _0138_
rlabel metal2 24248 26712 24248 26712 0 _0139_
rlabel metal2 20440 28392 20440 28392 0 _0140_
rlabel metal2 17192 27384 17192 27384 0 _0141_
rlabel metal3 18536 24920 18536 24920 0 _0142_
rlabel metal2 26656 29960 26656 29960 0 _0143_
rlabel metal3 23016 32536 23016 32536 0 _0144_
rlabel metal2 18984 32144 18984 32144 0 _0145_
rlabel metal3 13552 31864 13552 31864 0 _0146_
rlabel metal2 14280 33656 14280 33656 0 _0147_
rlabel metal2 24472 50792 24472 50792 0 _0148_
rlabel metal3 23744 54488 23744 54488 0 _0149_
rlabel metal2 24584 54544 24584 54544 0 _0150_
rlabel metal2 27160 52472 27160 52472 0 _0151_
rlabel metal2 34328 17192 34328 17192 0 _0152_
rlabel metal2 37576 15624 37576 15624 0 _0153_
rlabel metal2 16408 11984 16408 11984 0 _0154_
rlabel metal2 16856 12600 16856 12600 0 _0155_
rlabel metal2 9912 12600 9912 12600 0 _0156_
rlabel metal2 10360 11872 10360 11872 0 _0157_
rlabel metal3 32088 8344 32088 8344 0 _0158_
rlabel metal2 31416 9352 31416 9352 0 _0159_
rlabel metal2 19096 17192 19096 17192 0 _0160_
rlabel metal3 21112 14616 21112 14616 0 _0161_
rlabel metal2 32984 16296 32984 16296 0 _0162_
rlabel metal2 31752 14056 31752 14056 0 _0163_
rlabel metal2 33880 12488 33880 12488 0 _0164_
rlabel metal2 36008 11312 36008 11312 0 _0165_
rlabel metal3 9632 14392 9632 14392 0 _0166_
rlabel metal2 8008 14168 8008 14168 0 _0167_
rlabel metal2 26432 20104 26432 20104 0 _0168_
rlabel metal2 31080 19320 31080 19320 0 _0169_
rlabel metal2 31920 20888 31920 20888 0 _0170_
rlabel metal2 35000 20888 35000 20888 0 _0171_
rlabel metal2 21672 4144 21672 4144 0 _0172_
rlabel metal2 21784 5040 21784 5040 0 _0173_
rlabel metal2 26096 4536 26096 4536 0 _0174_
rlabel metal2 27496 5432 27496 5432 0 _0175_
rlabel metal2 21000 7784 21000 7784 0 _0176_
rlabel metal3 24192 8120 24192 8120 0 _0177_
rlabel metal2 26488 10920 26488 10920 0 _0178_
rlabel metal2 26488 8512 26488 8512 0 _0179_
rlabel metal2 27216 21784 27216 21784 0 _0180_
rlabel metal2 29400 23576 29400 23576 0 _0181_
rlabel metal2 32536 19712 32536 19712 0 _0182_
rlabel metal3 36792 17528 36792 17528 0 _0183_
rlabel metal2 5656 27328 5656 27328 0 _0184_
rlabel metal2 6776 28896 6776 28896 0 _0185_
rlabel metal2 26488 54600 26488 54600 0 _0186_
rlabel metal3 39592 53872 39592 53872 0 _0187_
rlabel metal2 30072 54936 30072 54936 0 _0188_
rlabel metal2 31192 52080 31192 52080 0 _0189_
rlabel metal2 31976 53368 31976 53368 0 _0190_
rlabel metal2 33208 54152 33208 54152 0 _0191_
rlabel metal2 35672 54824 35672 54824 0 _0192_
rlabel metal2 47096 30576 47096 30576 0 _0193_
rlabel metal2 43568 26488 43568 26488 0 _0194_
rlabel metal2 47880 32928 47880 32928 0 _0195_
rlabel metal3 47376 38584 47376 38584 0 _0196_
rlabel metal2 40376 31024 40376 31024 0 _0197_
rlabel metal3 46424 25592 46424 25592 0 _0198_
rlabel metal2 44912 36456 44912 36456 0 _0199_
rlabel metal2 43176 31976 43176 31976 0 _0200_
rlabel metal2 43288 29288 43288 29288 0 _0201_
rlabel metal3 47656 39480 47656 39480 0 _0202_
rlabel metal2 42728 39200 42728 39200 0 _0203_
rlabel metal2 43120 40376 43120 40376 0 _0204_
rlabel metal2 42504 39984 42504 39984 0 _0205_
rlabel metal2 44632 39088 44632 39088 0 _0206_
rlabel metal2 45584 38920 45584 38920 0 _0207_
rlabel metal2 46480 23240 46480 23240 0 _0208_
rlabel metal2 42840 26488 42840 26488 0 _0209_
rlabel metal3 45864 39592 45864 39592 0 _0210_
rlabel metal2 49784 42672 49784 42672 0 _0211_
rlabel metal2 42616 42728 42616 42728 0 _0212_
rlabel metal2 42728 42392 42728 42392 0 _0213_
rlabel metal3 42952 41048 42952 41048 0 _0214_
rlabel metal3 43960 40936 43960 40936 0 _0215_
rlabel metal2 43064 41608 43064 41608 0 _0216_
rlabel metal2 49448 41832 49448 41832 0 _0217_
rlabel metal2 49000 41216 49000 41216 0 _0218_
rlabel metal3 47432 23800 47432 23800 0 _0219_
rlabel metal3 48328 38920 48328 38920 0 _0220_
rlabel metal2 47376 39592 47376 39592 0 _0221_
rlabel metal2 48552 39592 48552 39592 0 _0222_
rlabel metal2 50344 40152 50344 40152 0 _0223_
rlabel metal3 49560 39592 49560 39592 0 _0224_
rlabel metal2 49224 39536 49224 39536 0 _0225_
rlabel metal2 51296 42616 51296 42616 0 _0226_
rlabel metal2 51800 42224 51800 42224 0 _0227_
rlabel metal3 52752 43288 52752 43288 0 _0228_
rlabel metal2 51352 41272 51352 41272 0 _0229_
rlabel metal2 51688 41216 51688 41216 0 _0230_
rlabel metal2 47768 38976 47768 38976 0 _0231_
rlabel metal3 49672 38920 49672 38920 0 _0232_
rlabel metal2 50120 40320 50120 40320 0 _0233_
rlabel metal2 47656 34888 47656 34888 0 _0234_
rlabel metal2 47768 37520 47768 37520 0 _0235_
rlabel metal2 52024 40768 52024 40768 0 _0236_
rlabel metal2 52248 41272 52248 41272 0 _0237_
rlabel metal2 51856 41384 51856 41384 0 _0238_
rlabel metal3 54096 38024 54096 38024 0 _0239_
rlabel metal2 55048 37688 55048 37688 0 _0240_
rlabel metal2 52696 36400 52696 36400 0 _0241_
rlabel metal2 45192 35168 45192 35168 0 _0242_
rlabel metal2 36456 22456 36456 22456 0 _0243_
rlabel metal2 44072 33936 44072 33936 0 _0244_
rlabel metal2 44072 33320 44072 33320 0 _0245_
rlabel metal2 45472 23912 45472 23912 0 _0246_
rlabel metal2 50792 35784 50792 35784 0 _0247_
rlabel metal2 51128 34888 51128 34888 0 _0248_
rlabel metal2 51688 36680 51688 36680 0 _0249_
rlabel metal3 48328 36568 48328 36568 0 _0250_
rlabel metal2 50456 37016 50456 37016 0 _0251_
rlabel metal2 48776 35952 48776 35952 0 _0252_
rlabel metal3 49224 34216 49224 34216 0 _0253_
rlabel metal2 49840 33992 49840 33992 0 _0254_
rlabel metal3 49112 35448 49112 35448 0 _0255_
rlabel metal2 47208 35728 47208 35728 0 _0256_
rlabel metal2 52920 35168 52920 35168 0 _0257_
rlabel metal3 52920 32536 52920 32536 0 _0258_
rlabel metal2 54320 31640 54320 31640 0 _0259_
rlabel metal2 51632 29624 51632 29624 0 _0260_
rlabel metal2 54600 36176 54600 36176 0 _0261_
rlabel metal2 54152 36400 54152 36400 0 _0262_
rlabel metal3 55104 35672 55104 35672 0 _0263_
rlabel metal2 50904 36008 50904 36008 0 _0264_
rlabel metal2 50456 35224 50456 35224 0 _0265_
rlabel metal3 50540 34216 50540 34216 0 _0266_
rlabel metal2 55160 35448 55160 35448 0 _0267_
rlabel metal2 56056 35952 56056 35952 0 _0268_
rlabel metal2 57232 35112 57232 35112 0 _0269_
rlabel metal2 54712 33936 54712 33936 0 _0270_
rlabel metal2 54152 34552 54152 34552 0 _0271_
rlabel metal2 56168 34776 56168 34776 0 _0272_
rlabel metal2 55944 35056 55944 35056 0 _0273_
rlabel metal2 57848 35448 57848 35448 0 _0274_
rlabel metal2 40600 29288 40600 29288 0 _0275_
rlabel metal2 51856 28840 51856 28840 0 _0276_
rlabel metal2 54152 30520 54152 30520 0 _0277_
rlabel metal2 53816 27496 53816 27496 0 _0278_
rlabel metal2 50456 30072 50456 30072 0 _0279_
rlabel metal3 53200 31304 53200 31304 0 _0280_
rlabel metal2 51240 33544 51240 33544 0 _0281_
rlabel metal2 53144 35168 53144 35168 0 _0282_
rlabel metal2 50120 32760 50120 32760 0 _0283_
rlabel metal2 50288 31528 50288 31528 0 _0284_
rlabel metal2 50120 31248 50120 31248 0 _0285_
rlabel metal2 50680 30856 50680 30856 0 _0286_
rlabel metal2 41608 21560 41608 21560 0 _0287_
rlabel metal2 48272 20888 48272 20888 0 _0288_
rlabel metal2 45416 24416 45416 24416 0 _0289_
rlabel metal3 47488 31192 47488 31192 0 _0290_
rlabel metal2 52136 29680 52136 29680 0 _0291_
rlabel metal2 53984 27944 53984 27944 0 _0292_
rlabel metal2 55384 28728 55384 28728 0 _0293_
rlabel metal2 53144 29456 53144 29456 0 _0294_
rlabel metal2 51576 30016 51576 30016 0 _0295_
rlabel metal2 45360 29400 45360 29400 0 _0296_
rlabel metal2 44352 31192 44352 31192 0 _0297_
rlabel metal2 42840 31752 42840 31752 0 _0298_
rlabel metal2 47768 28336 47768 28336 0 _0299_
rlabel metal2 51800 27216 51800 27216 0 _0300_
rlabel metal2 53816 29344 53816 29344 0 _0301_
rlabel metal2 52920 29736 52920 29736 0 _0302_
rlabel metal3 47936 26264 47936 26264 0 _0303_
rlabel metal2 45640 28952 45640 28952 0 _0304_
rlabel metal2 51688 28952 51688 28952 0 _0305_
rlabel metal2 53256 29120 53256 29120 0 _0306_
rlabel metal3 50904 25704 50904 25704 0 _0307_
rlabel metal3 49336 24696 49336 24696 0 _0308_
rlabel metal2 51016 25480 51016 25480 0 _0309_
rlabel metal2 52248 26880 52248 26880 0 _0310_
rlabel metal2 52472 25760 52472 25760 0 _0311_
rlabel metal2 49840 26264 49840 26264 0 _0312_
rlabel metal2 49448 26152 49448 26152 0 _0313_
rlabel metal2 49504 29400 49504 29400 0 _0314_
rlabel metal2 49112 29792 49112 29792 0 _0315_
rlabel metal2 51688 23576 51688 23576 0 _0316_
rlabel metal2 49672 23296 49672 23296 0 _0317_
rlabel metal2 51128 26096 51128 26096 0 _0318_
rlabel metal2 53480 27944 53480 27944 0 _0319_
rlabel metal2 53200 27608 53200 27608 0 _0320_
rlabel metal2 47880 22400 47880 22400 0 _0321_
rlabel metal3 51184 23912 51184 23912 0 _0322_
rlabel metal2 51688 22736 51688 22736 0 _0323_
rlabel metal2 51800 22960 51800 22960 0 _0324_
rlabel metal2 44968 24248 44968 24248 0 _0325_
rlabel metal3 41916 23912 41916 23912 0 _0326_
rlabel metal2 47880 24528 47880 24528 0 _0327_
rlabel metal3 49868 23128 49868 23128 0 _0328_
rlabel metal2 49224 23408 49224 23408 0 _0329_
rlabel metal2 45640 24024 45640 24024 0 _0330_
rlabel metal2 45976 24248 45976 24248 0 _0331_
rlabel metal2 49448 23856 49448 23856 0 _0332_
rlabel metal2 47208 24192 47208 24192 0 _0333_
rlabel metal2 47880 21672 47880 21672 0 _0334_
rlabel metal2 46592 22456 46592 22456 0 _0335_
rlabel metal2 47208 24920 47208 24920 0 _0336_
rlabel metal3 46144 25480 46144 25480 0 _0337_
rlabel metal2 45304 25704 45304 25704 0 _0338_
rlabel metal2 47320 21616 47320 21616 0 _0339_
rlabel metal2 47656 22064 47656 22064 0 _0340_
rlabel metal2 48776 22736 48776 22736 0 _0341_
rlabel metal2 46424 23856 46424 23856 0 _0342_
rlabel metal2 47012 29624 47012 29624 0 _0343_
rlabel metal3 46872 29400 46872 29400 0 _0344_
rlabel metal2 42728 25312 42728 25312 0 _0345_
rlabel metal2 44296 21112 44296 21112 0 _0346_
rlabel metal2 39816 23296 39816 23296 0 _0347_
rlabel metal2 41720 25200 41720 25200 0 _0348_
rlabel metal3 41832 22232 41832 22232 0 _0349_
rlabel metal3 41104 22456 41104 22456 0 _0350_
rlabel metal2 42616 24584 42616 24584 0 _0351_
rlabel metal3 42616 26824 42616 26824 0 _0352_
rlabel metal2 42504 23296 42504 23296 0 _0353_
rlabel metal3 42560 27048 42560 27048 0 _0354_
rlabel metal2 42392 27384 42392 27384 0 _0355_
rlabel metal2 41832 27384 41832 27384 0 _0356_
rlabel metal2 42056 21168 42056 21168 0 _0357_
rlabel metal2 42168 22064 42168 22064 0 _0358_
rlabel metal2 42168 24472 42168 24472 0 _0359_
rlabel metal2 39928 21616 39928 21616 0 _0360_
rlabel metal2 41832 21224 41832 21224 0 _0361_
rlabel metal2 38752 23240 38752 23240 0 _0362_
rlabel metal2 40488 22680 40488 22680 0 _0363_
rlabel metal2 39592 22848 39592 22848 0 _0364_
rlabel metal2 42056 23856 42056 23856 0 _0365_
rlabel metal2 40712 24304 40712 24304 0 _0366_
rlabel metal2 43064 23408 43064 23408 0 _0367_
rlabel metal2 35112 23072 35112 23072 0 _0368_
rlabel metal2 34776 23184 34776 23184 0 _0369_
rlabel metal2 38696 22736 38696 22736 0 _0370_
rlabel metal2 39032 27048 39032 27048 0 _0371_
rlabel metal3 36512 23800 36512 23800 0 _0372_
rlabel metal2 37800 24248 37800 24248 0 _0373_
rlabel metal2 36568 23184 36568 23184 0 _0374_
rlabel metal3 34944 24808 34944 24808 0 _0375_
rlabel metal2 35560 25816 35560 25816 0 _0376_
rlabel metal2 36120 23520 36120 23520 0 _0377_
rlabel metal2 36232 22512 36232 22512 0 _0378_
rlabel metal2 37464 24304 37464 24304 0 _0379_
rlabel metal2 33880 24920 33880 24920 0 _0380_
rlabel metal2 35616 23128 35616 23128 0 _0381_
rlabel metal2 36232 25200 36232 25200 0 _0382_
rlabel metal2 36120 26684 36120 26684 0 _0383_
rlabel metal2 32536 31696 32536 31696 0 _0384_
rlabel metal2 33096 25984 33096 25984 0 _0385_
rlabel metal2 33096 25144 33096 25144 0 _0386_
rlabel metal2 33656 25816 33656 25816 0 _0387_
rlabel metal2 33880 24024 33880 24024 0 _0388_
rlabel metal2 34216 25144 34216 25144 0 _0389_
rlabel metal2 14000 42728 14000 42728 0 _0390_
rlabel metal3 31976 27048 31976 27048 0 _0391_
rlabel metal2 32200 28392 32200 28392 0 _0392_
rlabel metal2 33824 27608 33824 27608 0 _0393_
rlabel metal2 33656 28952 33656 28952 0 _0394_
rlabel metal2 32984 27384 32984 27384 0 _0395_
rlabel metal2 34328 27720 34328 27720 0 _0396_
rlabel metal3 34664 29400 34664 29400 0 _0397_
rlabel metal3 32704 29400 32704 29400 0 _0398_
rlabel metal2 31976 30072 31976 30072 0 _0399_
rlabel metal2 33432 29344 33432 29344 0 _0400_
rlabel metal2 34888 29400 34888 29400 0 _0401_
rlabel metal2 34384 29288 34384 29288 0 _0402_
rlabel metal3 45808 43400 45808 43400 0 _0403_
rlabel metal2 19768 49840 19768 49840 0 _0404_
rlabel metal2 21112 49616 21112 49616 0 _0405_
rlabel metal2 34664 47768 34664 47768 0 _0406_
rlabel metal2 28616 35728 28616 35728 0 _0407_
rlabel metal2 21896 46256 21896 46256 0 _0408_
rlabel metal2 20664 52640 20664 52640 0 _0409_
rlabel metal3 25984 42728 25984 42728 0 _0410_
rlabel metal2 24360 45472 24360 45472 0 _0411_
rlabel metal3 17640 46088 17640 46088 0 _0412_
rlabel metal2 29512 30464 29512 30464 0 _0413_
rlabel metal2 28896 30184 28896 30184 0 _0414_
rlabel metal2 29512 49056 29512 49056 0 _0415_
rlabel metal2 22344 46368 22344 46368 0 _0416_
rlabel metal3 23744 48216 23744 48216 0 _0417_
rlabel metal2 26488 48328 26488 48328 0 _0418_
rlabel metal2 23464 46592 23464 46592 0 _0419_
rlabel metal3 15344 49560 15344 49560 0 _0420_
rlabel metal3 18872 50344 18872 50344 0 _0421_
rlabel metal2 16632 51800 16632 51800 0 _0422_
rlabel metal2 15904 45752 15904 45752 0 _0423_
rlabel metal2 23576 44632 23576 44632 0 _0424_
rlabel metal2 22288 45640 22288 45640 0 _0425_
rlabel metal2 22232 43960 22232 43960 0 _0426_
rlabel metal2 28504 46480 28504 46480 0 _0427_
rlabel metal3 28392 47432 28392 47432 0 _0428_
rlabel metal3 29008 48776 29008 48776 0 _0429_
rlabel metal3 28504 49000 28504 49000 0 _0430_
rlabel metal3 32536 45752 32536 45752 0 _0431_
rlabel metal3 28952 46760 28952 46760 0 _0432_
rlabel metal2 28952 46928 28952 46928 0 _0433_
rlabel metal2 23576 47432 23576 47432 0 _0434_
rlabel metal2 24360 47824 24360 47824 0 _0435_
rlabel metal2 27608 48496 27608 48496 0 _0436_
rlabel metal2 27888 48440 27888 48440 0 _0437_
rlabel metal2 28840 47208 28840 47208 0 _0438_
rlabel metal2 28224 46760 28224 46760 0 _0439_
rlabel metal3 30744 45192 30744 45192 0 _0440_
rlabel metal2 29624 46928 29624 46928 0 _0441_
rlabel metal2 19712 46872 19712 46872 0 _0442_
rlabel metal2 22904 44408 22904 44408 0 _0443_
rlabel metal2 21784 40656 21784 40656 0 _0444_
rlabel metal3 22792 41272 22792 41272 0 _0445_
rlabel metal2 23128 41048 23128 41048 0 _0446_
rlabel metal2 28672 40600 28672 40600 0 _0447_
rlabel metal2 34216 39592 34216 39592 0 _0448_
rlabel metal2 30072 46144 30072 46144 0 _0449_
rlabel metal2 31080 45808 31080 45808 0 _0450_
rlabel metal2 32536 46144 32536 46144 0 _0451_
rlabel metal2 29624 44744 29624 44744 0 _0452_
rlabel metal2 31192 43344 31192 43344 0 _0453_
rlabel metal2 26600 46648 26600 46648 0 _0454_
rlabel metal2 27384 46928 27384 46928 0 _0455_
rlabel metal2 28168 47096 28168 47096 0 _0456_
rlabel metal2 30408 41608 30408 41608 0 _0457_
rlabel metal2 30520 41020 30520 41020 0 _0458_
rlabel metal2 30520 35112 30520 35112 0 _0459_
rlabel metal2 28168 39928 28168 39928 0 _0460_
rlabel metal2 29400 40880 29400 40880 0 _0461_
rlabel metal2 26656 37912 26656 37912 0 _0462_
rlabel metal3 25984 39592 25984 39592 0 _0463_
rlabel metal2 23800 43176 23800 43176 0 _0464_
rlabel metal2 27160 40488 27160 40488 0 _0465_
rlabel metal2 26824 40600 26824 40600 0 _0466_
rlabel metal2 26488 41160 26488 41160 0 _0467_
rlabel metal2 25704 45360 25704 45360 0 _0468_
rlabel metal2 12600 44688 12600 44688 0 _0469_
rlabel metal2 14728 45528 14728 45528 0 _0470_
rlabel metal2 25928 45696 25928 45696 0 _0471_
rlabel metal2 26096 44184 26096 44184 0 _0472_
rlabel metal2 25592 43260 25592 43260 0 _0473_
rlabel metal2 24248 43960 24248 43960 0 _0474_
rlabel metal2 31416 46032 31416 46032 0 _0475_
rlabel metal2 26768 44184 26768 44184 0 _0476_
rlabel metal2 26600 42504 26600 42504 0 _0477_
rlabel metal2 29400 39592 29400 39592 0 _0478_
rlabel metal2 29568 35112 29568 35112 0 _0479_
rlabel metal3 16520 46760 16520 46760 0 _0480_
rlabel metal2 23408 46088 23408 46088 0 _0481_
rlabel metal2 29736 41048 29736 41048 0 _0482_
rlabel metal2 30072 40040 30072 40040 0 _0483_
rlabel metal3 29624 43512 29624 43512 0 _0484_
rlabel metal2 32536 39928 32536 39928 0 _0485_
rlabel metal2 22568 41440 22568 41440 0 _0486_
rlabel metal2 32872 40488 32872 40488 0 _0487_
rlabel metal2 32984 39480 32984 39480 0 _0488_
rlabel metal2 33320 42000 33320 42000 0 _0489_
rlabel metal3 30296 39816 30296 39816 0 _0490_
rlabel metal2 29344 39032 29344 39032 0 _0491_
rlabel metal3 23744 46648 23744 46648 0 _0492_
rlabel metal2 25032 46144 25032 46144 0 _0493_
rlabel metal2 25872 45192 25872 45192 0 _0494_
rlabel metal2 29288 45024 29288 45024 0 _0495_
rlabel metal2 18984 43624 18984 43624 0 _0496_
rlabel metal3 29008 42056 29008 42056 0 _0497_
rlabel metal2 26712 42056 26712 42056 0 _0498_
rlabel metal2 33768 39200 33768 39200 0 _0499_
rlabel metal2 33768 37072 33768 37072 0 _0500_
rlabel metal2 26264 40824 26264 40824 0 _0501_
rlabel metal2 26824 41496 26824 41496 0 _0502_
rlabel metal2 31864 41608 31864 41608 0 _0503_
rlabel metal2 26376 45920 26376 45920 0 _0504_
rlabel metal3 30520 44072 30520 44072 0 _0505_
rlabel metal2 30968 44744 30968 44744 0 _0506_
rlabel metal2 34664 44800 34664 44800 0 _0507_
rlabel metal2 26768 45864 26768 45864 0 _0508_
rlabel metal2 31640 44464 31640 44464 0 _0509_
rlabel metal2 33768 44352 33768 44352 0 _0510_
rlabel metal2 34440 43960 34440 43960 0 _0511_
rlabel metal3 29792 44296 29792 44296 0 _0512_
rlabel metal2 31360 40488 31360 40488 0 _0513_
rlabel metal3 35392 40600 35392 40600 0 _0514_
rlabel metal3 36288 42056 36288 42056 0 _0515_
rlabel metal2 38248 40600 38248 40600 0 _0516_
rlabel metal3 27944 42168 27944 42168 0 _0517_
rlabel metal2 28728 43456 28728 43456 0 _0518_
rlabel metal2 28840 42504 28840 42504 0 _0519_
rlabel metal2 28840 41720 28840 41720 0 _0520_
rlabel metal2 35784 41496 35784 41496 0 _0521_
rlabel metal3 15736 44184 15736 44184 0 _0522_
rlabel metal2 35336 41272 35336 41272 0 _0523_
rlabel metal2 29512 42784 29512 42784 0 _0524_
rlabel metal3 25732 43400 25732 43400 0 _0525_
rlabel metal2 28280 43120 28280 43120 0 _0526_
rlabel metal2 34552 43120 34552 43120 0 _0527_
rlabel metal3 35504 41944 35504 41944 0 _0528_
rlabel metal2 30632 43232 30632 43232 0 _0529_
rlabel metal2 27608 46144 27608 46144 0 _0530_
rlabel metal2 30072 43456 30072 43456 0 _0531_
rlabel metal2 31640 42392 31640 42392 0 _0532_
rlabel metal3 32648 41720 32648 41720 0 _0533_
rlabel metal2 14840 42280 14840 42280 0 _0534_
rlabel metal2 18928 42952 18928 42952 0 _0535_
rlabel metal2 17304 44128 17304 44128 0 _0536_
rlabel metal2 18984 45472 18984 45472 0 _0537_
rlabel metal2 14504 44128 14504 44128 0 _0538_
rlabel metal3 13496 42728 13496 42728 0 _0539_
rlabel metal3 6720 50344 6720 50344 0 _0540_
rlabel metal2 6944 47208 6944 47208 0 _0541_
rlabel metal2 3304 52864 3304 52864 0 _0542_
rlabel metal2 6160 49224 6160 49224 0 _0543_
rlabel metal2 6272 39816 6272 39816 0 _0544_
rlabel metal2 6552 44296 6552 44296 0 _0545_
rlabel metal2 5152 43736 5152 43736 0 _0546_
rlabel metal2 5656 45584 5656 45584 0 _0547_
rlabel metal3 7560 45192 7560 45192 0 _0548_
rlabel metal2 10360 43736 10360 43736 0 _0549_
rlabel metal2 12712 43344 12712 43344 0 _0550_
rlabel metal2 13384 42616 13384 42616 0 _0551_
rlabel metal2 11816 43680 11816 43680 0 _0552_
rlabel metal3 13104 44072 13104 44072 0 _0553_
rlabel metal3 16856 42840 16856 42840 0 _0554_
rlabel metal3 20384 40936 20384 40936 0 _0555_
rlabel metal2 18088 42504 18088 42504 0 _0556_
rlabel metal3 13440 43512 13440 43512 0 _0557_
rlabel metal2 12264 43596 12264 43596 0 _0558_
rlabel metal3 9520 47992 9520 47992 0 _0559_
rlabel metal3 12208 44296 12208 44296 0 _0560_
rlabel metal2 18200 44184 18200 44184 0 _0561_
rlabel metal2 16576 44408 16576 44408 0 _0562_
rlabel metal2 11872 51128 11872 51128 0 _0563_
rlabel metal3 9352 48104 9352 48104 0 _0564_
rlabel metal2 10584 49560 10584 49560 0 _0565_
rlabel metal2 14616 42840 14616 42840 0 _0566_
rlabel metal2 13664 51128 13664 51128 0 _0567_
rlabel metal2 10752 49784 10752 49784 0 _0568_
rlabel metal2 10584 52024 10584 52024 0 _0569_
rlabel metal3 11704 51128 11704 51128 0 _0570_
rlabel metal3 11480 52808 11480 52808 0 _0571_
rlabel metal3 17024 42728 17024 42728 0 _0572_
rlabel metal2 13720 52976 13720 52976 0 _0573_
rlabel metal2 12936 53480 12936 53480 0 _0574_
rlabel metal2 13720 51352 13720 51352 0 _0575_
rlabel metal2 14392 51632 14392 51632 0 _0576_
rlabel metal2 17864 50204 17864 50204 0 _0577_
rlabel metal2 17808 43624 17808 43624 0 _0578_
rlabel metal2 17304 49840 17304 49840 0 _0579_
rlabel metal2 17752 49000 17752 49000 0 _0580_
rlabel metal3 16016 39592 16016 39592 0 _0581_
rlabel metal4 16072 47712 16072 47712 0 _0582_
rlabel metal2 15848 52080 15848 52080 0 _0583_
rlabel metal3 6104 48216 6104 48216 0 _0584_
rlabel metal2 3080 48272 3080 48272 0 _0585_
rlabel metal2 2800 54488 2800 54488 0 _0586_
rlabel metal2 4872 51128 4872 51128 0 _0587_
rlabel metal2 6832 52136 6832 52136 0 _0588_
rlabel metal2 4200 52640 4200 52640 0 _0589_
rlabel metal2 7168 54488 7168 54488 0 _0590_
rlabel metal3 5040 50568 5040 50568 0 _0591_
rlabel metal2 7112 51240 7112 51240 0 _0592_
rlabel metal3 6888 49000 6888 49000 0 _0593_
rlabel metal2 4312 49000 4312 49000 0 _0594_
rlabel metal2 7224 49224 7224 49224 0 _0595_
rlabel metal2 6496 48776 6496 48776 0 _0596_
rlabel metal3 4480 43512 4480 43512 0 _0597_
rlabel metal2 5768 44464 5768 44464 0 _0598_
rlabel metal2 7560 43120 7560 43120 0 _0599_
rlabel metal2 6216 39200 6216 39200 0 _0600_
rlabel metal2 6720 38920 6720 38920 0 _0601_
rlabel metal2 3304 44800 3304 44800 0 _0602_
rlabel metal2 7560 38668 7560 38668 0 _0603_
rlabel metal2 5208 39144 5208 39144 0 _0604_
rlabel metal2 4088 37352 4088 37352 0 _0605_
rlabel metal2 5656 41552 5656 41552 0 _0606_
rlabel metal2 4368 39592 4368 39592 0 _0607_
rlabel metal3 6608 41160 6608 41160 0 _0608_
rlabel metal3 4424 41944 4424 41944 0 _0609_
rlabel metal2 3808 42952 3808 42952 0 _0610_
rlabel metal3 3584 41832 3584 41832 0 _0611_
rlabel metal2 3920 44520 3920 44520 0 _0612_
rlabel metal2 2296 44744 2296 44744 0 _0613_
rlabel metal2 2856 44800 2856 44800 0 _0614_
rlabel metal2 3584 46648 3584 46648 0 _0615_
rlabel metal2 2576 46760 2576 46760 0 _0616_
rlabel metal2 27216 28504 27216 28504 0 _0617_
rlabel metal2 22344 26432 22344 26432 0 _0618_
rlabel metal3 24752 26264 24752 26264 0 _0619_
rlabel metal2 27608 29008 27608 29008 0 _0620_
rlabel metal3 24640 26152 24640 26152 0 _0621_
rlabel metal3 21168 26488 21168 26488 0 _0622_
rlabel metal2 22008 25088 22008 25088 0 _0623_
rlabel metal2 22792 26544 22792 26544 0 _0624_
rlabel metal2 21336 27888 21336 27888 0 _0625_
rlabel metal3 21560 27048 21560 27048 0 _0626_
rlabel metal2 19656 27384 19656 27384 0 _0627_
rlabel metal2 20776 26320 20776 26320 0 _0628_
rlabel metal2 20888 25480 20888 25480 0 _0629_
rlabel metal2 25424 40712 25424 40712 0 _0630_
rlabel metal2 24752 50456 24752 50456 0 _0631_
rlabel metal2 22680 41272 22680 41272 0 _0632_
rlabel metal2 24584 51856 24584 51856 0 _0633_
rlabel metal2 22344 49784 22344 49784 0 _0634_
rlabel metal2 19600 42056 19600 42056 0 _0635_
rlabel metal3 21784 41720 21784 41720 0 _0636_
rlabel metal2 20664 47712 20664 47712 0 _0637_
rlabel metal2 20328 49784 20328 49784 0 _0638_
rlabel metal2 21336 48944 21336 48944 0 _0639_
rlabel metal3 21560 49560 21560 49560 0 _0640_
rlabel metal3 22960 50568 22960 50568 0 _0641_
rlabel metal2 26376 43176 26376 43176 0 _0642_
rlabel metal2 23688 47544 23688 47544 0 _0643_
rlabel metal2 23464 50568 23464 50568 0 _0644_
rlabel metal2 22904 49840 22904 49840 0 _0645_
rlabel metal2 22736 48776 22736 48776 0 _0646_
rlabel metal2 25368 41664 25368 41664 0 _0647_
rlabel metal2 24136 49504 24136 49504 0 _0648_
rlabel metal2 25144 40040 25144 40040 0 _0649_
rlabel metal3 24472 48888 24472 48888 0 _0650_
rlabel metal2 22624 49224 22624 49224 0 _0651_
rlabel metal3 21336 49672 21336 49672 0 _0652_
rlabel metal2 23128 50008 23128 50008 0 _0653_
rlabel metal2 23800 53872 23800 53872 0 _0654_
rlabel metal2 24192 49000 24192 49000 0 _0655_
rlabel metal2 24080 51688 24080 51688 0 _0656_
rlabel metal3 19432 50904 19432 50904 0 _0657_
rlabel metal3 21112 51240 21112 51240 0 _0658_
rlabel metal2 22232 52248 22232 52248 0 _0659_
rlabel metal2 23968 53144 23968 53144 0 _0660_
rlabel metal2 24248 50960 24248 50960 0 _0661_
rlabel metal3 19992 50624 19992 50624 0 _0662_
rlabel metal2 23800 51632 23800 51632 0 _0663_
rlabel metal3 24920 52248 24920 52248 0 _0664_
rlabel metal3 32928 15288 32928 15288 0 _0665_
rlabel metal2 34776 16016 34776 16016 0 _0666_
rlabel metal2 34104 16296 34104 16296 0 _0667_
rlabel metal2 35728 11592 35728 11592 0 _0668_
rlabel metal2 36064 16072 36064 16072 0 _0669_
rlabel metal3 19712 15960 19712 15960 0 _0670_
rlabel metal2 19768 13496 19768 13496 0 _0671_
rlabel metal2 18088 13048 18088 13048 0 _0672_
rlabel metal2 14448 12824 14448 12824 0 _0673_
rlabel metal2 16520 12936 16520 12936 0 _0674_
rlabel metal2 12936 12880 12936 12880 0 _0675_
rlabel metal3 11312 12152 11312 12152 0 _0676_
rlabel metal2 10920 12488 10920 12488 0 _0677_
rlabel metal2 23464 21672 23464 21672 0 _0678_
rlabel metal2 30632 11368 30632 11368 0 _0679_
rlabel metal2 31080 9856 31080 9856 0 _0680_
rlabel metal2 30016 9800 30016 9800 0 _0681_
rlabel metal2 22176 21560 22176 21560 0 _0682_
rlabel metal2 23072 20104 23072 20104 0 _0683_
rlabel metal2 20552 16128 20552 16128 0 _0684_
rlabel metal2 19544 16912 19544 16912 0 _0685_
rlabel metal3 20776 15288 20776 15288 0 _0686_
rlabel metal2 22736 20888 22736 20888 0 _0687_
rlabel metal2 31528 13832 31528 13832 0 _0688_
rlabel metal2 30856 15512 30856 15512 0 _0689_
rlabel metal2 30408 13832 30408 13832 0 _0690_
rlabel metal2 33880 11312 33880 11312 0 _0691_
rlabel metal2 33320 12264 33320 12264 0 _0692_
rlabel metal2 35672 10920 35672 10920 0 _0693_
rlabel metal2 12264 15624 12264 15624 0 _0694_
rlabel metal2 10584 14280 10584 14280 0 _0695_
rlabel metal3 9968 15848 9968 15848 0 _0696_
rlabel metal2 34104 20104 34104 20104 0 _0697_
rlabel metal2 29512 20048 29512 20048 0 _0698_
rlabel metal3 28000 20104 28000 20104 0 _0699_
rlabel metal2 36008 20552 36008 20552 0 _0700_
rlabel metal2 30744 19712 30744 19712 0 _0701_
rlabel metal3 25788 21672 25788 21672 0 _0702_
rlabel metal2 32760 21560 32760 21560 0 _0703_
rlabel metal2 35112 21280 35112 21280 0 _0704_
rlabel metal2 26600 6104 26600 6104 0 _0705_
rlabel metal2 24248 6216 24248 6216 0 _0706_
rlabel metal2 20552 5376 20552 5376 0 _0707_
rlabel metal2 23744 8232 23744 8232 0 _0708_
rlabel metal2 21560 5208 21560 5208 0 _0709_
rlabel metal2 27608 6272 27608 6272 0 _0710_
rlabel metal2 26264 4032 26264 4032 0 _0711_
rlabel metal2 26936 6328 26936 6328 0 _0712_
rlabel metal2 22456 9016 22456 9016 0 _0713_
rlabel metal2 20440 8512 20440 8512 0 _0714_
rlabel metal3 24360 8232 24360 8232 0 _0715_
rlabel metal2 27384 8680 27384 8680 0 _0716_
rlabel metal2 26488 10192 26488 10192 0 _0717_
rlabel metal2 26824 8176 26824 8176 0 _0718_
rlabel metal2 28504 22288 28504 22288 0 _0719_
rlabel metal2 26936 21504 26936 21504 0 _0720_
rlabel metal2 29288 22848 29288 22848 0 _0721_
rlabel metal2 25592 18760 25592 18760 0 _0722_
rlabel metal2 33768 18760 33768 18760 0 _0723_
rlabel metal2 33320 18312 33320 18312 0 _0724_
rlabel metal2 35896 18312 35896 18312 0 _0725_
rlabel metal2 8232 26376 8232 26376 0 _0726_
rlabel metal2 5992 27328 5992 27328 0 _0727_
rlabel metal2 7336 28616 7336 28616 0 _0728_
rlabel metal2 40096 51464 40096 51464 0 _0729_
rlabel metal2 49336 46368 49336 46368 0 _0730_
rlabel metal2 47544 51240 47544 51240 0 _0731_
rlabel metal3 48216 49896 48216 49896 0 _0732_
rlabel metal3 46536 49784 46536 49784 0 _0733_
rlabel metal2 43624 50176 43624 50176 0 _0734_
rlabel metal2 48104 51240 48104 51240 0 _0735_
rlabel metal2 46592 50568 46592 50568 0 _0736_
rlabel metal2 42952 51072 42952 51072 0 _0737_
rlabel metal2 49336 51240 49336 51240 0 _0738_
rlabel metal2 48216 50848 48216 50848 0 _0739_
rlabel metal2 43288 49952 43288 49952 0 _0740_
rlabel metal2 42280 51240 42280 51240 0 _0741_
rlabel metal2 42056 51800 42056 51800 0 _0742_
rlabel metal3 40236 52248 40236 52248 0 _0743_
rlabel metal2 40040 49896 40040 49896 0 _0744_
rlabel metal2 44072 49700 44072 49700 0 _0745_
rlabel metal2 41832 49392 41832 49392 0 _0746_
rlabel metal2 39144 49840 39144 49840 0 _0747_
rlabel metal2 40264 53088 40264 53088 0 _0748_
rlabel metal2 42672 50792 42672 50792 0 _0749_
rlabel metal3 43064 50008 43064 50008 0 _0750_
rlabel metal3 36904 49784 36904 49784 0 _0751_
rlabel metal2 42224 48888 42224 48888 0 _0752_
rlabel metal2 39368 50568 39368 50568 0 _0753_
rlabel metal2 41272 52752 41272 52752 0 _0754_
rlabel metal2 41888 49000 41888 49000 0 _0755_
rlabel metal2 41384 49280 41384 49280 0 _0756_
rlabel metal2 41272 49728 41272 49728 0 _0757_
rlabel metal2 39200 50120 39200 50120 0 _0758_
rlabel metal2 38976 49224 38976 49224 0 _0759_
rlabel metal2 39704 50344 39704 50344 0 _0760_
rlabel metal3 37128 50232 37128 50232 0 _0761_
rlabel metal2 38136 52976 38136 52976 0 _0762_
rlabel metal2 38696 50960 38696 50960 0 _0763_
rlabel metal2 38920 52920 38920 52920 0 _0764_
rlabel metal2 37912 53200 37912 53200 0 _0765_
rlabel metal2 38752 49560 38752 49560 0 _0766_
rlabel metal3 41552 52920 41552 52920 0 _0767_
rlabel metal2 39256 52024 39256 52024 0 _0768_
rlabel metal3 38248 51576 38248 51576 0 _0769_
rlabel metal3 39592 52024 39592 52024 0 _0770_
rlabel metal2 39368 52920 39368 52920 0 _0771_
rlabel metal2 39032 51576 39032 51576 0 _0772_
rlabel metal3 38080 52248 38080 52248 0 _0773_
rlabel metal3 34776 52920 34776 52920 0 _0774_
rlabel metal2 38024 52976 38024 52976 0 _0775_
rlabel metal2 36008 52752 36008 52752 0 _0776_
rlabel metal2 34328 53480 34328 53480 0 _0777_
rlabel metal2 39704 53928 39704 53928 0 _0778_
rlabel metal3 37072 48776 37072 48776 0 _0779_
rlabel metal3 40040 50568 40040 50568 0 _0780_
rlabel metal2 34664 50008 34664 50008 0 _0781_
rlabel metal2 36232 53200 36232 53200 0 _0782_
rlabel metal2 42392 49672 42392 49672 0 _0783_
rlabel metal2 36120 49392 36120 49392 0 _0784_
rlabel metal2 36456 52304 36456 52304 0 _0785_
rlabel metal2 36904 53592 36904 53592 0 _0786_
rlabel metal2 18312 40880 18312 40880 0 _0787_
rlabel metal3 30296 37912 30296 37912 0 _0788_
rlabel metal3 32144 36232 32144 36232 0 _0789_
rlabel metal2 45472 42504 45472 42504 0 _0790_
rlabel metal2 19992 41496 19992 41496 0 _0791_
rlabel metal2 22904 40656 22904 40656 0 _0792_
rlabel metal2 13440 47432 13440 47432 0 _0793_
rlabel metal2 16072 46816 16072 46816 0 _0794_
rlabel metal3 18704 51128 18704 51128 0 _0795_
rlabel metal3 18760 49896 18760 49896 0 _0796_
rlabel metal2 15960 49112 15960 49112 0 _0797_
rlabel metal2 15512 46368 15512 46368 0 _0798_
rlabel metal2 15176 46424 15176 46424 0 _0799_
rlabel metal2 15736 46928 15736 46928 0 _0800_
rlabel metal3 21896 47208 21896 47208 0 _0801_
rlabel metal2 14056 46928 14056 46928 0 _0802_
rlabel metal2 15064 51464 15064 51464 0 _0803_
rlabel metal3 13496 52136 13496 52136 0 _0804_
rlabel metal2 12600 48552 12600 48552 0 _0805_
rlabel metal2 16072 40600 16072 40600 0 _0806_
rlabel metal3 34104 48888 34104 48888 0 _0807_
rlabel metal2 21560 45472 21560 45472 0 _0808_
rlabel metal2 21784 47040 21784 47040 0 _0809_
rlabel metal2 17864 54880 17864 54880 0 _0810_
rlabel metal2 19656 47656 19656 47656 0 _0811_
rlabel metal2 19320 47320 19320 47320 0 _0812_
rlabel metal2 17976 42000 17976 42000 0 _0813_
rlabel metal2 13496 41608 13496 41608 0 _0814_
rlabel metal2 17752 44912 17752 44912 0 _0815_
rlabel metal2 14392 50848 14392 50848 0 _0816_
rlabel metal2 12488 52584 12488 52584 0 _0817_
rlabel metal2 12936 47880 12936 47880 0 _0818_
rlabel metal2 12824 46928 12824 46928 0 _0819_
rlabel metal2 18424 48160 18424 48160 0 _0820_
rlabel metal2 25144 48160 25144 48160 0 _0821_
rlabel metal2 10696 45752 10696 45752 0 _0822_
rlabel metal3 12376 46648 12376 46648 0 _0823_
rlabel metal2 18088 45472 18088 45472 0 _0824_
rlabel metal2 30744 49448 30744 49448 0 _0825_
rlabel metal2 17752 46704 17752 46704 0 _0826_
rlabel metal3 16800 41272 16800 41272 0 _0827_
rlabel metal2 17416 38360 17416 38360 0 _0828_
rlabel metal2 16688 34216 16688 34216 0 _0829_
rlabel metal2 17864 23016 17864 23016 0 _0830_
rlabel metal2 17864 31360 17864 31360 0 _0831_
rlabel metal3 18704 30856 18704 30856 0 _0832_
rlabel metal2 16184 30856 16184 30856 0 _0833_
rlabel metal2 16856 30744 16856 30744 0 _0834_
rlabel metal2 24136 28168 24136 28168 0 _0835_
rlabel metal2 26152 30240 26152 30240 0 _0836_
rlabel metal2 24360 28336 24360 28336 0 _0837_
rlabel metal2 24584 28168 24584 28168 0 _0838_
rlabel metal2 22120 30520 22120 30520 0 _0839_
rlabel metal2 22008 30016 22008 30016 0 _0840_
rlabel metal2 22792 28952 22792 28952 0 _0841_
rlabel metal2 25368 29344 25368 29344 0 _0842_
rlabel metal3 17024 29512 17024 29512 0 _0843_
rlabel metal3 17696 30856 17696 30856 0 _0844_
rlabel metal3 16184 30072 16184 30072 0 _0845_
rlabel metal2 17416 29680 17416 29680 0 _0846_
rlabel metal2 18424 29736 18424 29736 0 _0847_
rlabel metal2 17752 34888 17752 34888 0 _0848_
rlabel metal2 16184 36624 16184 36624 0 _0849_
rlabel metal3 24360 15512 24360 15512 0 _0850_
rlabel metal2 25256 15848 25256 15848 0 _0851_
rlabel metal3 16856 15848 16856 15848 0 _0852_
rlabel metal2 25592 13944 25592 13944 0 _0853_
rlabel metal2 27384 14784 27384 14784 0 _0854_
rlabel metal2 16856 16520 16856 16520 0 _0855_
rlabel metal2 17416 16744 17416 16744 0 _0856_
rlabel metal3 24304 15176 24304 15176 0 _0857_
rlabel metal2 28616 15540 28616 15540 0 _0858_
rlabel metal2 26824 15960 26824 15960 0 _0859_
rlabel metal3 29120 16296 29120 16296 0 _0860_
rlabel metal2 16968 17696 16968 17696 0 _0861_
rlabel metal2 28056 17192 28056 17192 0 _0862_
rlabel metal2 28224 15288 28224 15288 0 _0863_
rlabel metal3 25256 16800 25256 16800 0 _0864_
rlabel metal2 27048 17360 27048 17360 0 _0865_
rlabel metal2 35168 13160 35168 13160 0 _0866_
rlabel metal2 28616 7336 28616 7336 0 _0867_
rlabel metal2 25368 11424 25368 11424 0 _0868_
rlabel metal2 29568 11144 29568 11144 0 _0869_
rlabel metal3 28728 13608 28728 13608 0 _0870_
rlabel metal2 15624 15904 15624 15904 0 _0871_
rlabel metal3 22792 12992 22792 12992 0 _0872_
rlabel metal2 27272 17304 27272 17304 0 _0873_
rlabel metal3 15624 17528 15624 17528 0 _0874_
rlabel metal2 25424 15512 25424 15512 0 _0875_
rlabel metal2 33880 15568 33880 15568 0 _0876_
rlabel metal2 28728 19152 28728 19152 0 _0877_
rlabel metal2 28168 17192 28168 17192 0 _0878_
rlabel metal3 27440 16072 27440 16072 0 _0879_
rlabel metal2 24584 15512 24584 15512 0 _0880_
rlabel metal3 23688 12376 23688 12376 0 _0881_
rlabel metal2 23016 12600 23016 12600 0 _0882_
rlabel metal2 25592 13104 25592 13104 0 _0883_
rlabel metal3 24752 12936 24752 12936 0 _0884_
rlabel metal2 24696 15204 24696 15204 0 _0885_
rlabel metal2 17528 18032 17528 18032 0 _0886_
rlabel metal3 24920 15288 24920 15288 0 _0887_
rlabel metal2 25592 15904 25592 15904 0 _0888_
rlabel metal3 13496 16856 13496 16856 0 _0889_
rlabel metal3 13216 8120 13216 8120 0 _0890_
rlabel metal3 13496 13944 13496 13944 0 _0891_
rlabel metal2 9912 17976 9912 17976 0 _0892_
rlabel metal2 11032 16576 11032 16576 0 _0893_
rlabel metal2 14616 11312 14616 11312 0 _0894_
rlabel metal2 11648 18200 11648 18200 0 _0895_
rlabel metal2 11592 18816 11592 18816 0 _0896_
rlabel metal2 12488 18312 12488 18312 0 _0897_
rlabel metal2 15288 20720 15288 20720 0 _0898_
rlabel metal2 12936 18424 12936 18424 0 _0899_
rlabel metal2 12824 10696 12824 10696 0 _0900_
rlabel metal2 6832 17080 6832 17080 0 _0901_
rlabel metal2 16184 22176 16184 22176 0 _0902_
rlabel metal3 9576 18424 9576 18424 0 _0903_
rlabel metal2 13272 17472 13272 17472 0 _0904_
rlabel metal2 13608 16464 13608 16464 0 _0905_
rlabel metal3 13664 16632 13664 16632 0 _0906_
rlabel metal2 16520 18144 16520 18144 0 _0907_
rlabel metal3 11704 8344 11704 8344 0 _0908_
rlabel metal2 9912 19040 9912 19040 0 _0909_
rlabel metal2 10360 19600 10360 19600 0 _0910_
rlabel metal2 13832 18704 13832 18704 0 _0911_
rlabel metal2 14728 18928 14728 18928 0 _0912_
rlabel metal2 15176 16856 15176 16856 0 _0913_
rlabel metal3 13272 20776 13272 20776 0 _0914_
rlabel metal3 8568 17528 8568 17528 0 _0915_
rlabel metal2 9576 24276 9576 24276 0 _0916_
rlabel metal2 9968 21560 9968 21560 0 _0917_
rlabel metal2 8904 21616 8904 21616 0 _0918_
rlabel metal2 12376 21224 12376 21224 0 _0919_
rlabel metal2 14504 19320 14504 19320 0 _0920_
rlabel metal3 15400 19208 15400 19208 0 _0921_
rlabel metal2 16744 19320 16744 19320 0 _0922_
rlabel metal2 26656 37128 26656 37128 0 _0923_
rlabel metal2 24976 37240 24976 37240 0 _0924_
rlabel metal2 25816 16240 25816 16240 0 _0925_
rlabel metal3 28392 15400 28392 15400 0 _0926_
rlabel metal2 22008 12768 22008 12768 0 _0927_
rlabel metal2 27608 12264 27608 12264 0 _0928_
rlabel metal2 21224 18536 21224 18536 0 _0929_
rlabel metal2 27328 16744 27328 16744 0 _0930_
rlabel metal2 24696 17472 24696 17472 0 _0931_
rlabel metal2 26992 16296 26992 16296 0 _0932_
rlabel metal2 26152 15736 26152 15736 0 _0933_
rlabel metal3 26852 13720 26852 13720 0 _0934_
rlabel metal2 26320 6104 26320 6104 0 _0935_
rlabel metal2 27664 13160 27664 13160 0 _0936_
rlabel metal2 26936 13272 26936 13272 0 _0937_
rlabel metal2 26488 15848 26488 15848 0 _0938_
rlabel metal2 26264 16576 26264 16576 0 _0939_
rlabel metal3 28672 16968 28672 16968 0 _0940_
rlabel metal2 25368 18592 25368 18592 0 _0941_
rlabel metal2 24920 18032 24920 18032 0 _0942_
rlabel metal2 25592 16520 25592 16520 0 _0943_
rlabel metal2 24360 16632 24360 16632 0 _0944_
rlabel metal2 23464 6664 23464 6664 0 _0945_
rlabel metal2 21672 12600 21672 12600 0 _0946_
rlabel metal3 21504 13160 21504 13160 0 _0947_
rlabel metal2 22456 12936 22456 12936 0 _0948_
rlabel metal3 23800 13832 23800 13832 0 _0949_
rlabel metal2 24248 16408 24248 16408 0 _0950_
rlabel metal2 25816 19320 25816 19320 0 _0951_
rlabel metal3 11928 16296 11928 16296 0 _0952_
rlabel metal2 11368 18088 11368 18088 0 _0953_
rlabel metal3 12656 19768 12656 19768 0 _0954_
rlabel metal2 11928 19488 11928 19488 0 _0955_
rlabel metal3 12264 17864 12264 17864 0 _0956_
rlabel metal2 12936 17584 12936 17584 0 _0957_
rlabel metal2 15120 11592 15120 11592 0 _0958_
rlabel metal2 6440 17304 6440 17304 0 _0959_
rlabel metal2 7784 16968 7784 16968 0 _0960_
rlabel metal3 11368 17416 11368 17416 0 _0961_
rlabel metal3 14952 17640 14952 17640 0 _0962_
rlabel metal2 15792 17864 15792 17864 0 _0963_
rlabel metal2 14952 6216 14952 6216 0 _0964_
rlabel metal2 9128 22232 9128 22232 0 _0965_
rlabel metal3 8288 21000 8288 21000 0 _0966_
rlabel metal2 14616 19880 14616 19880 0 _0967_
rlabel metal3 15400 19992 15400 19992 0 _0968_
rlabel metal2 14952 22232 14952 22232 0 _0969_
rlabel metal2 7672 26544 7672 26544 0 _0970_
rlabel metal3 8288 21448 8288 21448 0 _0971_
rlabel metal3 11704 21000 11704 21000 0 _0972_
rlabel metal2 15512 20048 15512 20048 0 _0973_
rlabel metal2 16072 19600 16072 19600 0 _0974_
rlabel metal2 16408 19040 16408 19040 0 _0975_
rlabel metal2 26264 38696 26264 38696 0 _0976_
rlabel metal2 24360 37632 24360 37632 0 _0977_
rlabel metal3 21784 35784 21784 35784 0 _0978_
rlabel metal3 20384 37240 20384 37240 0 _0979_
rlabel metal2 12936 51408 12936 51408 0 _0980_
rlabel metal2 13832 49728 13832 49728 0 _0981_
rlabel metal2 14168 49336 14168 49336 0 _0982_
rlabel metal3 17640 47432 17640 47432 0 _0983_
rlabel metal2 22456 40544 22456 40544 0 _0984_
rlabel metal2 18704 37016 18704 37016 0 _0985_
rlabel metal2 16688 39592 16688 39592 0 _0986_
rlabel metal2 16464 35448 16464 35448 0 _0987_
rlabel metal2 31304 38724 31304 38724 0 _0988_
rlabel metal2 22624 37800 22624 37800 0 _0989_
rlabel metal3 22456 41944 22456 41944 0 _0990_
rlabel metal2 22008 42504 22008 42504 0 _0991_
rlabel metal2 23128 39312 23128 39312 0 _0992_
rlabel metal2 18592 41720 18592 41720 0 _0993_
rlabel metal3 22344 45864 22344 45864 0 _0994_
rlabel metal2 22288 40936 22288 40936 0 _0995_
rlabel metal2 18984 36176 18984 36176 0 _0996_
rlabel metal2 19936 36456 19936 36456 0 _0997_
rlabel metal2 16520 38976 16520 38976 0 _0998_
rlabel metal2 20552 38864 20552 38864 0 _0999_
rlabel metal2 19768 41104 19768 41104 0 _1000_
rlabel metal2 22792 47600 22792 47600 0 _1001_
rlabel metal2 14952 42952 14952 42952 0 _1002_
rlabel metal2 15288 41552 15288 41552 0 _1003_
rlabel metal3 18480 40152 18480 40152 0 _1004_
rlabel metal2 16184 39312 16184 39312 0 _1005_
rlabel metal3 25256 35896 25256 35896 0 _1006_
rlabel metal2 19096 32760 19096 32760 0 _1007_
rlabel metal2 25032 40264 25032 40264 0 _1008_
rlabel metal2 23464 36344 23464 36344 0 _1009_
rlabel metal2 18760 43344 18760 43344 0 _1010_
rlabel metal2 23576 42896 23576 42896 0 _1011_
rlabel metal2 17416 54544 17416 54544 0 _1012_
rlabel metal2 16912 54712 16912 54712 0 _1013_
rlabel metal2 19712 54600 19712 54600 0 _1014_
rlabel metal3 18592 54712 18592 54712 0 _1015_
rlabel metal2 17864 42672 17864 42672 0 _1016_
rlabel metal2 17360 41944 17360 41944 0 _1017_
rlabel metal3 17696 45752 17696 45752 0 _1018_
rlabel metal2 24024 43120 24024 43120 0 _1019_
rlabel metal2 16520 39368 16520 39368 0 _1020_
rlabel metal2 20664 45920 20664 45920 0 _1021_
rlabel metal3 19040 45864 19040 45864 0 _1022_
rlabel metal3 19096 42952 19096 42952 0 _1023_
rlabel metal2 15624 39200 15624 39200 0 _1024_
rlabel metal2 15400 39312 15400 39312 0 _1025_
rlabel metal2 15176 43680 15176 43680 0 _1026_
rlabel metal2 15288 42896 15288 42896 0 _1027_
rlabel metal2 16856 40600 16856 40600 0 _1028_
rlabel metal2 14784 38808 14784 38808 0 _1029_
rlabel metal2 15288 38724 15288 38724 0 _1030_
rlabel metal3 17248 36456 17248 36456 0 _1031_
rlabel metal2 13664 34776 13664 34776 0 _1032_
rlabel metal3 17360 38696 17360 38696 0 _1033_
rlabel metal2 17416 41216 17416 41216 0 _1034_
rlabel metal2 14616 36456 14616 36456 0 _1035_
rlabel metal2 14168 36288 14168 36288 0 _1036_
rlabel metal2 43064 53312 43064 53312 0 _1037_
rlabel metal3 36288 51464 36288 51464 0 _1038_
rlabel metal2 34776 50792 34776 50792 0 _1039_
rlabel metal3 34888 50568 34888 50568 0 _1040_
rlabel metal2 35056 50792 35056 50792 0 _1041_
rlabel metal2 34664 51072 34664 51072 0 _1042_
rlabel metal2 39816 53480 39816 53480 0 _1043_
rlabel metal2 38752 52920 38752 52920 0 _1044_
rlabel metal2 39536 53144 39536 53144 0 _1045_
rlabel metal2 35224 53256 35224 53256 0 _1046_
rlabel metal2 34776 53368 34776 53368 0 _1047_
rlabel metal2 29288 30576 29288 30576 0 _1048_
rlabel metal2 17416 37576 17416 37576 0 _1049_
rlabel metal3 18928 38808 18928 38808 0 _1050_
rlabel metal2 21896 40096 21896 40096 0 _1051_
rlabel metal2 19208 40376 19208 40376 0 _1052_
rlabel metal2 19432 43204 19432 43204 0 _1053_
rlabel metal2 19656 40320 19656 40320 0 _1054_
rlabel metal3 15064 39480 15064 39480 0 _1055_
rlabel metal2 18088 38024 18088 38024 0 _1056_
rlabel metal2 20328 25424 20328 25424 0 _1057_
rlabel metal2 20552 34328 20552 34328 0 _1058_
rlabel metal3 28616 26264 28616 26264 0 _1059_
rlabel metal3 16072 24696 16072 24696 0 _1060_
rlabel metal2 15512 25256 15512 25256 0 _1061_
rlabel metal2 23576 25536 23576 25536 0 _1062_
rlabel metal2 25592 23128 25592 23128 0 _1063_
rlabel metal3 25088 23912 25088 23912 0 _1064_
rlabel metal2 19880 21728 19880 21728 0 _1065_
rlabel metal2 25816 23576 25816 23576 0 _1066_
rlabel metal2 26152 21112 26152 21112 0 _1067_
rlabel metal2 20552 21728 20552 21728 0 _1068_
rlabel metal2 21336 24024 21336 24024 0 _1069_
rlabel metal2 18648 24024 18648 24024 0 _1070_
rlabel metal2 19208 20216 19208 20216 0 _1071_
rlabel metal3 16828 24808 16828 24808 0 _1072_
rlabel metal2 5992 25760 5992 25760 0 _1073_
rlabel metal3 29568 30072 29568 30072 0 _1074_
rlabel metal2 29512 25592 29512 25592 0 _1075_
rlabel metal2 13720 8792 13720 8792 0 _1076_
rlabel metal2 10696 26096 10696 26096 0 _1077_
rlabel metal2 8120 25032 8120 25032 0 _1078_
rlabel metal2 18536 21336 18536 21336 0 _1079_
rlabel metal2 18312 20496 18312 20496 0 _1080_
rlabel metal2 23016 22624 23016 22624 0 _1081_
rlabel metal3 22960 11704 22960 11704 0 _1082_
rlabel metal3 16884 20552 16884 20552 0 _1083_
rlabel metal3 3304 20664 3304 20664 0 _1084_
rlabel metal2 17416 20888 17416 20888 0 _1085_
rlabel metal2 17640 20384 17640 20384 0 _1086_
rlabel metal2 6552 20048 6552 20048 0 _1087_
rlabel metal2 19992 23800 19992 23800 0 _1088_
rlabel metal2 19656 23408 19656 23408 0 _1089_
rlabel metal2 17752 23576 17752 23576 0 _1090_
rlabel metal2 18312 23576 18312 23576 0 _1091_
rlabel metal2 23128 23296 23128 23296 0 _1092_
rlabel metal2 23744 20552 23744 20552 0 _1093_
rlabel metal3 14560 14392 14560 14392 0 _1094_
rlabel metal2 12152 24640 12152 24640 0 _1095_
rlabel metal2 13608 26292 13608 26292 0 _1096_
rlabel metal2 11200 24136 11200 24136 0 _1097_
rlabel metal3 25648 24808 25648 24808 0 _1098_
rlabel metal2 24920 22008 24920 22008 0 _1099_
rlabel metal2 13496 14000 13496 14000 0 _1100_
rlabel metal2 13552 22568 13552 22568 0 _1101_
rlabel metal2 14168 22176 14168 22176 0 _1102_
rlabel metal3 11592 21672 11592 21672 0 _1103_
rlabel metal2 15512 42392 15512 42392 0 _1104_
rlabel metal2 18648 45024 18648 45024 0 _1105_
rlabel metal2 11592 29568 11592 29568 0 _1106_
rlabel metal2 10136 27048 10136 27048 0 _1107_
rlabel metal2 10584 29120 10584 29120 0 _1108_
rlabel metal2 8232 19208 8232 19208 0 _1109_
rlabel metal2 19880 22736 19880 22736 0 _1110_
rlabel metal3 21392 21560 21392 21560 0 _1111_
rlabel metal2 24584 21672 24584 21672 0 _1112_
rlabel metal3 21672 20104 21672 20104 0 _1113_
rlabel metal2 18872 19992 18872 19992 0 _1114_
rlabel metal2 22680 19936 22680 19936 0 _1115_
rlabel metal2 14392 7644 14392 7644 0 _1116_
rlabel metal2 14840 7392 14840 7392 0 _1117_
rlabel metal2 13832 6216 13832 6216 0 _1118_
rlabel metal2 12600 7840 12600 7840 0 _1119_
rlabel metal2 11480 6552 11480 6552 0 _1120_
rlabel metal2 19880 8232 19880 8232 0 _1121_
rlabel metal2 18312 6720 18312 6720 0 _1122_
rlabel metal3 17080 5880 17080 5880 0 _1123_
rlabel metal3 17192 7448 17192 7448 0 _1124_
rlabel metal2 7672 22736 7672 22736 0 _1125_
rlabel metal2 2744 22848 2744 22848 0 _1126_
rlabel metal3 5600 23352 5600 23352 0 _1127_
rlabel metal2 48216 46928 48216 46928 0 _1128_
rlabel metal2 50624 52136 50624 52136 0 _1129_
rlabel metal2 24920 25760 24920 25760 0 _1130_
rlabel metal2 22008 15512 22008 15512 0 _1131_
rlabel metal3 16744 15624 16744 15624 0 _1132_
rlabel metal2 14840 12936 14840 12936 0 _1133_
rlabel metal2 14392 9912 14392 9912 0 _1134_
rlabel metal2 10696 8316 10696 8316 0 _1135_
rlabel metal2 6888 12264 6888 12264 0 _1136_
rlabel metal2 8232 11928 8232 11928 0 _1137_
rlabel metal2 6888 10584 6888 10584 0 _1138_
rlabel metal2 9576 17416 9576 17416 0 _1139_
rlabel metal2 6664 9744 6664 9744 0 _1140_
rlabel metal2 25256 24528 25256 24528 0 _1141_
rlabel metal2 7336 14420 7336 14420 0 _1142_
rlabel metal2 2744 16744 2744 16744 0 _1143_
rlabel metal2 6216 14168 6216 14168 0 _1144_
rlabel metal2 6664 18480 6664 18480 0 _1145_
rlabel metal3 4704 17864 4704 17864 0 _1146_
rlabel metal2 2856 18760 2856 18760 0 _1147_
rlabel metal3 16184 14504 16184 14504 0 _1148_
rlabel metal2 6440 12936 6440 12936 0 _1149_
rlabel metal3 4536 13160 4536 13160 0 _1150_
rlabel metal3 4592 12376 4592 12376 0 _1151_
rlabel metal2 20608 21000 20608 21000 0 _1152_
rlabel metal2 21280 17976 21280 17976 0 _1153_
rlabel metal3 19656 10808 19656 10808 0 _1154_
rlabel metal2 18424 9912 18424 9912 0 _1155_
rlabel metal3 20048 9800 20048 9800 0 _1156_
rlabel metal2 21448 43512 21448 43512 0 _1157_
rlabel metal3 18088 40264 18088 40264 0 _1158_
rlabel metal2 21448 40712 21448 40712 0 _1159_
rlabel metal2 18760 40488 18760 40488 0 _1160_
rlabel metal3 22736 33096 22736 33096 0 _1161_
rlabel metal3 25536 31640 25536 31640 0 _1162_
rlabel metal3 18760 35112 18760 35112 0 _1163_
rlabel metal3 23128 34104 23128 34104 0 _1164_
rlabel metal2 26096 31864 26096 31864 0 _1165_
rlabel metal2 52696 35000 52696 35000 0 _1166_
rlabel metal2 16520 31640 16520 31640 0 _1167_
rlabel metal2 17752 31472 17752 31472 0 _1168_
rlabel metal2 22736 30408 22736 30408 0 _1169_
rlabel metal3 18872 31864 18872 31864 0 _1170_
rlabel metal3 19600 31640 19600 31640 0 _1171_
rlabel metal3 15624 31808 15624 31808 0 _1172_
rlabel metal2 24696 34216 24696 34216 0 _1173_
rlabel metal2 17640 32704 17640 32704 0 _1174_
rlabel metal2 44968 47040 44968 47040 0 _1175_
rlabel metal2 45192 47936 45192 47936 0 _1176_
rlabel metal2 45864 46032 45864 46032 0 _1177_
rlabel via2 48552 47544 48552 47544 0 _1178_
rlabel metal2 46088 47880 46088 47880 0 _1179_
rlabel metal3 48328 48216 48328 48216 0 _1180_
rlabel metal2 46424 47880 46424 47880 0 _1181_
rlabel metal2 46088 46872 46088 46872 0 _1182_
rlabel metal3 47768 46536 47768 46536 0 _1183_
rlabel metal2 47320 47712 47320 47712 0 _1184_
rlabel metal3 49112 47432 49112 47432 0 _1185_
rlabel metal2 49952 46648 49952 46648 0 _1186_
rlabel metal2 51352 47824 51352 47824 0 _1187_
rlabel metal2 51912 52192 51912 52192 0 _1188_
rlabel metal2 50904 51128 50904 51128 0 _1189_
rlabel metal2 49896 51968 49896 51968 0 _1190_
rlabel metal2 49952 50792 49952 50792 0 _1191_
rlabel metal2 49896 51184 49896 51184 0 _1192_
rlabel metal2 49896 52584 49896 52584 0 _1193_
rlabel metal2 49392 52808 49392 52808 0 _1194_
rlabel metal2 50232 50624 50232 50624 0 _1195_
rlabel metal2 51016 51408 51016 51408 0 _1196_
rlabel metal2 51128 51016 51128 51016 0 _1197_
rlabel metal3 32144 35784 32144 35784 0 _1198_
rlabel metal2 40824 44688 40824 44688 0 _1199_
rlabel metal2 33712 32648 33712 32648 0 _1200_
rlabel metal3 35840 33208 35840 33208 0 _1201_
rlabel metal2 37184 34664 37184 34664 0 _1202_
rlabel metal2 36904 32984 36904 32984 0 _1203_
rlabel metal3 38808 34048 38808 34048 0 _1204_
rlabel metal2 38024 38780 38024 38780 0 _1205_
rlabel metal2 37016 37184 37016 37184 0 _1206_
rlabel metal2 39312 35672 39312 35672 0 _1207_
rlabel metal2 37128 37408 37128 37408 0 _1208_
rlabel metal2 36456 37520 36456 37520 0 _1209_
rlabel metal2 37352 38724 37352 38724 0 _1210_
rlabel metal2 38136 39144 38136 39144 0 _1211_
rlabel metal2 38528 38920 38528 38920 0 _1212_
rlabel metal3 38472 38808 38472 38808 0 _1213_
rlabel metal2 38584 37576 38584 37576 0 _1214_
rlabel metal2 39032 37240 39032 37240 0 _1215_
rlabel metal2 39872 46648 39872 46648 0 _1216_
rlabel metal3 37856 37352 37856 37352 0 _1217_
rlabel metal3 37744 38024 37744 38024 0 _1218_
rlabel metal2 39816 37408 39816 37408 0 _1219_
rlabel metal2 43288 41440 43288 41440 0 _1220_
rlabel metal3 40208 45864 40208 45864 0 _1221_
rlabel metal2 40320 45976 40320 45976 0 _1222_
rlabel metal3 41944 45192 41944 45192 0 _1223_
rlabel metal2 39872 43736 39872 43736 0 _1224_
rlabel metal2 41496 43456 41496 43456 0 _1225_
rlabel metal2 40824 43400 40824 43400 0 _1226_
rlabel metal2 41720 44408 41720 44408 0 _1227_
rlabel metal3 42056 45080 42056 45080 0 _1228_
rlabel metal2 43624 40768 43624 40768 0 _1229_
rlabel metal2 45752 37408 45752 37408 0 _1230_
rlabel metal2 41608 31752 41608 31752 0 _1231_
rlabel metal2 46648 42728 46648 42728 0 _1232_
rlabel metal2 39704 41384 39704 41384 0 _1233_
rlabel metal3 42112 40936 42112 40936 0 _1234_
rlabel metal2 43848 40768 43848 40768 0 _1235_
rlabel metal2 39144 43904 39144 43904 0 _1236_
rlabel metal2 39592 41440 39592 41440 0 _1237_
rlabel metal3 40712 39928 40712 39928 0 _1238_
rlabel metal2 40040 31416 40040 31416 0 _1239_
rlabel metal2 49504 24472 49504 24472 0 _1240_
rlabel metal2 44296 28896 44296 28896 0 _1241_
rlabel metal2 50568 27104 50568 27104 0 _1242_
rlabel metal3 49728 22232 49728 22232 0 _1243_
rlabel metal2 48776 21896 48776 21896 0 _1244_
rlabel metal2 49896 22736 49896 22736 0 _1245_
rlabel metal3 52360 31192 52360 31192 0 _1246_
rlabel metal2 52136 31360 52136 31360 0 _1247_
rlabel metal2 45640 40376 45640 40376 0 _1248_
rlabel metal2 49000 34496 49000 34496 0 _1249_
rlabel metal2 49896 39648 49896 39648 0 _1250_
rlabel metal2 50456 34384 50456 34384 0 _1251_
rlabel metal2 52024 31892 52024 31892 0 _1252_
rlabel metal2 49224 33432 49224 33432 0 _1253_
rlabel metal2 53592 33264 53592 33264 0 _1254_
rlabel metal2 53368 35392 53368 35392 0 _1255_
rlabel metal2 47992 32256 47992 32256 0 _1256_
rlabel metal2 48328 30408 48328 30408 0 _1257_
rlabel metal2 52080 28392 52080 28392 0 _1258_
rlabel metal3 53704 27832 53704 27832 0 _1259_
rlabel metal2 46760 27216 46760 27216 0 _1260_
rlabel metal2 46592 25704 46592 25704 0 _1261_
rlabel metal2 47208 29288 47208 29288 0 _1262_
rlabel metal2 46928 30744 46928 30744 0 _1263_
rlabel metal2 47096 33488 47096 33488 0 _1264_
rlabel metal2 47208 33432 47208 33432 0 _1265_
rlabel metal2 47208 32816 47208 32816 0 _1266_
rlabel metal2 50456 27944 50456 27944 0 _1267_
rlabel metal2 47544 32648 47544 32648 0 _1268_
rlabel metal2 46760 32984 46760 32984 0 _1269_
rlabel metal2 46984 32032 46984 32032 0 _1270_
rlabel metal2 37856 31976 37856 31976 0 _1271_
rlabel metal3 37016 30184 37016 30184 0 _1272_
rlabel metal2 41720 23744 41720 23744 0 _1273_
rlabel metal2 39592 26488 39592 26488 0 _1274_
rlabel metal2 38472 29064 38472 29064 0 _1275_
rlabel metal2 46536 30688 46536 30688 0 _1276_
rlabel metal2 49336 32704 49336 32704 0 _1277_
rlabel metal2 48776 23128 48776 23128 0 _1278_
rlabel metal3 42280 39704 42280 39704 0 _1279_
rlabel metal2 42392 44240 42392 44240 0 _1280_
rlabel metal3 38696 43512 38696 43512 0 _1281_
rlabel metal2 38808 43120 38808 43120 0 _1282_
rlabel metal2 41832 42448 41832 42448 0 _1283_
rlabel metal2 42224 40376 42224 40376 0 _1284_
rlabel metal2 43960 38752 43960 38752 0 _1285_
rlabel metal2 45136 37240 45136 37240 0 _1286_
rlabel metal2 12488 13216 12488 13216 0 clknet_0_wb_clk_i
rlabel metal3 5320 13552 5320 13552 0 clknet_4_0_0_wb_clk_i
rlabel metal3 54096 26936 54096 26936 0 clknet_4_10_0_wb_clk_i
rlabel metal3 55160 30968 55160 30968 0 clknet_4_11_0_wb_clk_i
rlabel metal2 33992 49336 33992 49336 0 clknet_4_12_0_wb_clk_i
rlabel metal2 23912 54432 23912 54432 0 clknet_4_13_0_wb_clk_i
rlabel metal2 48272 40936 48272 40936 0 clknet_4_14_0_wb_clk_i
rlabel metal2 52696 50960 52696 50960 0 clknet_4_15_0_wb_clk_i
rlabel metal2 1848 21952 1848 21952 0 clknet_4_1_0_wb_clk_i
rlabel metal2 15736 11424 15736 11424 0 clknet_4_2_0_wb_clk_i
rlabel metal2 17528 18816 17528 18816 0 clknet_4_3_0_wb_clk_i
rlabel metal2 1848 38416 1848 38416 0 clknet_4_4_0_wb_clk_i
rlabel metal2 1848 54488 1848 54488 0 clknet_4_5_0_wb_clk_i
rlabel metal2 15736 26684 15736 26684 0 clknet_4_6_0_wb_clk_i
rlabel metal2 21000 48720 21000 48720 0 clknet_4_7_0_wb_clk_i
rlabel metal2 39424 12376 39424 12376 0 clknet_4_8_0_wb_clk_i
rlabel metal2 32648 24024 32648 24024 0 clknet_4_9_0_wb_clk_i
rlabel metal2 18984 56392 18984 56392 0 io_in[10]
rlabel metal2 20104 56168 20104 56168 0 io_in[11]
rlabel metal2 39200 55272 39200 55272 0 io_in[26]
rlabel metal2 14840 55720 14840 55720 0 io_in[8]
rlabel metal2 17192 56168 17192 56168 0 io_in[9]
rlabel metal3 21896 53704 21896 53704 0 io_out[12]
rlabel metal2 22120 56392 22120 56392 0 io_out[13]
rlabel metal2 23688 56392 23688 56392 0 io_out[14]
rlabel metal2 25592 57610 25592 57610 0 io_out[15]
rlabel metal2 26992 56280 26992 56280 0 io_out[16]
rlabel metal3 28784 54712 28784 54712 0 io_out[17]
rlabel metal2 30744 56112 30744 56112 0 io_out[18]
rlabel metal2 32648 56112 32648 56112 0 io_out[19]
rlabel metal2 34216 56504 34216 56504 0 io_out[20]
rlabel metal2 36456 56448 36456 56448 0 io_out[21]
rlabel metal2 38024 56504 38024 56504 0 io_out[22]
rlabel metal3 36904 55384 36904 55384 0 io_out[23]
rlabel metal2 40488 56336 40488 56336 0 io_out[24]
rlabel metal2 42056 56392 42056 56392 0 io_out[25]
rlabel metal2 18648 55328 18648 55328 0 net1
rlabel metal2 25088 52248 25088 52248 0 net10
rlabel metal2 44856 44520 44856 44520 0 net11
rlabel metal2 28616 54936 28616 54936 0 net12
rlabel metal2 30352 52808 30352 52808 0 net13
rlabel metal2 32088 55720 32088 55720 0 net14
rlabel metal2 33320 53256 33320 53256 0 net15
rlabel metal2 33768 54376 33768 54376 0 net16
rlabel metal2 35336 55440 35336 55440 0 net17
rlabel metal2 37800 54824 37800 54824 0 net18
rlabel metal2 39704 55720 39704 55720 0 net19
rlabel metal3 19208 55384 19208 55384 0 net2
rlabel metal2 42728 55216 42728 55216 0 net20
rlabel metal2 21840 55160 21840 55160 0 net21
rlabel metal2 22176 55160 22176 55160 0 net22
rlabel metal2 24696 57778 24696 57778 0 net23
rlabel metal2 26152 54712 26152 54712 0 net24
rlabel metal2 28392 56448 28392 56448 0 net25
rlabel metal2 28840 56280 28840 56280 0 net26
rlabel metal2 29512 56448 29512 56448 0 net27
rlabel metal2 31472 56280 31472 56280 0 net28
rlabel metal2 32928 54712 32928 54712 0 net29
rlabel metal3 40824 53704 40824 53704 0 net3
rlabel metal3 34720 56280 34720 56280 0 net30
rlabel metal2 36288 55160 36288 55160 0 net31
rlabel metal2 36792 57778 36792 57778 0 net32
rlabel metal2 38584 56224 38584 56224 0 net33
rlabel metal2 39592 54712 39592 54712 0 net34
rlabel metal2 4984 56336 4984 56336 0 net35
rlabel metal2 6888 56280 6888 56280 0 net36
rlabel metal2 8176 56280 8176 56280 0 net37
rlabel metal2 9576 56280 9576 56280 0 net38
rlabel metal2 10920 56280 10920 56280 0 net39
rlabel metal2 16296 55328 16296 55328 0 net4
rlabel metal2 12264 56280 12264 56280 0 net40
rlabel metal2 13608 56280 13608 56280 0 net41
rlabel metal2 14784 56280 14784 56280 0 net42
rlabel metal2 15176 56672 15176 56672 0 net43
rlabel metal2 15624 56672 15624 56672 0 net44
rlabel metal2 18312 56336 18312 56336 0 net45
rlabel metal2 20440 56168 20440 56168 0 net46
rlabel metal2 40936 55832 40936 55832 0 net47
rlabel metal3 42672 56280 42672 56280 0 net48
rlabel metal2 43400 55664 43400 55664 0 net49
rlabel metal2 18424 55160 18424 55160 0 net5
rlabel metal2 44968 56672 44968 56672 0 net50
rlabel metal2 45864 56280 45864 56280 0 net51
rlabel metal2 47432 57008 47432 57008 0 net52
rlabel metal2 48552 56280 48552 56280 0 net53
rlabel metal2 49896 56280 49896 56280 0 net54
rlabel metal2 51240 56280 51240 56280 0 net55
rlabel metal2 52584 56280 52584 56280 0 net56
rlabel metal2 53928 56280 53928 56280 0 net57
rlabel metal2 55160 57778 55160 57778 0 net58
rlabel metal2 6216 56728 6216 56728 0 net59
rlabel metal2 8456 55804 8456 55804 0 net6
rlabel metal2 7336 55944 7336 55944 0 net60
rlabel metal2 8624 55944 8624 55944 0 net61
rlabel metal2 10024 55944 10024 55944 0 net62
rlabel metal2 11368 55944 11368 55944 0 net63
rlabel metal2 13160 56280 13160 56280 0 net64
rlabel metal2 14056 55944 14056 55944 0 net65
rlabel metal2 15400 55496 15400 55496 0 net66
rlabel metal2 16184 56448 16184 56448 0 net67
rlabel metal3 18592 55496 18592 55496 0 net68
rlabel metal2 19376 55944 19376 55944 0 net69
rlabel metal2 25256 51464 25256 51464 0 net7
rlabel metal2 20720 55944 20720 55944 0 net70
rlabel metal2 42952 56504 42952 56504 0 net71
rlabel metal2 44072 56448 44072 56448 0 net72
rlabel metal3 44016 55944 44016 55944 0 net73
rlabel metal3 45136 55832 45136 55832 0 net74
rlabel metal2 46312 55944 46312 55944 0 net75
rlabel metal2 47712 55944 47712 55944 0 net76
rlabel metal2 49000 55944 49000 55944 0 net77
rlabel metal2 50232 57610 50232 57610 0 net78
rlabel metal2 51688 55944 51688 55944 0 net79
rlabel metal2 21000 53984 21000 53984 0 net8
rlabel metal2 53032 55944 53032 55944 0 net80
rlabel metal2 55048 56280 55048 56280 0 net81
rlabel metal2 55944 56728 55944 56728 0 net82
rlabel metal2 22456 54208 22456 54208 0 net9
rlabel metal2 11256 44576 11256 44576 0 simon1.millis_counter\[0\]
rlabel metal2 12040 45864 12040 45864 0 simon1.millis_counter\[1\]
rlabel metal2 12152 48664 12152 48664 0 simon1.millis_counter\[2\]
rlabel metal2 15176 48664 15176 48664 0 simon1.millis_counter\[3\]
rlabel metal3 13664 50456 13664 50456 0 simon1.millis_counter\[4\]
rlabel metal2 11368 51408 11368 51408 0 simon1.millis_counter\[5\]
rlabel metal2 12824 52976 12824 52976 0 simon1.millis_counter\[6\]
rlabel metal2 14840 52192 14840 52192 0 simon1.millis_counter\[7\]
rlabel metal2 18592 48328 18592 48328 0 simon1.millis_counter\[8\]
rlabel metal2 18368 48440 18368 48440 0 simon1.millis_counter\[9\]
rlabel metal2 29176 32144 29176 32144 0 simon1.next_random\[0\]
rlabel metal2 30744 30072 30744 30072 0 simon1.next_random\[1\]
rlabel metal2 32536 33936 32536 33936 0 simon1.play1.freq\[0\]
rlabel metal2 29288 34720 29288 34720 0 simon1.play1.freq\[1\]
rlabel metal2 38696 37464 38696 37464 0 simon1.play1.freq\[2\]
rlabel metal2 36064 36456 36064 36456 0 simon1.play1.freq\[3\]
rlabel metal2 38360 45472 38360 45472 0 simon1.play1.freq\[4\]
rlabel metal2 38024 43848 38024 43848 0 simon1.play1.freq\[5\]
rlabel metal2 39928 39648 39928 39648 0 simon1.play1.freq\[6\]
rlabel metal2 39256 40656 39256 40656 0 simon1.play1.freq\[7\]
rlabel metal2 46872 42672 46872 42672 0 simon1.play1.freq\[8\]
rlabel metal2 39872 41944 39872 41944 0 simon1.play1.freq\[9\]
rlabel metal3 42056 33992 42056 33992 0 simon1.play1.tick_counter\[0\]
rlabel metal2 52920 37352 52920 37352 0 simon1.play1.tick_counter\[10\]
rlabel metal2 51800 38136 51800 38136 0 simon1.play1.tick_counter\[11\]
rlabel metal3 53256 32648 53256 32648 0 simon1.play1.tick_counter\[12\]
rlabel metal2 54264 32928 54264 32928 0 simon1.play1.tick_counter\[13\]
rlabel metal2 54656 30296 54656 30296 0 simon1.play1.tick_counter\[14\]
rlabel metal2 53480 31024 53480 31024 0 simon1.play1.tick_counter\[15\]
rlabel metal2 54096 27048 54096 27048 0 simon1.play1.tick_counter\[16\]
rlabel metal2 54040 25648 54040 25648 0 simon1.play1.tick_counter\[17\]
rlabel metal2 51464 29344 51464 29344 0 simon1.play1.tick_counter\[18\]
rlabel metal2 53368 25424 53368 25424 0 simon1.play1.tick_counter\[19\]
rlabel metal2 39928 33768 39928 33768 0 simon1.play1.tick_counter\[1\]
rlabel metal2 44184 25424 44184 25424 0 simon1.play1.tick_counter\[20\]
rlabel metal2 43960 22680 43960 22680 0 simon1.play1.tick_counter\[21\]
rlabel metal2 45752 25424 45752 25424 0 simon1.play1.tick_counter\[22\]
rlabel metal3 43288 25480 43288 25480 0 simon1.play1.tick_counter\[23\]
rlabel metal2 41272 21224 41272 21224 0 simon1.play1.tick_counter\[24\]
rlabel metal2 39928 25816 39928 25816 0 simon1.play1.tick_counter\[25\]
rlabel metal2 38920 22120 38920 22120 0 simon1.play1.tick_counter\[26\]
rlabel metal2 37352 27496 37352 27496 0 simon1.play1.tick_counter\[27\]
rlabel metal2 32648 25984 32648 25984 0 simon1.play1.tick_counter\[28\]
rlabel metal2 35112 28168 35112 28168 0 simon1.play1.tick_counter\[29\]
rlabel metal2 38808 36792 38808 36792 0 simon1.play1.tick_counter\[2\]
rlabel metal2 35952 30184 35952 30184 0 simon1.play1.tick_counter\[30\]
rlabel metal2 39256 31248 39256 31248 0 simon1.play1.tick_counter\[31\]
rlabel metal2 42504 36624 42504 36624 0 simon1.play1.tick_counter\[3\]
rlabel metal2 43848 46312 43848 46312 0 simon1.play1.tick_counter\[4\]
rlabel metal3 45024 44072 45024 44072 0 simon1.play1.tick_counter\[5\]
rlabel metal2 42504 37520 42504 37520 0 simon1.play1.tick_counter\[6\]
rlabel metal2 44968 41272 44968 41272 0 simon1.play1.tick_counter\[7\]
rlabel metal2 49896 43624 49896 43624 0 simon1.play1.tick_counter\[8\]
rlabel metal2 51688 39088 51688 39088 0 simon1.play1.tick_counter\[9\]
rlabel metal2 47880 52472 47880 52472 0 simon1.score1.active_digit
rlabel metal3 45696 50232 45696 50232 0 simon1.score1.ena
rlabel metal2 44520 46872 44520 46872 0 simon1.score1.inc
rlabel metal2 44744 47320 44744 47320 0 simon1.score1.ones\[0\]
rlabel metal2 47712 47432 47712 47432 0 simon1.score1.ones\[1\]
rlabel metal3 47992 49224 47992 49224 0 simon1.score1.ones\[2\]
rlabel metal3 52024 44968 52024 44968 0 simon1.score1.ones\[3\]
rlabel metal2 49672 47992 49672 47992 0 simon1.score1.tens\[0\]
rlabel metal2 51744 51912 51744 51912 0 simon1.score1.tens\[1\]
rlabel via2 51464 52920 51464 52920 0 simon1.score1.tens\[2\]
rlabel metal2 50792 51016 50792 51016 0 simon1.score1.tens\[3\]
rlabel metal3 30520 37128 30520 37128 0 simon1.score_rst
rlabel metal2 11928 20048 11928 20048 0 simon1.seq\[0\]\[0\]
rlabel metal2 11816 21280 11816 21280 0 simon1.seq\[0\]\[1\]
rlabel metal2 15512 23184 15512 23184 0 simon1.seq\[10\]\[0\]
rlabel metal3 13384 21560 13384 21560 0 simon1.seq\[10\]\[1\]
rlabel metal2 15288 25760 15288 25760 0 simon1.seq\[11\]\[0\]
rlabel metal2 12264 23520 12264 23520 0 simon1.seq\[11\]\[1\]
rlabel metal2 4648 21392 4648 21392 0 simon1.seq\[12\]\[0\]
rlabel metal3 8624 19880 8624 19880 0 simon1.seq\[12\]\[1\]
rlabel metal2 7112 24304 7112 24304 0 simon1.seq\[13\]\[0\]
rlabel metal3 9408 25592 9408 25592 0 simon1.seq\[13\]\[1\]
rlabel metal3 17304 5992 17304 5992 0 simon1.seq\[14\]\[0\]
rlabel metal2 14728 7840 14728 7840 0 simon1.seq\[14\]\[1\]
rlabel metal2 15288 6216 15288 6216 0 simon1.seq\[15\]\[0\]
rlabel metal3 13664 7560 13664 7560 0 simon1.seq\[15\]\[1\]
rlabel metal2 20440 19544 20440 19544 0 simon1.seq\[16\]\[0\]
rlabel metal2 24248 19040 24248 19040 0 simon1.seq\[16\]\[1\]
rlabel via2 26488 22344 26488 22344 0 simon1.seq\[17\]\[0\]
rlabel metal2 29400 24024 29400 24024 0 simon1.seq\[17\]\[1\]
rlabel metal3 32984 21336 32984 21336 0 simon1.seq\[18\]\[0\]
rlabel metal2 35448 20272 35448 20272 0 simon1.seq\[18\]\[1\]
rlabel metal2 35112 16296 35112 16296 0 simon1.seq\[19\]\[0\]
rlabel metal3 34832 15176 34832 15176 0 simon1.seq\[19\]\[1\]
rlabel metal2 11144 15736 11144 15736 0 simon1.seq\[1\]\[0\]
rlabel metal3 11424 14616 11424 14616 0 simon1.seq\[1\]\[1\]
rlabel metal3 19488 12152 19488 12152 0 simon1.seq\[20\]\[0\]
rlabel metal2 19432 12880 19432 12880 0 simon1.seq\[20\]\[1\]
rlabel metal2 20104 10136 20104 10136 0 simon1.seq\[21\]\[0\]
rlabel via2 22904 11256 22904 11256 0 simon1.seq\[21\]\[1\]
rlabel metal2 22568 6104 22568 6104 0 simon1.seq\[22\]\[0\]
rlabel metal2 24416 5992 24416 5992 0 simon1.seq\[22\]\[1\]
rlabel metal2 23128 8512 23128 8512 0 simon1.seq\[23\]\[0\]
rlabel metal3 22904 8288 22904 8288 0 simon1.seq\[23\]\[1\]
rlabel metal2 28504 19208 28504 19208 0 simon1.seq\[24\]\[0\]
rlabel metal2 30184 18536 30184 18536 0 simon1.seq\[24\]\[1\]
rlabel via2 27720 10472 27720 10472 0 simon1.seq\[25\]\[0\]
rlabel metal3 28280 8344 28280 8344 0 simon1.seq\[25\]\[1\]
rlabel metal3 31360 16184 31360 16184 0 simon1.seq\[26\]\[0\]
rlabel metal2 29624 13552 29624 13552 0 simon1.seq\[26\]\[1\]
rlabel metal2 21224 16632 21224 16632 0 simon1.seq\[27\]\[0\]
rlabel metal2 24248 14560 24248 14560 0 simon1.seq\[27\]\[1\]
rlabel metal3 29568 10696 29568 10696 0 simon1.seq\[28\]\[0\]
rlabel metal2 29288 10080 29288 10080 0 simon1.seq\[28\]\[1\]
rlabel metal2 28280 5488 28280 5488 0 simon1.seq\[29\]\[0\]
rlabel metal2 27944 5096 27944 5096 0 simon1.seq\[29\]\[1\]
rlabel metal2 11704 13104 11704 13104 0 simon1.seq\[2\]\[0\]
rlabel metal2 13944 12376 13944 12376 0 simon1.seq\[2\]\[1\]
rlabel metal2 34328 12544 34328 12544 0 simon1.seq\[30\]\[0\]
rlabel metal2 36344 11648 36344 11648 0 simon1.seq\[30\]\[1\]
rlabel metal3 34104 19320 34104 19320 0 simon1.seq\[31\]\[0\]
rlabel metal2 35336 18256 35336 18256 0 simon1.seq\[31\]\[1\]
rlabel metal2 4984 12992 4984 12992 0 simon1.seq\[3\]\[0\]
rlabel metal2 5432 12376 5432 12376 0 simon1.seq\[3\]\[1\]
rlabel metal2 6048 17640 6048 17640 0 simon1.seq\[4\]\[0\]
rlabel metal3 7448 18424 7448 18424 0 simon1.seq\[4\]\[1\]
rlabel metal2 6160 16296 6160 16296 0 simon1.seq\[5\]\[0\]
rlabel metal2 6664 16856 6664 16856 0 simon1.seq\[5\]\[1\]
rlabel metal2 7448 11088 7448 11088 0 simon1.seq\[6\]\[0\]
rlabel metal2 7672 9352 7672 9352 0 simon1.seq\[6\]\[1\]
rlabel metal2 15064 10304 15064 10304 0 simon1.seq\[7\]\[0\]
rlabel metal2 12488 10360 12488 10360 0 simon1.seq\[7\]\[1\]
rlabel metal2 6104 22120 6104 22120 0 simon1.seq\[8\]\[0\]
rlabel metal2 6888 22736 6888 22736 0 simon1.seq\[8\]\[1\]
rlabel metal2 7448 27832 7448 27832 0 simon1.seq\[9\]\[0\]
rlabel via2 8568 28616 8568 28616 0 simon1.seq\[9\]\[1\]
rlabel metal2 25256 30632 25256 30632 0 simon1.seq_counter\[0\]
rlabel metal2 21560 32032 21560 32032 0 simon1.seq_counter\[1\]
rlabel metal2 21448 30520 21448 30520 0 simon1.seq_counter\[2\]
rlabel metal2 15288 32368 15288 32368 0 simon1.seq_counter\[3\]
rlabel metal2 16632 32536 16632 32536 0 simon1.seq_counter\[4\]
rlabel metal3 25536 24920 25536 24920 0 simon1.seq_length\[0\]
rlabel via2 26264 27832 26264 27832 0 simon1.seq_length\[1\]
rlabel metal2 21616 25480 21616 25480 0 simon1.seq_length\[2\]
rlabel metal2 19656 24584 19656 24584 0 simon1.seq_length\[3\]
rlabel metal2 19992 21168 19992 21168 0 simon1.seq_length\[4\]
rlabel metal3 22008 38472 22008 38472 0 simon1.state\[0\]
rlabel metal2 19040 41720 19040 41720 0 simon1.state\[1\]
rlabel metal2 21336 39648 21336 39648 0 simon1.state\[2\]
rlabel metal2 18200 37744 18200 37744 0 simon1.state\[3\]
rlabel metal2 12488 39928 12488 39928 0 simon1.state\[4\]
rlabel metal2 25648 36232 25648 36232 0 simon1.state\[5\]
rlabel metal2 19656 37184 19656 37184 0 simon1.state\[6\]
rlabel metal2 20216 46480 20216 46480 0 simon1.state\[7\]
rlabel metal2 4648 53872 4648 53872 0 simon1.tick_counter\[0\]
rlabel metal2 5320 39256 5320 39256 0 simon1.tick_counter\[10\]
rlabel via2 5880 41048 5880 41048 0 simon1.tick_counter\[11\]
rlabel metal2 4984 42672 4984 42672 0 simon1.tick_counter\[12\]
rlabel metal2 4648 43344 4648 43344 0 simon1.tick_counter\[13\]
rlabel metal2 2744 44688 2744 44688 0 simon1.tick_counter\[14\]
rlabel metal2 3192 46536 3192 46536 0 simon1.tick_counter\[15\]
rlabel metal2 4312 52528 4312 52528 0 simon1.tick_counter\[1\]
rlabel metal2 4648 50736 4648 50736 0 simon1.tick_counter\[2\]
rlabel metal2 7224 51800 7224 51800 0 simon1.tick_counter\[3\]
rlabel metal2 7560 51240 7560 51240 0 simon1.tick_counter\[4\]
rlabel metal2 3976 49000 3976 49000 0 simon1.tick_counter\[5\]
rlabel metal2 7112 47936 7112 47936 0 simon1.tick_counter\[6\]
rlabel metal3 7952 44408 7952 44408 0 simon1.tick_counter\[7\]
rlabel metal3 8120 38808 8120 38808 0 simon1.tick_counter\[8\]
rlabel metal2 5824 39144 5824 39144 0 simon1.tick_counter\[9\]
rlabel metal2 31696 49896 31696 49896 0 simon1.tone_sequence_counter\[0\]
rlabel metal3 30912 49672 30912 49672 0 simon1.tone_sequence_counter\[1\]
rlabel metal2 33208 47880 33208 47880 0 simon1.tone_sequence_counter\[2\]
rlabel metal2 24920 45080 24920 45080 0 simon1.user_input\[0\]
rlabel metal2 25368 44016 25368 44016 0 simon1.user_input\[1\]
rlabel metal2 4088 56546 4088 56546 0 wb_clk_i
rlabel metal2 4592 56280 4592 56280 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
