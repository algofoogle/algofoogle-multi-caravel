magic
tech gf180mcuD
magscale 1 10
timestamp 1702302759
<< metal1 >>
rect 27010 50318 27022 50370
rect 27074 50367 27086 50370
rect 27906 50367 27918 50370
rect 27074 50321 27918 50367
rect 27074 50318 27086 50321
rect 27906 50318 27918 50321
rect 27970 50318 27982 50370
rect 1344 50202 48720 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 48720 50202
rect 1344 50116 48720 50150
rect 27022 50034 27074 50046
rect 27022 49970 27074 49982
rect 29486 49922 29538 49934
rect 29486 49858 29538 49870
rect 32846 49922 32898 49934
rect 32846 49858 32898 49870
rect 29822 49810 29874 49822
rect 26786 49758 26798 49810
rect 26850 49758 26862 49810
rect 32610 49758 32622 49810
rect 32674 49758 32686 49810
rect 29822 49746 29874 49758
rect 21086 49698 21138 49710
rect 21086 49634 21138 49646
rect 21534 49698 21586 49710
rect 21534 49634 21586 49646
rect 28926 49698 28978 49710
rect 28926 49634 28978 49646
rect 1344 49418 48720 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 48720 49418
rect 1344 49332 48720 49366
rect 14466 48974 14478 49026
rect 14530 48974 14542 49026
rect 15026 48974 15038 49026
rect 15090 48974 15102 49026
rect 17602 48974 17614 49026
rect 17666 48974 17678 49026
rect 18274 48974 18286 49026
rect 18338 48974 18350 49026
rect 21410 48974 21422 49026
rect 21474 48974 21486 49026
rect 21858 48974 21870 49026
rect 21922 48974 21934 49026
rect 27906 48974 27918 49026
rect 27970 48974 27982 49026
rect 28690 48974 28702 49026
rect 28754 48974 28766 49026
rect 29250 48974 29262 49026
rect 29314 48974 29326 49026
rect 29698 48974 29710 49026
rect 29762 48974 29774 49026
rect 32610 48974 32622 49026
rect 32674 48974 32686 49026
rect 33282 48974 33294 49026
rect 33346 48974 33358 49026
rect 37090 48974 37102 49026
rect 37154 48974 37166 49026
rect 37538 48974 37550 49026
rect 37602 48974 37614 49026
rect 36206 48802 36258 48814
rect 40462 48802 40514 48814
rect 17378 48750 17390 48802
rect 17442 48750 17454 48802
rect 20738 48750 20750 48802
rect 20802 48750 20814 48802
rect 24322 48750 24334 48802
rect 24386 48750 24398 48802
rect 25554 48750 25566 48802
rect 25618 48750 25630 48802
rect 32162 48750 32174 48802
rect 32226 48750 32238 48802
rect 35746 48750 35758 48802
rect 35810 48750 35822 48802
rect 40002 48750 40014 48802
rect 40066 48750 40078 48802
rect 36206 48738 36258 48750
rect 40462 48738 40514 48750
rect 1344 48634 48720 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 48720 48634
rect 1344 48548 48720 48582
rect 16270 48466 16322 48478
rect 16270 48402 16322 48414
rect 17614 48466 17666 48478
rect 17614 48402 17666 48414
rect 18174 48466 18226 48478
rect 18174 48402 18226 48414
rect 27358 48466 27410 48478
rect 27358 48402 27410 48414
rect 29934 48466 29986 48478
rect 29934 48402 29986 48414
rect 33182 48466 33234 48478
rect 33182 48402 33234 48414
rect 37550 48466 37602 48478
rect 37550 48402 37602 48414
rect 22654 48354 22706 48366
rect 19842 48302 19854 48354
rect 19906 48302 19918 48354
rect 21522 48302 21534 48354
rect 21586 48302 21598 48354
rect 21970 48302 21982 48354
rect 22034 48302 22046 48354
rect 22654 48290 22706 48302
rect 24110 48354 24162 48366
rect 39902 48354 39954 48366
rect 28242 48302 28254 48354
rect 28306 48302 28318 48354
rect 30818 48302 30830 48354
rect 30882 48302 30894 48354
rect 33730 48302 33742 48354
rect 33794 48302 33806 48354
rect 34066 48302 34078 48354
rect 34130 48302 34142 48354
rect 38882 48302 38894 48354
rect 38946 48302 38958 48354
rect 24110 48290 24162 48302
rect 39902 48290 39954 48302
rect 16606 48242 16658 48254
rect 16606 48178 16658 48190
rect 18510 48242 18562 48254
rect 18510 48178 18562 48190
rect 18958 48242 19010 48254
rect 24446 48242 24498 48254
rect 30270 48242 30322 48254
rect 37998 48242 38050 48254
rect 39566 48242 39618 48254
rect 20066 48190 20078 48242
rect 20130 48190 20142 48242
rect 28466 48190 28478 48242
rect 28530 48190 28542 48242
rect 30706 48190 30718 48242
rect 30770 48190 30782 48242
rect 37314 48190 37326 48242
rect 37378 48190 37390 48242
rect 38770 48190 38782 48242
rect 38834 48190 38846 48242
rect 18958 48178 19010 48190
rect 24446 48178 24498 48190
rect 30270 48178 30322 48190
rect 37998 48178 38050 48190
rect 39566 48178 39618 48190
rect 32398 48130 32450 48142
rect 32398 48066 32450 48078
rect 40350 48130 40402 48142
rect 40350 48066 40402 48078
rect 19294 48018 19346 48030
rect 19294 47954 19346 47966
rect 20974 48018 21026 48030
rect 20974 47954 21026 47966
rect 21310 48018 21362 48030
rect 21310 47954 21362 47966
rect 27694 48018 27746 48030
rect 27694 47954 27746 47966
rect 33518 48018 33570 48030
rect 33518 47954 33570 47966
rect 38334 48018 38386 48030
rect 40114 47966 40126 48018
rect 40178 48015 40190 48018
rect 40338 48015 40350 48018
rect 40178 47969 40350 48015
rect 40178 47966 40190 47969
rect 40338 47966 40350 47969
rect 40402 47966 40414 48018
rect 38334 47954 38386 47966
rect 1344 47850 48720 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 48720 47850
rect 1344 47764 48720 47798
rect 17278 47682 17330 47694
rect 17278 47618 17330 47630
rect 38894 47682 38946 47694
rect 38894 47618 38946 47630
rect 17614 47458 17666 47470
rect 21310 47458 21362 47470
rect 38558 47458 38610 47470
rect 9986 47406 9998 47458
rect 10050 47406 10062 47458
rect 10546 47406 10558 47458
rect 10610 47406 10622 47458
rect 18386 47406 18398 47458
rect 18450 47406 18462 47458
rect 23202 47406 23214 47458
rect 23266 47406 23278 47458
rect 23986 47406 23998 47458
rect 24050 47406 24062 47458
rect 32610 47406 32622 47458
rect 32674 47406 32686 47458
rect 33058 47406 33070 47458
rect 33122 47406 33134 47458
rect 39218 47406 39230 47458
rect 39282 47406 39294 47458
rect 39890 47406 39902 47458
rect 39954 47406 39966 47458
rect 17614 47394 17666 47406
rect 21310 47394 21362 47406
rect 38558 47394 38610 47406
rect 21646 47346 21698 47358
rect 18162 47294 18174 47346
rect 18226 47294 18238 47346
rect 21646 47282 21698 47294
rect 31838 47346 31890 47358
rect 31838 47282 31890 47294
rect 32174 47346 32226 47358
rect 37986 47294 37998 47346
rect 38050 47294 38062 47346
rect 38210 47294 38222 47346
rect 38274 47294 38286 47346
rect 32174 47282 32226 47294
rect 13582 47234 13634 47246
rect 12898 47182 12910 47234
rect 12962 47182 12974 47234
rect 13582 47170 13634 47182
rect 22990 47234 23042 47246
rect 35982 47234 36034 47246
rect 26338 47182 26350 47234
rect 26402 47182 26414 47234
rect 35522 47182 35534 47234
rect 35586 47182 35598 47234
rect 42354 47182 42366 47234
rect 42418 47182 42430 47234
rect 22990 47170 23042 47182
rect 35982 47170 36034 47182
rect 1344 47066 48720 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 48720 47066
rect 1344 46980 48720 47014
rect 10894 46898 10946 46910
rect 10894 46834 10946 46846
rect 11678 46898 11730 46910
rect 11678 46834 11730 46846
rect 12910 46898 12962 46910
rect 12910 46834 12962 46846
rect 25342 46898 25394 46910
rect 25342 46834 25394 46846
rect 31278 46898 31330 46910
rect 31278 46834 31330 46846
rect 39454 46898 39506 46910
rect 39454 46834 39506 46846
rect 40238 46898 40290 46910
rect 40238 46834 40290 46846
rect 9550 46786 9602 46798
rect 9550 46722 9602 46734
rect 17390 46786 17442 46798
rect 27806 46786 27858 46798
rect 26338 46734 26350 46786
rect 26402 46734 26414 46786
rect 31938 46734 31950 46786
rect 32002 46734 32014 46786
rect 32386 46734 32398 46786
rect 32450 46734 32462 46786
rect 35186 46734 35198 46786
rect 35250 46734 35262 46786
rect 35746 46734 35758 46786
rect 35810 46734 35822 46786
rect 38658 46734 38670 46786
rect 38722 46734 38734 46786
rect 17390 46722 17442 46734
rect 27806 46722 27858 46734
rect 9886 46674 9938 46686
rect 9886 46610 9938 46622
rect 11230 46674 11282 46686
rect 27470 46674 27522 46686
rect 13122 46622 13134 46674
rect 13186 46622 13198 46674
rect 13906 46622 13918 46674
rect 13970 46622 13982 46674
rect 17602 46622 17614 46674
rect 17666 46622 17678 46674
rect 26114 46622 26126 46674
rect 26178 46622 26190 46674
rect 11230 46610 11282 46622
rect 27470 46610 27522 46622
rect 30606 46674 30658 46686
rect 38882 46622 38894 46674
rect 38946 46622 38958 46674
rect 30606 46610 30658 46622
rect 34974 46562 35026 46574
rect 16258 46510 16270 46562
rect 16322 46510 16334 46562
rect 30146 46510 30158 46562
rect 30210 46510 30222 46562
rect 34974 46498 35026 46510
rect 25678 46450 25730 46462
rect 25678 46386 25730 46398
rect 31614 46450 31666 46462
rect 31614 46386 31666 46398
rect 34638 46450 34690 46462
rect 34638 46386 34690 46398
rect 37774 46450 37826 46462
rect 37774 46386 37826 46398
rect 38110 46450 38162 46462
rect 38110 46386 38162 46398
rect 1344 46282 48720 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48720 46282
rect 1344 46196 48720 46230
rect 11678 46114 11730 46126
rect 11678 46050 11730 46062
rect 27358 46114 27410 46126
rect 27358 46050 27410 46062
rect 27694 46114 27746 46126
rect 27694 46050 27746 46062
rect 41134 46114 41186 46126
rect 41134 46050 41186 46062
rect 19630 46002 19682 46014
rect 19630 45938 19682 45950
rect 26910 46002 26962 46014
rect 40002 45950 40014 46002
rect 40066 45950 40078 46002
rect 26910 45938 26962 45950
rect 12014 45890 12066 45902
rect 14030 45890 14082 45902
rect 8306 45838 8318 45890
rect 8370 45838 8382 45890
rect 8866 45838 8878 45890
rect 8930 45838 8942 45890
rect 12674 45838 12686 45890
rect 12738 45838 12750 45890
rect 16258 45838 16270 45890
rect 16322 45838 16334 45890
rect 16706 45838 16718 45890
rect 16770 45838 16782 45890
rect 20514 45838 20526 45890
rect 20578 45838 20590 45890
rect 21186 45838 21198 45890
rect 21250 45838 21262 45890
rect 21858 45838 21870 45890
rect 21922 45838 21934 45890
rect 28354 45838 28366 45890
rect 28418 45838 28430 45890
rect 37090 45838 37102 45890
rect 37154 45838 37166 45890
rect 37650 45838 37662 45890
rect 37714 45838 37726 45890
rect 43026 45838 43038 45890
rect 43090 45838 43102 45890
rect 12014 45826 12066 45838
rect 14030 45826 14082 45838
rect 20750 45778 20802 45790
rect 12786 45726 12798 45778
rect 12850 45726 12862 45778
rect 14354 45726 14366 45778
rect 14418 45726 14430 45778
rect 14802 45726 14814 45778
rect 14866 45726 14878 45778
rect 20750 45714 20802 45726
rect 25006 45778 25058 45790
rect 28466 45726 28478 45778
rect 28530 45726 28542 45778
rect 41346 45726 41358 45778
rect 41410 45726 41422 45778
rect 41682 45726 41694 45778
rect 41746 45726 41758 45778
rect 25006 45714 25058 45726
rect 13694 45666 13746 45678
rect 24670 45666 24722 45678
rect 11218 45614 11230 45666
rect 11282 45614 11294 45666
rect 19170 45614 19182 45666
rect 19234 45614 19246 45666
rect 24322 45614 24334 45666
rect 24386 45614 24398 45666
rect 13694 45602 13746 45614
rect 24670 45602 24722 45614
rect 40798 45666 40850 45678
rect 40798 45602 40850 45614
rect 42814 45666 42866 45678
rect 42814 45602 42866 45614
rect 1344 45498 48720 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48720 45498
rect 1344 45412 48720 45446
rect 10222 45330 10274 45342
rect 10222 45266 10274 45278
rect 13918 45330 13970 45342
rect 13918 45266 13970 45278
rect 17502 45330 17554 45342
rect 17502 45266 17554 45278
rect 20974 45330 21026 45342
rect 20974 45266 21026 45278
rect 25342 45330 25394 45342
rect 31502 45330 31554 45342
rect 37774 45330 37826 45342
rect 29922 45278 29934 45330
rect 29986 45278 29998 45330
rect 37426 45278 37438 45330
rect 37490 45278 37502 45330
rect 25342 45266 25394 45278
rect 31502 45266 31554 45278
rect 37774 45266 37826 45278
rect 40910 45218 40962 45230
rect 11330 45166 11342 45218
rect 11394 45166 11406 45218
rect 18498 45166 18510 45218
rect 18562 45166 18574 45218
rect 26226 45166 26238 45218
rect 26290 45166 26302 45218
rect 40910 45154 40962 45166
rect 30270 45106 30322 45118
rect 11106 45054 11118 45106
rect 11170 45054 11182 45106
rect 13682 45054 13694 45106
rect 13746 45054 13758 45106
rect 18274 45054 18286 45106
rect 18338 45054 18350 45106
rect 26114 45054 26126 45106
rect 26178 45054 26190 45106
rect 27010 45054 27022 45106
rect 27074 45054 27086 45106
rect 27570 45054 27582 45106
rect 27634 45054 27646 45106
rect 31266 45054 31278 45106
rect 31330 45054 31342 45106
rect 34290 45054 34302 45106
rect 34354 45054 34366 45106
rect 35074 45054 35086 45106
rect 35138 45054 35150 45106
rect 37986 45054 37998 45106
rect 38050 45054 38062 45106
rect 39778 45054 39790 45106
rect 39842 45054 39854 45106
rect 42018 45054 42030 45106
rect 42082 45054 42094 45106
rect 42802 45054 42814 45106
rect 42866 45054 42878 45106
rect 30270 45042 30322 45054
rect 33406 44994 33458 45006
rect 30706 44942 30718 44994
rect 30770 44942 30782 44994
rect 33406 44930 33458 44942
rect 33854 44994 33906 45006
rect 33854 44930 33906 44942
rect 39342 44994 39394 45006
rect 39342 44930 39394 44942
rect 41470 44994 41522 45006
rect 45154 44942 45166 44994
rect 45218 44942 45230 44994
rect 41470 44930 41522 44942
rect 10558 44882 10610 44894
rect 10558 44818 10610 44830
rect 17838 44882 17890 44894
rect 25678 44882 25730 44894
rect 20738 44830 20750 44882
rect 20802 44879 20814 44882
rect 21074 44879 21086 44882
rect 20802 44833 21086 44879
rect 20802 44830 20814 44833
rect 21074 44830 21086 44833
rect 21138 44830 21150 44882
rect 17838 44818 17890 44830
rect 25678 44818 25730 44830
rect 1344 44714 48720 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48720 44714
rect 1344 44628 48720 44662
rect 21646 44546 21698 44558
rect 21646 44482 21698 44494
rect 42478 44546 42530 44558
rect 42478 44482 42530 44494
rect 10894 44434 10946 44446
rect 30158 44434 30210 44446
rect 10434 44382 10446 44434
rect 10498 44382 10510 44434
rect 11666 44382 11678 44434
rect 11730 44382 11742 44434
rect 18386 44382 18398 44434
rect 18450 44382 18462 44434
rect 10894 44370 10946 44382
rect 30158 44370 30210 44382
rect 41806 44434 41858 44446
rect 41806 44370 41858 44382
rect 21982 44322 22034 44334
rect 34414 44322 34466 44334
rect 42814 44322 42866 44334
rect 7522 44270 7534 44322
rect 7586 44270 7598 44322
rect 8082 44270 8094 44322
rect 8146 44270 8158 44322
rect 22418 44270 22430 44322
rect 22482 44270 22494 44322
rect 23314 44270 23326 44322
rect 23378 44270 23390 44322
rect 24098 44270 24110 44322
rect 24162 44270 24174 44322
rect 30482 44270 30494 44322
rect 30546 44270 30558 44322
rect 31154 44270 31166 44322
rect 31218 44270 31230 44322
rect 34850 44270 34862 44322
rect 34914 44270 34926 44322
rect 35858 44270 35870 44322
rect 35922 44270 35934 44322
rect 21982 44258 22034 44270
rect 34414 44258 34466 44270
rect 42814 44258 42866 44270
rect 20190 44210 20242 44222
rect 22754 44158 22766 44210
rect 22818 44158 22830 44210
rect 27906 44158 27918 44210
rect 27970 44158 27982 44210
rect 34962 44158 34974 44210
rect 35026 44158 35038 44210
rect 43026 44158 43038 44210
rect 43090 44158 43102 44210
rect 43362 44158 43374 44210
rect 43426 44158 43438 44210
rect 20190 44146 20242 44158
rect 12126 44098 12178 44110
rect 12126 44034 12178 44046
rect 17950 44098 18002 44110
rect 17950 44034 18002 44046
rect 19854 44098 19906 44110
rect 27358 44098 27410 44110
rect 26450 44046 26462 44098
rect 26514 44046 26526 44098
rect 19854 44034 19906 44046
rect 27358 44034 27410 44046
rect 27582 44098 27634 44110
rect 34078 44098 34130 44110
rect 33618 44046 33630 44098
rect 33682 44046 33694 44098
rect 27582 44034 27634 44046
rect 34078 44034 34130 44046
rect 35646 44098 35698 44110
rect 35646 44034 35698 44046
rect 40238 44098 40290 44110
rect 40238 44034 40290 44046
rect 1344 43930 48720 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48720 43930
rect 1344 43844 48720 43878
rect 8094 43762 8146 43774
rect 8094 43698 8146 43710
rect 23102 43762 23154 43774
rect 23102 43698 23154 43710
rect 31166 43762 31218 43774
rect 31166 43698 31218 43710
rect 12238 43650 12290 43662
rect 18734 43650 18786 43662
rect 17938 43598 17950 43650
rect 18002 43598 18014 43650
rect 12238 43586 12290 43598
rect 18734 43586 18786 43598
rect 25230 43650 25282 43662
rect 25230 43586 25282 43598
rect 28254 43650 28306 43662
rect 35198 43650 35250 43662
rect 29250 43598 29262 43650
rect 29314 43598 29326 43650
rect 29810 43598 29822 43650
rect 29874 43598 29886 43650
rect 32274 43598 32286 43650
rect 32338 43598 32350 43650
rect 34290 43598 34302 43650
rect 34354 43598 34366 43650
rect 28254 43586 28306 43598
rect 35198 43586 35250 43598
rect 37998 43650 38050 43662
rect 43150 43650 43202 43662
rect 39330 43598 39342 43650
rect 39394 43598 39406 43650
rect 39890 43598 39902 43650
rect 39954 43598 39966 43650
rect 41458 43598 41470 43650
rect 41522 43598 41534 43650
rect 37998 43586 38050 43598
rect 43150 43586 43202 43598
rect 8430 43538 8482 43550
rect 28702 43538 28754 43550
rect 34862 43538 34914 43550
rect 4722 43486 4734 43538
rect 4786 43486 4798 43538
rect 5282 43486 5294 43538
rect 5346 43486 5358 43538
rect 12002 43486 12014 43538
rect 12066 43486 12078 43538
rect 12674 43486 12686 43538
rect 12738 43486 12750 43538
rect 13122 43486 13134 43538
rect 13186 43486 13198 43538
rect 18162 43486 18174 43538
rect 18226 43486 18238 43538
rect 18946 43486 18958 43538
rect 19010 43486 19022 43538
rect 19618 43486 19630 43538
rect 19682 43486 19694 43538
rect 25442 43486 25454 43538
rect 25506 43486 25518 43538
rect 28018 43486 28030 43538
rect 28082 43486 28094 43538
rect 32050 43486 32062 43538
rect 32114 43486 32126 43538
rect 34066 43486 34078 43538
rect 34130 43486 34142 43538
rect 8430 43474 8482 43486
rect 28702 43474 28754 43486
rect 34862 43474 34914 43486
rect 38334 43538 38386 43550
rect 38334 43474 38386 43486
rect 38782 43538 38834 43550
rect 42814 43538 42866 43550
rect 41346 43486 41358 43538
rect 41410 43486 41422 43538
rect 38782 43474 38834 43486
rect 42814 43474 42866 43486
rect 8878 43426 8930 43438
rect 7634 43374 7646 43426
rect 7698 43374 7710 43426
rect 8878 43362 8930 43374
rect 11566 43426 11618 43438
rect 17614 43426 17666 43438
rect 15586 43374 15598 43426
rect 15650 43374 15662 43426
rect 22082 43374 22094 43426
rect 22146 43374 22158 43426
rect 11566 43362 11618 43374
rect 17614 43362 17666 43374
rect 29038 43314 29090 43326
rect 29038 43250 29090 43262
rect 31502 43314 31554 43326
rect 31502 43250 31554 43262
rect 39118 43314 39170 43326
rect 39118 43250 39170 43262
rect 42030 43314 42082 43326
rect 42030 43250 42082 43262
rect 42366 43314 42418 43326
rect 42366 43250 42418 43262
rect 1344 43146 48720 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48720 43146
rect 1344 43060 48720 43094
rect 8654 42978 8706 42990
rect 8654 42914 8706 42926
rect 13582 42978 13634 42990
rect 13582 42914 13634 42926
rect 21422 42978 21474 42990
rect 21422 42914 21474 42926
rect 42702 42978 42754 42990
rect 42702 42914 42754 42926
rect 18846 42866 18898 42878
rect 10658 42814 10670 42866
rect 10722 42814 10734 42866
rect 18846 42802 18898 42814
rect 23550 42866 23602 42878
rect 23550 42802 23602 42814
rect 36318 42866 36370 42878
rect 36318 42802 36370 42814
rect 8990 42754 9042 42766
rect 11118 42754 11170 42766
rect 9762 42702 9774 42754
rect 9826 42702 9838 42754
rect 8990 42690 9042 42702
rect 11118 42690 11170 42702
rect 11454 42754 11506 42766
rect 11454 42690 11506 42702
rect 12014 42754 12066 42766
rect 12014 42690 12066 42702
rect 13918 42754 13970 42766
rect 21758 42754 21810 42766
rect 43038 42754 43090 42766
rect 14354 42702 14366 42754
rect 14418 42702 14430 42754
rect 15474 42702 15486 42754
rect 15538 42702 15550 42754
rect 16034 42702 16046 42754
rect 16098 42702 16110 42754
rect 18386 42702 18398 42754
rect 18450 42702 18462 42754
rect 22194 42702 22206 42754
rect 22258 42702 22270 42754
rect 23762 42702 23774 42754
rect 23826 42702 23838 42754
rect 24546 42702 24558 42754
rect 24610 42702 24622 42754
rect 37762 42702 37774 42754
rect 37826 42702 37838 42754
rect 38210 42702 38222 42754
rect 38274 42702 38286 42754
rect 43474 42702 43486 42754
rect 43538 42702 43550 42754
rect 13918 42690 13970 42702
rect 21758 42690 21810 42702
rect 43038 42690 43090 42702
rect 5630 42642 5682 42654
rect 5630 42578 5682 42590
rect 5966 42642 6018 42654
rect 35310 42642 35362 42654
rect 9650 42590 9662 42642
rect 9714 42590 9726 42642
rect 14690 42590 14702 42642
rect 14754 42590 14766 42642
rect 22530 42590 22542 42642
rect 22594 42590 22606 42642
rect 43810 42590 43822 42642
rect 43874 42590 43886 42642
rect 5966 42578 6018 42590
rect 35310 42578 35362 42590
rect 35646 42530 35698 42542
rect 41134 42530 41186 42542
rect 26898 42478 26910 42530
rect 26962 42478 26974 42530
rect 40674 42478 40686 42530
rect 40738 42478 40750 42530
rect 35646 42466 35698 42478
rect 41134 42466 41186 42478
rect 1344 42362 48720 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48720 42362
rect 1344 42276 48720 42310
rect 6526 42194 6578 42206
rect 6526 42130 6578 42142
rect 18958 42194 19010 42206
rect 18958 42130 19010 42142
rect 25342 42194 25394 42206
rect 45714 42142 45726 42194
rect 45778 42142 45790 42194
rect 25342 42130 25394 42142
rect 9998 42082 10050 42094
rect 31054 42082 31106 42094
rect 7634 42030 7646 42082
rect 7698 42030 7710 42082
rect 26226 42030 26238 42082
rect 26290 42030 26302 42082
rect 9998 42018 10050 42030
rect 31054 42018 31106 42030
rect 39790 42082 39842 42094
rect 39790 42018 39842 42030
rect 9662 41970 9714 41982
rect 41022 41970 41074 41982
rect 7522 41918 7534 41970
rect 7586 41918 7598 41970
rect 19170 41918 19182 41970
rect 19234 41918 19246 41970
rect 19954 41918 19966 41970
rect 20018 41918 20030 41970
rect 26114 41918 26126 41970
rect 26178 41918 26190 41970
rect 27794 41918 27806 41970
rect 27858 41918 27870 41970
rect 28242 41918 28254 41970
rect 28306 41918 28318 41970
rect 31266 41918 31278 41970
rect 31330 41918 31342 41970
rect 32946 41918 32958 41970
rect 33010 41918 33022 41970
rect 33618 41918 33630 41970
rect 33682 41918 33694 41970
rect 38770 41918 38782 41970
rect 38834 41918 38846 41970
rect 39330 41918 39342 41970
rect 39394 41918 39406 41970
rect 40002 41918 40014 41970
rect 40066 41918 40078 41970
rect 9662 41906 9714 41918
rect 41022 41906 41074 41918
rect 42366 41970 42418 41982
rect 42578 41918 42590 41970
rect 42642 41918 42654 41970
rect 43250 41918 43262 41970
rect 43314 41918 43326 41970
rect 42366 41906 42418 41918
rect 31838 41858 31890 41870
rect 22306 41806 22318 41858
rect 22370 41806 22382 41858
rect 30706 41806 30718 41858
rect 30770 41806 30782 41858
rect 36082 41806 36094 41858
rect 36146 41806 36158 41858
rect 36418 41806 36430 41858
rect 36482 41806 36494 41858
rect 31838 41794 31890 41806
rect 6862 41746 6914 41758
rect 6862 41682 6914 41694
rect 25678 41746 25730 41758
rect 25678 41682 25730 41694
rect 1344 41578 48720 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48720 41578
rect 1344 41492 48720 41526
rect 34974 41410 35026 41422
rect 34974 41346 35026 41358
rect 35310 41410 35362 41422
rect 35310 41346 35362 41358
rect 19630 41298 19682 41310
rect 19170 41246 19182 41298
rect 19234 41246 19246 41298
rect 19630 41234 19682 41246
rect 26686 41298 26738 41310
rect 26686 41234 26738 41246
rect 27694 41298 27746 41310
rect 27694 41234 27746 41246
rect 15038 41186 15090 41198
rect 21758 41186 21810 41198
rect 33406 41186 33458 41198
rect 38446 41186 38498 41198
rect 42590 41186 42642 41198
rect 6626 41134 6638 41186
rect 6690 41134 6702 41186
rect 9314 41134 9326 41186
rect 9378 41134 9390 41186
rect 9986 41134 9998 41186
rect 10050 41134 10062 41186
rect 16258 41134 16270 41186
rect 16322 41134 16334 41186
rect 16818 41134 16830 41186
rect 16882 41134 16894 41186
rect 22194 41134 22206 41186
rect 22258 41134 22270 41186
rect 29586 41134 29598 41186
rect 29650 41134 29662 41186
rect 30146 41134 30158 41186
rect 30210 41134 30222 41186
rect 34066 41134 34078 41186
rect 34130 41134 34142 41186
rect 38882 41134 38894 41186
rect 38946 41134 38958 41186
rect 39442 41134 39454 41186
rect 39506 41134 39518 41186
rect 15038 41122 15090 41134
rect 21758 41122 21810 41134
rect 33406 41122 33458 41134
rect 38446 41122 38498 41134
rect 42590 41122 42642 41134
rect 15262 41074 15314 41086
rect 15262 41010 15314 41022
rect 20190 41074 20242 41086
rect 20190 41010 20242 41022
rect 20526 41074 20578 41086
rect 20526 41010 20578 41022
rect 21422 41074 21474 41086
rect 24446 41074 24498 41086
rect 22418 41022 22430 41074
rect 22482 41022 22494 41074
rect 34178 41022 34190 41074
rect 34242 41022 34254 41074
rect 35522 41022 35534 41074
rect 35586 41022 35598 41074
rect 36082 41022 36094 41074
rect 36146 41022 36158 41074
rect 42802 41022 42814 41074
rect 42866 41022 42878 41074
rect 43138 41022 43150 41074
rect 43202 41022 43214 41074
rect 21422 41010 21474 41022
rect 24446 41010 24498 41022
rect 6414 40962 6466 40974
rect 12910 40962 12962 40974
rect 12450 40910 12462 40962
rect 12514 40910 12526 40962
rect 6414 40898 6466 40910
rect 12910 40898 12962 40910
rect 14366 40962 14418 40974
rect 14366 40898 14418 40910
rect 14478 40962 14530 40974
rect 14478 40898 14530 40910
rect 14590 40962 14642 40974
rect 14590 40898 14642 40910
rect 15374 40962 15426 40974
rect 15374 40898 15426 40910
rect 23102 40962 23154 40974
rect 23102 40898 23154 40910
rect 24110 40962 24162 40974
rect 24110 40898 24162 40910
rect 27246 40962 27298 40974
rect 33070 40962 33122 40974
rect 42254 40962 42306 40974
rect 32498 40910 32510 40962
rect 32562 40910 32574 40962
rect 41794 40910 41806 40962
rect 41858 40910 41870 40962
rect 27246 40898 27298 40910
rect 33070 40898 33122 40910
rect 42254 40898 42306 40910
rect 1344 40794 48720 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48720 40794
rect 1344 40708 48720 40742
rect 9662 40626 9714 40638
rect 15486 40626 15538 40638
rect 15250 40574 15262 40626
rect 15314 40574 15326 40626
rect 9662 40562 9714 40574
rect 15486 40562 15538 40574
rect 22990 40626 23042 40638
rect 22990 40562 23042 40574
rect 25342 40626 25394 40638
rect 25342 40562 25394 40574
rect 30718 40626 30770 40638
rect 30718 40562 30770 40574
rect 33406 40626 33458 40638
rect 33406 40562 33458 40574
rect 39118 40626 39170 40638
rect 39118 40562 39170 40574
rect 41694 40626 41746 40638
rect 41694 40562 41746 40574
rect 15710 40514 15762 40526
rect 33070 40514 33122 40526
rect 8978 40462 8990 40514
rect 9042 40462 9054 40514
rect 10546 40462 10558 40514
rect 10610 40462 10622 40514
rect 17602 40462 17614 40514
rect 17666 40462 17678 40514
rect 26450 40462 26462 40514
rect 26514 40462 26526 40514
rect 31602 40462 31614 40514
rect 31666 40462 31678 40514
rect 40002 40462 40014 40514
rect 40066 40462 40078 40514
rect 15710 40450 15762 40462
rect 33070 40450 33122 40462
rect 15822 40402 15874 40414
rect 2370 40350 2382 40402
rect 2434 40350 2446 40402
rect 3154 40350 3166 40402
rect 3218 40350 3230 40402
rect 5506 40350 5518 40402
rect 5570 40350 5582 40402
rect 5842 40350 5854 40402
rect 5906 40350 5918 40402
rect 6514 40350 6526 40402
rect 6578 40350 6590 40402
rect 10658 40350 10670 40402
rect 10722 40350 10734 40402
rect 12114 40350 12126 40402
rect 12178 40350 12190 40402
rect 12786 40350 12798 40402
rect 12850 40350 12862 40402
rect 15822 40338 15874 40350
rect 16270 40402 16322 40414
rect 18286 40402 18338 40414
rect 17490 40350 17502 40402
rect 17554 40350 17566 40402
rect 16270 40338 16322 40350
rect 18286 40338 18338 40350
rect 19182 40402 19234 40414
rect 19182 40338 19234 40350
rect 20190 40402 20242 40414
rect 20190 40338 20242 40350
rect 23550 40402 23602 40414
rect 32510 40402 32562 40414
rect 26338 40350 26350 40402
rect 26402 40350 26414 40402
rect 27346 40350 27358 40402
rect 27410 40350 27422 40402
rect 27906 40350 27918 40402
rect 27970 40350 27982 40402
rect 31714 40350 31726 40402
rect 31778 40350 31790 40402
rect 40114 40350 40126 40402
rect 40178 40350 40190 40402
rect 41906 40350 41918 40402
rect 41970 40350 41982 40402
rect 42578 40350 42590 40402
rect 42642 40350 42654 40402
rect 45042 40350 45054 40402
rect 45106 40350 45118 40402
rect 23550 40338 23602 40350
rect 32510 40338 32562 40350
rect 19742 40290 19794 40302
rect 19742 40226 19794 40238
rect 20974 40290 21026 40302
rect 20974 40226 21026 40238
rect 21758 40290 21810 40302
rect 21758 40226 21810 40238
rect 24222 40290 24274 40302
rect 24222 40226 24274 40238
rect 24670 40290 24722 40302
rect 30258 40238 30270 40290
rect 30322 40238 30334 40290
rect 24670 40226 24722 40238
rect 9998 40178 10050 40190
rect 9998 40114 10050 40126
rect 18622 40178 18674 40190
rect 25678 40178 25730 40190
rect 19170 40126 19182 40178
rect 19234 40175 19246 40178
rect 19730 40175 19742 40178
rect 19234 40129 19742 40175
rect 19234 40126 19246 40129
rect 19730 40126 19742 40129
rect 19794 40126 19806 40178
rect 18622 40114 18674 40126
rect 25678 40114 25730 40126
rect 31054 40178 31106 40190
rect 31054 40114 31106 40126
rect 39454 40178 39506 40190
rect 39454 40114 39506 40126
rect 1344 40010 48720 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48720 40010
rect 1344 39924 48720 39958
rect 6750 39842 6802 39854
rect 6750 39778 6802 39790
rect 7086 39842 7138 39854
rect 7086 39778 7138 39790
rect 12238 39842 12290 39854
rect 12238 39778 12290 39790
rect 30494 39730 30546 39742
rect 34962 39678 34974 39730
rect 35026 39678 35038 39730
rect 30494 39666 30546 39678
rect 22094 39618 22146 39630
rect 42254 39618 42306 39630
rect 7522 39566 7534 39618
rect 7586 39566 7598 39618
rect 16930 39566 16942 39618
rect 16994 39566 17006 39618
rect 17490 39566 17502 39618
rect 17554 39566 17566 39618
rect 20514 39566 20526 39618
rect 20578 39566 20590 39618
rect 23314 39566 23326 39618
rect 23378 39566 23390 39618
rect 24098 39566 24110 39618
rect 24162 39566 24174 39618
rect 28130 39566 28142 39618
rect 28194 39566 28206 39618
rect 37090 39566 37102 39618
rect 37154 39566 37166 39618
rect 22094 39554 22146 39566
rect 42254 39554 42306 39566
rect 3278 39506 3330 39518
rect 3278 39442 3330 39454
rect 3614 39506 3666 39518
rect 12462 39506 12514 39518
rect 7634 39454 7646 39506
rect 7698 39454 7710 39506
rect 3614 39442 3666 39454
rect 12462 39442 12514 39454
rect 14030 39506 14082 39518
rect 14030 39442 14082 39454
rect 14702 39506 14754 39518
rect 14702 39442 14754 39454
rect 21758 39506 21810 39518
rect 27918 39506 27970 39518
rect 22306 39454 22318 39506
rect 22370 39454 22382 39506
rect 22866 39454 22878 39506
rect 22930 39454 22942 39506
rect 21758 39442 21810 39454
rect 27918 39442 27970 39454
rect 42590 39506 42642 39518
rect 42590 39442 42642 39454
rect 5742 39394 5794 39406
rect 5742 39330 5794 39342
rect 9214 39394 9266 39406
rect 9214 39330 9266 39342
rect 11678 39394 11730 39406
rect 13022 39394 13074 39406
rect 11890 39342 11902 39394
rect 11954 39342 11966 39394
rect 11678 39330 11730 39342
rect 13022 39330 13074 39342
rect 13694 39394 13746 39406
rect 13694 39330 13746 39342
rect 14366 39394 14418 39406
rect 14366 39330 14418 39342
rect 14590 39394 14642 39406
rect 20750 39394 20802 39406
rect 27134 39394 27186 39406
rect 34526 39394 34578 39406
rect 19842 39342 19854 39394
rect 19906 39342 19918 39394
rect 26450 39342 26462 39394
rect 26514 39342 26526 39394
rect 27458 39342 27470 39394
rect 27522 39342 27534 39394
rect 14590 39330 14642 39342
rect 20750 39330 20802 39342
rect 27134 39330 27186 39342
rect 34526 39330 34578 39342
rect 37326 39394 37378 39406
rect 37326 39330 37378 39342
rect 40350 39394 40402 39406
rect 40350 39330 40402 39342
rect 1344 39226 48720 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48720 39226
rect 1344 39140 48720 39174
rect 11566 39058 11618 39070
rect 8978 39006 8990 39058
rect 9042 39006 9054 39058
rect 11566 38994 11618 39006
rect 11790 39058 11842 39070
rect 11790 38994 11842 39006
rect 17502 39058 17554 39070
rect 28142 39058 28194 39070
rect 23202 39006 23214 39058
rect 23266 39006 23278 39058
rect 17502 38994 17554 39006
rect 28142 38994 28194 39006
rect 11902 38946 11954 38958
rect 11902 38882 11954 38894
rect 17614 38946 17666 38958
rect 17614 38882 17666 38894
rect 18510 38946 18562 38958
rect 18510 38882 18562 38894
rect 18622 38946 18674 38958
rect 18622 38882 18674 38894
rect 19630 38946 19682 38958
rect 30830 38946 30882 38958
rect 39566 38946 39618 38958
rect 28690 38894 28702 38946
rect 28754 38894 28766 38946
rect 29026 38894 29038 38946
rect 29090 38894 29102 38946
rect 31938 38894 31950 38946
rect 32002 38894 32014 38946
rect 32274 38894 32286 38946
rect 32338 38894 32350 38946
rect 34738 38894 34750 38946
rect 34802 38894 34814 38946
rect 35074 38894 35086 38946
rect 35138 38894 35150 38946
rect 19630 38882 19682 38894
rect 30830 38882 30882 38894
rect 39566 38882 39618 38894
rect 41246 38946 41298 38958
rect 41246 38882 41298 38894
rect 5182 38834 5234 38846
rect 9662 38834 9714 38846
rect 1810 38782 1822 38834
rect 1874 38782 1886 38834
rect 2258 38782 2270 38834
rect 2322 38782 2334 38834
rect 5842 38782 5854 38834
rect 5906 38782 5918 38834
rect 6626 38782 6638 38834
rect 6690 38782 6702 38834
rect 5182 38770 5234 38782
rect 9662 38770 9714 38782
rect 10782 38834 10834 38846
rect 17390 38834 17442 38846
rect 12226 38782 12238 38834
rect 12290 38782 12302 38834
rect 12674 38782 12686 38834
rect 12738 38782 12750 38834
rect 13346 38782 13358 38834
rect 13410 38782 13422 38834
rect 10782 38770 10834 38782
rect 17390 38770 17442 38782
rect 18062 38834 18114 38846
rect 18062 38770 18114 38782
rect 18846 38834 18898 38846
rect 18846 38770 18898 38782
rect 19518 38834 19570 38846
rect 24334 38834 24386 38846
rect 20178 38782 20190 38834
rect 20242 38782 20254 38834
rect 20738 38782 20750 38834
rect 20802 38782 20814 38834
rect 19518 38770 19570 38782
rect 24334 38770 24386 38782
rect 26014 38834 26066 38846
rect 31614 38834 31666 38846
rect 27234 38782 27246 38834
rect 27298 38782 27310 38834
rect 30594 38782 30606 38834
rect 30658 38782 30670 38834
rect 26014 38770 26066 38782
rect 31614 38770 31666 38782
rect 34526 38834 34578 38846
rect 39230 38834 39282 38846
rect 38210 38782 38222 38834
rect 38274 38782 38286 38834
rect 38994 38782 39006 38834
rect 39058 38782 39070 38834
rect 41010 38782 41022 38834
rect 41074 38782 41086 38834
rect 34526 38770 34578 38782
rect 39230 38770 39282 38782
rect 11342 38722 11394 38734
rect 16046 38722 16098 38734
rect 4722 38670 4734 38722
rect 4786 38670 4798 38722
rect 12338 38670 12350 38722
rect 12402 38670 12414 38722
rect 15698 38670 15710 38722
rect 15762 38670 15774 38722
rect 11342 38658 11394 38670
rect 16046 38658 16098 38670
rect 16158 38722 16210 38734
rect 16158 38658 16210 38670
rect 19294 38722 19346 38734
rect 19294 38658 19346 38670
rect 23774 38722 23826 38734
rect 23774 38658 23826 38670
rect 24110 38722 24162 38734
rect 24110 38658 24162 38670
rect 25454 38722 25506 38734
rect 25454 38658 25506 38670
rect 25790 38722 25842 38734
rect 25790 38658 25842 38670
rect 26798 38722 26850 38734
rect 26798 38658 26850 38670
rect 27694 38722 27746 38734
rect 27694 38658 27746 38670
rect 31278 38722 31330 38734
rect 40014 38722 40066 38734
rect 35858 38670 35870 38722
rect 35922 38670 35934 38722
rect 31278 38658 31330 38670
rect 40014 38658 40066 38670
rect 24670 38610 24722 38622
rect 24670 38546 24722 38558
rect 26350 38610 26402 38622
rect 26350 38546 26402 38558
rect 28478 38610 28530 38622
rect 28478 38546 28530 38558
rect 34190 38610 34242 38622
rect 34190 38546 34242 38558
rect 1344 38442 48720 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48720 38442
rect 1344 38356 48720 38390
rect 3838 38274 3890 38286
rect 3838 38210 3890 38222
rect 10558 38274 10610 38286
rect 10558 38210 10610 38222
rect 37102 38274 37154 38286
rect 37102 38210 37154 38222
rect 37438 38274 37490 38286
rect 37438 38210 37490 38222
rect 38782 38274 38834 38286
rect 38782 38210 38834 38222
rect 6078 38162 6130 38174
rect 6078 38098 6130 38110
rect 9662 38162 9714 38174
rect 14142 38162 14194 38174
rect 12226 38110 12238 38162
rect 12290 38110 12302 38162
rect 9662 38098 9714 38110
rect 14142 38098 14194 38110
rect 14814 38162 14866 38174
rect 14814 38098 14866 38110
rect 16718 38162 16770 38174
rect 16718 38098 16770 38110
rect 17614 38162 17666 38174
rect 17614 38098 17666 38110
rect 21646 38162 21698 38174
rect 22990 38162 23042 38174
rect 22418 38110 22430 38162
rect 22482 38110 22494 38162
rect 21646 38098 21698 38110
rect 22990 38098 23042 38110
rect 24110 38162 24162 38174
rect 27794 38110 27806 38162
rect 27858 38110 27870 38162
rect 33842 38110 33854 38162
rect 33906 38110 33918 38162
rect 24110 38098 24162 38110
rect 4174 38050 4226 38062
rect 13694 38050 13746 38062
rect 17166 38050 17218 38062
rect 19742 38050 19794 38062
rect 23214 38050 23266 38062
rect 26686 38050 26738 38062
rect 28142 38050 28194 38062
rect 39118 38050 39170 38062
rect 4834 37998 4846 38050
rect 4898 37998 4910 38050
rect 11442 37998 11454 38050
rect 11506 37998 11518 38050
rect 12338 37998 12350 38050
rect 12402 37998 12414 38050
rect 14354 37998 14366 38050
rect 14418 37998 14430 38050
rect 18946 37998 18958 38050
rect 19010 37998 19022 38050
rect 19170 37998 19182 38050
rect 19234 37998 19246 38050
rect 20066 37998 20078 38050
rect 20130 37998 20142 38050
rect 25330 37998 25342 38050
rect 25394 37998 25406 38050
rect 25666 37998 25678 38050
rect 25730 37998 25742 38050
rect 27458 37998 27470 38050
rect 27522 37998 27534 38050
rect 27682 37998 27694 38050
rect 27746 37998 27758 38050
rect 30930 37998 30942 38050
rect 30994 37998 31006 38050
rect 31378 37998 31390 38050
rect 31442 37998 31454 38050
rect 35410 37998 35422 38050
rect 35474 37998 35486 38050
rect 39778 37998 39790 38050
rect 39842 37998 39854 38050
rect 40562 37998 40574 38050
rect 40626 37998 40638 38050
rect 41234 37998 41246 38050
rect 41298 37998 41310 38050
rect 4174 37986 4226 37998
rect 13694 37986 13746 37998
rect 17166 37986 17218 37998
rect 19742 37986 19794 37998
rect 23214 37986 23266 37998
rect 26686 37986 26738 37998
rect 28142 37986 28194 37998
rect 39118 37986 39170 37998
rect 2270 37938 2322 37950
rect 2270 37874 2322 37886
rect 2606 37938 2658 37950
rect 5742 37938 5794 37950
rect 7422 37938 7474 37950
rect 4946 37886 4958 37938
rect 5010 37886 5022 37938
rect 6290 37886 6302 37938
rect 6354 37886 6366 37938
rect 6850 37886 6862 37938
rect 6914 37886 6926 37938
rect 2606 37874 2658 37886
rect 5742 37874 5794 37886
rect 7422 37874 7474 37886
rect 7758 37938 7810 37950
rect 7758 37874 7810 37886
rect 9438 37938 9490 37950
rect 9438 37874 9490 37886
rect 10334 37938 10386 37950
rect 10334 37874 10386 37886
rect 11230 37938 11282 37950
rect 16270 37938 16322 37950
rect 12450 37886 12462 37938
rect 12514 37886 12526 37938
rect 11230 37874 11282 37886
rect 16270 37874 16322 37886
rect 16606 37938 16658 37950
rect 16606 37874 16658 37886
rect 16942 37938 16994 37950
rect 16942 37874 16994 37886
rect 17502 37938 17554 37950
rect 17502 37874 17554 37886
rect 17726 37938 17778 37950
rect 17726 37874 17778 37886
rect 20414 37938 20466 37950
rect 20414 37874 20466 37886
rect 20526 37938 20578 37950
rect 20526 37874 20578 37886
rect 24558 37938 24610 37950
rect 24558 37874 24610 37886
rect 24670 37938 24722 37950
rect 24670 37874 24722 37886
rect 26574 37938 26626 37950
rect 26574 37874 26626 37886
rect 35870 37938 35922 37950
rect 37650 37886 37662 37938
rect 37714 37886 37726 37938
rect 37986 37886 37998 37938
rect 38050 37886 38062 37938
rect 39890 37886 39902 37938
rect 39954 37886 39966 37938
rect 35870 37874 35922 37886
rect 14702 37826 14754 37838
rect 9986 37774 9998 37826
rect 10050 37774 10062 37826
rect 10882 37774 10894 37826
rect 10946 37774 10958 37826
rect 14702 37762 14754 37774
rect 14926 37826 14978 37838
rect 14926 37762 14978 37774
rect 15486 37826 15538 37838
rect 15486 37762 15538 37774
rect 18734 37826 18786 37838
rect 18734 37762 18786 37774
rect 19406 37826 19458 37838
rect 19406 37762 19458 37774
rect 19518 37826 19570 37838
rect 19518 37762 19570 37774
rect 19854 37826 19906 37838
rect 19854 37762 19906 37774
rect 20750 37826 20802 37838
rect 20750 37762 20802 37774
rect 21982 37826 22034 37838
rect 24334 37826 24386 37838
rect 23538 37774 23550 37826
rect 23602 37774 23614 37826
rect 21982 37762 22034 37774
rect 24334 37762 24386 37774
rect 25902 37826 25954 37838
rect 25902 37762 25954 37774
rect 26014 37826 26066 37838
rect 26014 37762 26066 37774
rect 26126 37826 26178 37838
rect 26126 37762 26178 37774
rect 26350 37826 26402 37838
rect 26350 37762 26402 37774
rect 27918 37826 27970 37838
rect 27918 37762 27970 37774
rect 29710 37826 29762 37838
rect 29710 37762 29762 37774
rect 34302 37826 34354 37838
rect 44158 37826 44210 37838
rect 43698 37774 43710 37826
rect 43762 37774 43774 37826
rect 34302 37762 34354 37774
rect 44158 37762 44210 37774
rect 1344 37658 48720 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48720 37658
rect 1344 37572 48720 37606
rect 5182 37490 5234 37502
rect 5182 37426 5234 37438
rect 10222 37490 10274 37502
rect 10222 37426 10274 37438
rect 15486 37490 15538 37502
rect 15486 37426 15538 37438
rect 16382 37490 16434 37502
rect 16382 37426 16434 37438
rect 24334 37490 24386 37502
rect 24334 37426 24386 37438
rect 24558 37490 24610 37502
rect 24558 37426 24610 37438
rect 25566 37490 25618 37502
rect 25566 37426 25618 37438
rect 25790 37490 25842 37502
rect 25790 37426 25842 37438
rect 26462 37490 26514 37502
rect 26462 37426 26514 37438
rect 41134 37490 41186 37502
rect 41134 37426 41186 37438
rect 10110 37378 10162 37390
rect 10110 37314 10162 37326
rect 10894 37378 10946 37390
rect 10894 37314 10946 37326
rect 11006 37378 11058 37390
rect 13918 37378 13970 37390
rect 12002 37326 12014 37378
rect 12066 37326 12078 37378
rect 11006 37314 11058 37326
rect 13918 37314 13970 37326
rect 15038 37378 15090 37390
rect 29486 37378 29538 37390
rect 43150 37378 43202 37390
rect 18274 37326 18286 37378
rect 18338 37326 18350 37378
rect 42242 37326 42254 37378
rect 42306 37326 42318 37378
rect 15038 37314 15090 37326
rect 29486 37314 29538 37326
rect 43150 37314 43202 37326
rect 9102 37266 9154 37278
rect 1810 37214 1822 37266
rect 1874 37214 1886 37266
rect 2370 37214 2382 37266
rect 2434 37214 2446 37266
rect 9102 37202 9154 37214
rect 10446 37266 10498 37278
rect 10446 37202 10498 37214
rect 10670 37266 10722 37278
rect 11790 37266 11842 37278
rect 13470 37266 13522 37278
rect 11330 37214 11342 37266
rect 11394 37214 11406 37266
rect 12450 37214 12462 37266
rect 12514 37214 12526 37266
rect 13234 37214 13246 37266
rect 13298 37214 13310 37266
rect 10670 37202 10722 37214
rect 11790 37202 11842 37214
rect 13470 37202 13522 37214
rect 14142 37266 14194 37278
rect 14142 37202 14194 37214
rect 15598 37266 15650 37278
rect 15598 37202 15650 37214
rect 16046 37266 16098 37278
rect 16046 37202 16098 37214
rect 16382 37266 16434 37278
rect 16382 37202 16434 37214
rect 16718 37266 16770 37278
rect 22766 37266 22818 37278
rect 25342 37266 25394 37278
rect 20066 37214 20078 37266
rect 20130 37214 20142 37266
rect 22194 37214 22206 37266
rect 22258 37214 22270 37266
rect 23090 37214 23102 37266
rect 23154 37214 23166 37266
rect 23874 37214 23886 37266
rect 23938 37214 23950 37266
rect 24098 37214 24110 37266
rect 24162 37214 24174 37266
rect 16718 37202 16770 37214
rect 22766 37202 22818 37214
rect 25342 37202 25394 37214
rect 26014 37266 26066 37278
rect 26014 37202 26066 37214
rect 27022 37266 27074 37278
rect 27022 37202 27074 37214
rect 28926 37266 28978 37278
rect 30046 37266 30098 37278
rect 41470 37266 41522 37278
rect 29250 37214 29262 37266
rect 29314 37214 29326 37266
rect 33058 37214 33070 37266
rect 33122 37214 33134 37266
rect 39666 37214 39678 37266
rect 39730 37214 39742 37266
rect 40450 37214 40462 37266
rect 40514 37214 40526 37266
rect 41906 37214 41918 37266
rect 41970 37214 41982 37266
rect 42914 37214 42926 37266
rect 42978 37214 42990 37266
rect 43362 37214 43374 37266
rect 43426 37214 43438 37266
rect 44034 37214 44046 37266
rect 44098 37214 44110 37266
rect 28926 37202 28978 37214
rect 30046 37202 30098 37214
rect 41470 37202 41522 37214
rect 9886 37154 9938 37166
rect 13694 37154 13746 37166
rect 4722 37102 4734 37154
rect 4786 37102 4798 37154
rect 11442 37102 11454 37154
rect 11506 37102 11518 37154
rect 9886 37090 9938 37102
rect 13694 37090 13746 37102
rect 14702 37154 14754 37166
rect 14702 37090 14754 37102
rect 20638 37154 20690 37166
rect 20638 37090 20690 37102
rect 21310 37154 21362 37166
rect 26126 37154 26178 37166
rect 22306 37102 22318 37154
rect 22370 37102 22382 37154
rect 23762 37102 23774 37154
rect 23826 37102 23838 37154
rect 21310 37090 21362 37102
rect 26126 37090 26178 37102
rect 28254 37154 28306 37166
rect 28254 37090 28306 37102
rect 28702 37154 28754 37166
rect 28702 37090 28754 37102
rect 29822 37154 29874 37166
rect 29822 37090 29874 37102
rect 30830 37154 30882 37166
rect 30830 37090 30882 37102
rect 31726 37154 31778 37166
rect 31726 37090 31778 37102
rect 32062 37154 32114 37166
rect 32062 37090 32114 37102
rect 32510 37154 32562 37166
rect 34514 37102 34526 37154
rect 34578 37102 34590 37154
rect 37314 37102 37326 37154
rect 37378 37102 37390 37154
rect 46498 37102 46510 37154
rect 46562 37102 46574 37154
rect 32510 37090 32562 37102
rect 13358 37042 13410 37054
rect 13358 36978 13410 36990
rect 15710 37042 15762 37054
rect 29150 37042 29202 37054
rect 22082 36990 22094 37042
rect 22146 36990 22158 37042
rect 15710 36978 15762 36990
rect 29150 36978 29202 36990
rect 30382 37042 30434 37054
rect 30382 36978 30434 36990
rect 1344 36874 48720 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48720 36874
rect 1344 36788 48720 36822
rect 8206 36706 8258 36718
rect 8206 36642 8258 36654
rect 19854 36706 19906 36718
rect 19854 36642 19906 36654
rect 24894 36706 24946 36718
rect 24894 36642 24946 36654
rect 32398 36706 32450 36718
rect 32398 36642 32450 36654
rect 43038 36706 43090 36718
rect 43038 36642 43090 36654
rect 43374 36706 43426 36718
rect 43374 36642 43426 36654
rect 37438 36594 37490 36606
rect 11218 36542 11230 36594
rect 11282 36542 11294 36594
rect 33170 36542 33182 36594
rect 33234 36542 33246 36594
rect 37438 36530 37490 36542
rect 6078 36482 6130 36494
rect 6078 36418 6130 36430
rect 8542 36482 8594 36494
rect 8542 36418 8594 36430
rect 10670 36482 10722 36494
rect 10670 36418 10722 36430
rect 12350 36482 12402 36494
rect 12350 36418 12402 36430
rect 12574 36482 12626 36494
rect 12574 36418 12626 36430
rect 12798 36482 12850 36494
rect 12798 36418 12850 36430
rect 12910 36482 12962 36494
rect 19406 36482 19458 36494
rect 23326 36482 23378 36494
rect 14018 36430 14030 36482
rect 14082 36430 14094 36482
rect 15138 36430 15150 36482
rect 15202 36430 15214 36482
rect 15586 36430 15598 36482
rect 15650 36430 15662 36482
rect 16146 36430 16158 36482
rect 16210 36430 16222 36482
rect 19954 36430 19966 36482
rect 20018 36430 20030 36482
rect 21522 36430 21534 36482
rect 21586 36430 21598 36482
rect 22082 36430 22094 36482
rect 22146 36430 22158 36482
rect 22530 36430 22542 36482
rect 22594 36430 22606 36482
rect 12910 36418 12962 36430
rect 19406 36418 19458 36430
rect 23326 36418 23378 36430
rect 23550 36482 23602 36494
rect 23550 36418 23602 36430
rect 25118 36482 25170 36494
rect 25118 36418 25170 36430
rect 26014 36482 26066 36494
rect 26014 36418 26066 36430
rect 26238 36482 26290 36494
rect 26238 36418 26290 36430
rect 27582 36482 27634 36494
rect 27582 36418 27634 36430
rect 27806 36482 27858 36494
rect 27806 36418 27858 36430
rect 28142 36482 28194 36494
rect 28142 36418 28194 36430
rect 29710 36482 29762 36494
rect 30370 36430 30382 36482
rect 30434 36430 30446 36482
rect 33506 36430 33518 36482
rect 33570 36430 33582 36482
rect 34402 36430 34414 36482
rect 34466 36430 34478 36482
rect 35298 36430 35310 36482
rect 35362 36430 35374 36482
rect 29710 36418 29762 36430
rect 2494 36370 2546 36382
rect 2494 36306 2546 36318
rect 2830 36370 2882 36382
rect 2830 36306 2882 36318
rect 5742 36370 5794 36382
rect 11566 36370 11618 36382
rect 6290 36318 6302 36370
rect 6354 36318 6366 36370
rect 6850 36318 6862 36370
rect 6914 36318 6926 36370
rect 8754 36318 8766 36370
rect 8818 36318 8830 36370
rect 9090 36318 9102 36370
rect 9154 36318 9166 36370
rect 5742 36306 5794 36318
rect 11566 36306 11618 36318
rect 11902 36370 11954 36382
rect 18958 36370 19010 36382
rect 23102 36370 23154 36382
rect 14242 36318 14254 36370
rect 14306 36318 14318 36370
rect 18498 36318 18510 36370
rect 18562 36318 18574 36370
rect 19618 36318 19630 36370
rect 19682 36318 19694 36370
rect 21410 36318 21422 36370
rect 21474 36318 21486 36370
rect 11902 36306 11954 36318
rect 18958 36306 19010 36318
rect 23102 36306 23154 36318
rect 23774 36370 23826 36382
rect 23774 36306 23826 36318
rect 24782 36370 24834 36382
rect 24782 36306 24834 36318
rect 26574 36370 26626 36382
rect 26574 36306 26626 36318
rect 27918 36370 27970 36382
rect 27918 36306 27970 36318
rect 29374 36370 29426 36382
rect 29374 36306 29426 36318
rect 29934 36370 29986 36382
rect 29934 36306 29986 36318
rect 30046 36370 30098 36382
rect 30046 36306 30098 36318
rect 32174 36370 32226 36382
rect 34078 36370 34130 36382
rect 33730 36318 33742 36370
rect 33794 36318 33806 36370
rect 43698 36318 43710 36370
rect 43762 36318 43774 36370
rect 44146 36318 44158 36370
rect 44210 36318 44222 36370
rect 32174 36306 32226 36318
rect 34078 36306 34130 36318
rect 10110 36258 10162 36270
rect 10110 36194 10162 36206
rect 10558 36258 10610 36270
rect 10558 36194 10610 36206
rect 11006 36258 11058 36270
rect 11006 36194 11058 36206
rect 11230 36258 11282 36270
rect 11230 36194 11282 36206
rect 13694 36258 13746 36270
rect 18846 36258 18898 36270
rect 15026 36206 15038 36258
rect 15090 36206 15102 36258
rect 13694 36194 13746 36206
rect 18846 36194 18898 36206
rect 19518 36258 19570 36270
rect 19518 36194 19570 36206
rect 20862 36258 20914 36270
rect 20862 36194 20914 36206
rect 22654 36258 22706 36270
rect 22654 36194 22706 36206
rect 23886 36258 23938 36270
rect 23886 36194 23938 36206
rect 24222 36258 24274 36270
rect 24222 36194 24274 36206
rect 24558 36258 24610 36270
rect 24558 36194 24610 36206
rect 25454 36258 25506 36270
rect 25454 36194 25506 36206
rect 26350 36258 26402 36270
rect 26350 36194 26402 36206
rect 27022 36258 27074 36270
rect 27022 36194 27074 36206
rect 28590 36258 28642 36270
rect 28590 36194 28642 36206
rect 29822 36258 29874 36270
rect 29822 36194 29874 36206
rect 31166 36258 31218 36270
rect 31166 36194 31218 36206
rect 31614 36258 31666 36270
rect 35086 36258 35138 36270
rect 32722 36206 32734 36258
rect 32786 36206 32798 36258
rect 31614 36194 31666 36206
rect 35086 36194 35138 36206
rect 40574 36258 40626 36270
rect 40574 36194 40626 36206
rect 44942 36258 44994 36270
rect 44942 36194 44994 36206
rect 1344 36090 48720 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48720 36090
rect 1344 36004 48720 36038
rect 10782 35922 10834 35934
rect 14590 35922 14642 35934
rect 8530 35870 8542 35922
rect 8594 35870 8606 35922
rect 14242 35870 14254 35922
rect 14306 35870 14318 35922
rect 10782 35858 10834 35870
rect 14590 35858 14642 35870
rect 15374 35922 15426 35934
rect 15374 35858 15426 35870
rect 15822 35922 15874 35934
rect 15822 35858 15874 35870
rect 16158 35922 16210 35934
rect 16158 35858 16210 35870
rect 16270 35922 16322 35934
rect 16270 35858 16322 35870
rect 16382 35922 16434 35934
rect 23102 35922 23154 35934
rect 21634 35870 21646 35922
rect 21698 35870 21710 35922
rect 16382 35858 16434 35870
rect 23102 35858 23154 35870
rect 28142 35922 28194 35934
rect 28142 35858 28194 35870
rect 29486 35922 29538 35934
rect 29486 35858 29538 35870
rect 30942 35922 30994 35934
rect 30942 35858 30994 35870
rect 32286 35922 32338 35934
rect 32286 35858 32338 35870
rect 43262 35922 43314 35934
rect 43262 35858 43314 35870
rect 16606 35810 16658 35822
rect 9650 35758 9662 35810
rect 9714 35758 9726 35810
rect 10210 35758 10222 35810
rect 10274 35758 10286 35810
rect 16606 35746 16658 35758
rect 22206 35810 22258 35822
rect 22206 35746 22258 35758
rect 22542 35810 22594 35822
rect 22542 35746 22594 35758
rect 22990 35810 23042 35822
rect 22990 35746 23042 35758
rect 24110 35810 24162 35822
rect 24110 35746 24162 35758
rect 26462 35810 26514 35822
rect 26462 35746 26514 35758
rect 27806 35810 27858 35822
rect 27806 35746 27858 35758
rect 28366 35810 28418 35822
rect 28366 35746 28418 35758
rect 29038 35810 29090 35822
rect 29038 35746 29090 35758
rect 29934 35810 29986 35822
rect 29934 35746 29986 35758
rect 31950 35810 32002 35822
rect 31950 35746 32002 35758
rect 32510 35810 32562 35822
rect 32510 35746 32562 35758
rect 33854 35810 33906 35822
rect 42690 35758 42702 35810
rect 42754 35758 42766 35810
rect 33854 35746 33906 35758
rect 21982 35698 22034 35710
rect 28142 35698 28194 35710
rect 5618 35646 5630 35698
rect 5682 35646 5694 35698
rect 6178 35646 6190 35698
rect 6242 35646 6254 35698
rect 13906 35646 13918 35698
rect 13970 35646 13982 35698
rect 18722 35646 18734 35698
rect 18786 35646 18798 35698
rect 22754 35646 22766 35698
rect 22818 35646 22830 35698
rect 23650 35646 23662 35698
rect 23714 35646 23726 35698
rect 21982 35634 22034 35646
rect 28142 35634 28194 35646
rect 29262 35698 29314 35710
rect 29262 35634 29314 35646
rect 29598 35698 29650 35710
rect 29598 35634 29650 35646
rect 30158 35698 30210 35710
rect 30158 35634 30210 35646
rect 30494 35698 30546 35710
rect 30494 35634 30546 35646
rect 32286 35698 32338 35710
rect 32286 35634 32338 35646
rect 33630 35698 33682 35710
rect 41918 35698 41970 35710
rect 34514 35646 34526 35698
rect 34578 35646 34590 35698
rect 35074 35646 35086 35698
rect 35138 35646 35150 35698
rect 39778 35646 39790 35698
rect 39842 35646 39854 35698
rect 42354 35646 42366 35698
rect 42418 35646 42430 35698
rect 33630 35634 33682 35646
rect 41918 35634 41970 35646
rect 10446 35586 10498 35598
rect 18174 35586 18226 35598
rect 25678 35586 25730 35598
rect 12674 35534 12686 35586
rect 12738 35534 12750 35586
rect 20178 35534 20190 35586
rect 20242 35534 20254 35586
rect 23538 35534 23550 35586
rect 23602 35534 23614 35586
rect 10446 35522 10498 35534
rect 18174 35522 18226 35534
rect 25678 35522 25730 35534
rect 26126 35586 26178 35598
rect 26126 35522 26178 35534
rect 26686 35586 26738 35598
rect 26686 35522 26738 35534
rect 27470 35586 27522 35598
rect 27470 35522 27522 35534
rect 30046 35586 30098 35598
rect 30046 35522 30098 35534
rect 31390 35586 31442 35598
rect 41246 35586 41298 35598
rect 37426 35534 37438 35586
rect 37490 35534 37502 35586
rect 39218 35534 39230 35586
rect 39282 35534 39294 35586
rect 31390 35522 31442 35534
rect 41246 35522 41298 35534
rect 23326 35474 23378 35486
rect 23326 35410 23378 35422
rect 27022 35474 27074 35486
rect 33294 35474 33346 35486
rect 30818 35422 30830 35474
rect 30882 35471 30894 35474
rect 31602 35471 31614 35474
rect 30882 35425 31614 35471
rect 30882 35422 30894 35425
rect 31602 35422 31614 35425
rect 31666 35422 31678 35474
rect 27022 35410 27074 35422
rect 33294 35410 33346 35422
rect 41582 35474 41634 35486
rect 41582 35410 41634 35422
rect 1344 35306 48720 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48720 35306
rect 1344 35220 48720 35254
rect 20190 35138 20242 35150
rect 18834 35086 18846 35138
rect 18898 35086 18910 35138
rect 20190 35074 20242 35086
rect 35198 35138 35250 35150
rect 35198 35074 35250 35086
rect 10334 35026 10386 35038
rect 10334 34962 10386 34974
rect 10558 35026 10610 35038
rect 10558 34962 10610 34974
rect 11118 35026 11170 35038
rect 14254 35026 14306 35038
rect 12226 34974 12238 35026
rect 12290 34974 12302 35026
rect 11118 34962 11170 34974
rect 14254 34962 14306 34974
rect 21646 35026 21698 35038
rect 34526 35026 34578 35038
rect 26226 34974 26238 35026
rect 26290 34974 26302 35026
rect 32610 34974 32622 35026
rect 32674 34974 32686 35026
rect 21646 34962 21698 34974
rect 34526 34962 34578 34974
rect 42142 35026 42194 35038
rect 42142 34962 42194 34974
rect 8318 34914 8370 34926
rect 1810 34862 1822 34914
rect 1874 34862 1886 34914
rect 2370 34862 2382 34914
rect 2434 34862 2446 34914
rect 4722 34862 4734 34914
rect 4786 34862 4798 34914
rect 8318 34850 8370 34862
rect 10782 34914 10834 34926
rect 10782 34850 10834 34862
rect 13806 34914 13858 34926
rect 13806 34850 13858 34862
rect 16606 34914 16658 34926
rect 16606 34850 16658 34862
rect 16942 34914 16994 34926
rect 16942 34850 16994 34862
rect 18062 34914 18114 34926
rect 18062 34850 18114 34862
rect 18286 34914 18338 34926
rect 18286 34850 18338 34862
rect 18622 34914 18674 34926
rect 19742 34914 19794 34926
rect 18946 34862 18958 34914
rect 19010 34862 19022 34914
rect 18622 34850 18674 34862
rect 19742 34850 19794 34862
rect 20078 34914 20130 34926
rect 22878 34914 22930 34926
rect 20514 34862 20526 34914
rect 20578 34862 20590 34914
rect 20078 34850 20130 34862
rect 22878 34850 22930 34862
rect 25006 34914 25058 34926
rect 25006 34850 25058 34862
rect 25118 34914 25170 34926
rect 27470 34914 27522 34926
rect 28142 34914 28194 34926
rect 26674 34862 26686 34914
rect 26738 34862 26750 34914
rect 27010 34862 27022 34914
rect 27074 34862 27086 34914
rect 25118 34850 25170 34862
rect 27246 34858 27298 34870
rect 6414 34802 6466 34814
rect 6414 34738 6466 34750
rect 6750 34802 6802 34814
rect 6750 34738 6802 34750
rect 7982 34802 8034 34814
rect 11678 34802 11730 34814
rect 8530 34750 8542 34802
rect 8594 34750 8606 34802
rect 8866 34750 8878 34802
rect 8930 34750 8942 34802
rect 7982 34738 8034 34750
rect 11678 34738 11730 34750
rect 11790 34802 11842 34814
rect 12574 34802 12626 34814
rect 12002 34750 12014 34802
rect 12066 34750 12078 34802
rect 11790 34738 11842 34750
rect 12574 34738 12626 34750
rect 12910 34802 12962 34814
rect 22318 34802 22370 34814
rect 14578 34750 14590 34802
rect 14642 34750 14654 34802
rect 12910 34738 12962 34750
rect 22318 34738 22370 34750
rect 25454 34802 25506 34814
rect 28018 34862 28030 34914
rect 28082 34862 28094 34914
rect 27470 34850 27522 34862
rect 28142 34850 28194 34862
rect 28254 34914 28306 34926
rect 28254 34850 28306 34862
rect 28590 34914 28642 34926
rect 35534 34914 35586 34926
rect 29698 34862 29710 34914
rect 29762 34862 29774 34914
rect 30482 34862 30494 34914
rect 30546 34862 30558 34914
rect 31042 34862 31054 34914
rect 31106 34862 31118 34914
rect 31490 34862 31502 34914
rect 31554 34862 31566 34914
rect 36194 34862 36206 34914
rect 36258 34862 36270 34914
rect 37650 34862 37662 34914
rect 37714 34862 37726 34914
rect 38210 34862 38222 34914
rect 38274 34862 38286 34914
rect 40562 34862 40574 34914
rect 40626 34862 40638 34914
rect 41234 34862 41246 34914
rect 41298 34862 41310 34914
rect 28590 34850 28642 34862
rect 35534 34850 35586 34862
rect 27246 34794 27298 34806
rect 27358 34802 27410 34814
rect 37102 34802 37154 34814
rect 25454 34738 25506 34750
rect 29810 34750 29822 34802
rect 29874 34750 29886 34802
rect 36082 34750 36094 34802
rect 36146 34750 36158 34802
rect 27358 34738 27410 34750
rect 37102 34738 37154 34750
rect 43038 34802 43090 34814
rect 43038 34738 43090 34750
rect 43374 34802 43426 34814
rect 43374 34738 43426 34750
rect 46510 34802 46562 34814
rect 46510 34738 46562 34750
rect 9662 34690 9714 34702
rect 9662 34626 9714 34638
rect 11454 34690 11506 34702
rect 14926 34690 14978 34702
rect 13458 34638 13470 34690
rect 13522 34638 13534 34690
rect 11454 34626 11506 34638
rect 14926 34626 14978 34638
rect 15374 34690 15426 34702
rect 15374 34626 15426 34638
rect 16830 34690 16882 34702
rect 16830 34626 16882 34638
rect 19070 34690 19122 34702
rect 19070 34626 19122 34638
rect 20526 34690 20578 34702
rect 20526 34626 20578 34638
rect 21982 34690 22034 34702
rect 21982 34626 22034 34638
rect 23214 34690 23266 34702
rect 23214 34626 23266 34638
rect 24558 34690 24610 34702
rect 24558 34626 24610 34638
rect 25342 34690 25394 34702
rect 25342 34626 25394 34638
rect 25790 34690 25842 34702
rect 25790 34626 25842 34638
rect 27806 34690 27858 34702
rect 27806 34626 27858 34638
rect 29262 34690 29314 34702
rect 29262 34626 29314 34638
rect 31054 34690 31106 34702
rect 31054 34626 31106 34638
rect 37886 34690 37938 34702
rect 37886 34626 37938 34638
rect 41582 34690 41634 34702
rect 41582 34626 41634 34638
rect 42478 34690 42530 34702
rect 42478 34626 42530 34638
rect 43710 34690 43762 34702
rect 43710 34626 43762 34638
rect 44158 34690 44210 34702
rect 44158 34626 44210 34638
rect 46174 34690 46226 34702
rect 46174 34626 46226 34638
rect 1344 34522 48720 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48720 34522
rect 1344 34436 48720 34470
rect 2382 34354 2434 34366
rect 2382 34290 2434 34302
rect 10446 34354 10498 34366
rect 10446 34290 10498 34302
rect 17390 34354 17442 34366
rect 19518 34354 19570 34366
rect 18050 34302 18062 34354
rect 18114 34302 18126 34354
rect 17390 34290 17442 34302
rect 19518 34290 19570 34302
rect 20638 34354 20690 34366
rect 20638 34290 20690 34302
rect 21086 34354 21138 34366
rect 21086 34290 21138 34302
rect 31614 34354 31666 34366
rect 31614 34290 31666 34302
rect 33854 34354 33906 34366
rect 33854 34290 33906 34302
rect 34190 34354 34242 34366
rect 34190 34290 34242 34302
rect 35086 34354 35138 34366
rect 35086 34290 35138 34302
rect 37998 34354 38050 34366
rect 37998 34290 38050 34302
rect 39678 34354 39730 34366
rect 39678 34290 39730 34302
rect 41022 34354 41074 34366
rect 41022 34290 41074 34302
rect 46622 34354 46674 34366
rect 46622 34290 46674 34302
rect 5742 34242 5794 34254
rect 5058 34190 5070 34242
rect 5122 34190 5134 34242
rect 5742 34178 5794 34190
rect 17726 34242 17778 34254
rect 27582 34242 27634 34254
rect 25554 34190 25566 34242
rect 25618 34190 25630 34242
rect 26226 34190 26238 34242
rect 26290 34190 26302 34242
rect 17726 34178 17778 34190
rect 27582 34178 27634 34190
rect 28590 34242 28642 34254
rect 31950 34242 32002 34254
rect 33630 34242 33682 34254
rect 30930 34190 30942 34242
rect 30994 34190 31006 34242
rect 33282 34190 33294 34242
rect 33346 34190 33358 34242
rect 34514 34190 34526 34242
rect 34578 34190 34590 34242
rect 35858 34190 35870 34242
rect 35922 34190 35934 34242
rect 36194 34190 36206 34242
rect 36258 34190 36270 34242
rect 38658 34190 38670 34242
rect 38722 34190 38734 34242
rect 38882 34190 38894 34242
rect 38946 34190 38958 34242
rect 42130 34190 42142 34242
rect 42194 34190 42206 34242
rect 42690 34190 42702 34242
rect 42754 34190 42766 34242
rect 46162 34190 46174 34242
rect 46226 34190 46238 34242
rect 47170 34190 47182 34242
rect 47234 34190 47246 34242
rect 47506 34190 47518 34242
rect 47570 34190 47582 34242
rect 28590 34178 28642 34190
rect 31950 34178 32002 34190
rect 33630 34178 33682 34190
rect 2718 34130 2770 34142
rect 2718 34066 2770 34078
rect 4174 34130 4226 34142
rect 4174 34066 4226 34078
rect 4510 34130 4562 34142
rect 18398 34130 18450 34142
rect 5282 34078 5294 34130
rect 5346 34078 5358 34130
rect 6178 34078 6190 34130
rect 6242 34078 6254 34130
rect 13346 34078 13358 34130
rect 13410 34078 13422 34130
rect 13906 34078 13918 34130
rect 13970 34078 13982 34130
rect 14466 34078 14478 34130
rect 14530 34078 14542 34130
rect 16818 34078 16830 34130
rect 16882 34078 16894 34130
rect 4510 34066 4562 34078
rect 18398 34066 18450 34078
rect 18734 34130 18786 34142
rect 19182 34130 19234 34142
rect 27470 34130 27522 34142
rect 18946 34078 18958 34130
rect 19010 34078 19022 34130
rect 19394 34078 19406 34130
rect 19458 34078 19470 34130
rect 21298 34078 21310 34130
rect 21362 34078 21374 34130
rect 21970 34078 21982 34130
rect 22034 34078 22046 34130
rect 25442 34078 25454 34130
rect 25506 34078 25518 34130
rect 26674 34078 26686 34130
rect 26738 34078 26750 34130
rect 18734 34066 18786 34078
rect 19182 34066 19234 34078
rect 27470 34066 27522 34078
rect 28030 34130 28082 34142
rect 28030 34066 28082 34078
rect 28926 34130 28978 34142
rect 28926 34066 28978 34078
rect 29038 34130 29090 34142
rect 29038 34066 29090 34078
rect 29262 34130 29314 34142
rect 32286 34130 32338 34142
rect 29810 34078 29822 34130
rect 29874 34078 29886 34130
rect 31042 34078 31054 34130
rect 31106 34078 31118 34130
rect 29262 34066 29314 34078
rect 32286 34066 32338 34078
rect 32510 34130 32562 34142
rect 38334 34130 38386 34142
rect 46958 34130 47010 34142
rect 33394 34078 33406 34130
rect 33458 34078 33470 34130
rect 43250 34078 43262 34130
rect 43314 34078 43326 34130
rect 43698 34078 43710 34130
rect 43762 34078 43774 34130
rect 32510 34066 32562 34078
rect 38334 34066 38386 34078
rect 46958 34066 47010 34078
rect 6750 34018 6802 34030
rect 6750 33954 6802 33966
rect 9886 34018 9938 34030
rect 19966 34018 20018 34030
rect 26238 34018 26290 34030
rect 11106 33966 11118 34018
rect 11170 33966 11182 34018
rect 24434 33966 24446 34018
rect 24498 33966 24510 34018
rect 9886 33954 9938 33966
rect 19966 33954 20018 33966
rect 26238 33954 26290 33966
rect 27806 34018 27858 34030
rect 27806 33954 27858 33966
rect 30270 34018 30322 34030
rect 30270 33954 30322 33966
rect 30382 34018 30434 34030
rect 30382 33954 30434 33966
rect 32062 34018 32114 34030
rect 33506 33966 33518 34018
rect 33570 33966 33582 34018
rect 32062 33954 32114 33966
rect 36430 33906 36482 33918
rect 36430 33842 36482 33854
rect 36766 33906 36818 33918
rect 36766 33842 36818 33854
rect 41582 33906 41634 33918
rect 41582 33842 41634 33854
rect 41918 33906 41970 33918
rect 41918 33842 41970 33854
rect 1344 33738 48720 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48720 33738
rect 1344 33652 48720 33686
rect 3838 33570 3890 33582
rect 3838 33506 3890 33518
rect 16382 33570 16434 33582
rect 22542 33570 22594 33582
rect 17154 33518 17166 33570
rect 17218 33567 17230 33570
rect 18050 33567 18062 33570
rect 17218 33521 18062 33567
rect 17218 33518 17230 33521
rect 18050 33518 18062 33521
rect 18114 33518 18126 33570
rect 18274 33518 18286 33570
rect 18338 33567 18350 33570
rect 18722 33567 18734 33570
rect 18338 33521 18734 33567
rect 18338 33518 18350 33521
rect 18722 33518 18734 33521
rect 18786 33518 18798 33570
rect 16382 33506 16434 33518
rect 22542 33506 22594 33518
rect 24558 33570 24610 33582
rect 24558 33506 24610 33518
rect 25006 33570 25058 33582
rect 25006 33506 25058 33518
rect 34750 33570 34802 33582
rect 34750 33506 34802 33518
rect 43038 33570 43090 33582
rect 43038 33506 43090 33518
rect 15598 33458 15650 33470
rect 8978 33406 8990 33458
rect 9042 33406 9054 33458
rect 15598 33394 15650 33406
rect 17166 33458 17218 33470
rect 17166 33394 17218 33406
rect 17726 33458 17778 33470
rect 17726 33394 17778 33406
rect 19406 33458 19458 33470
rect 19406 33394 19458 33406
rect 24334 33458 24386 33470
rect 24334 33394 24386 33406
rect 29374 33458 29426 33470
rect 29374 33394 29426 33406
rect 33966 33458 34018 33470
rect 38546 33406 38558 33458
rect 38610 33406 38622 33458
rect 41234 33406 41246 33458
rect 41298 33406 41310 33458
rect 33966 33394 34018 33406
rect 10334 33346 10386 33358
rect 4386 33294 4398 33346
rect 4450 33294 4462 33346
rect 6066 33294 6078 33346
rect 6130 33294 6142 33346
rect 6626 33294 6638 33346
rect 6690 33294 6702 33346
rect 10334 33282 10386 33294
rect 15822 33346 15874 33358
rect 19518 33346 19570 33358
rect 16706 33294 16718 33346
rect 16770 33294 16782 33346
rect 15822 33282 15874 33294
rect 19518 33282 19570 33294
rect 19966 33346 20018 33358
rect 19966 33282 20018 33294
rect 22878 33346 22930 33358
rect 22878 33282 22930 33294
rect 24110 33346 24162 33358
rect 24110 33282 24162 33294
rect 25342 33346 25394 33358
rect 25342 33282 25394 33294
rect 28702 33346 28754 33358
rect 32734 33346 32786 33358
rect 29922 33294 29934 33346
rect 29986 33294 29998 33346
rect 30930 33294 30942 33346
rect 30994 33294 31006 33346
rect 28702 33282 28754 33294
rect 32734 33282 32786 33294
rect 33294 33346 33346 33358
rect 33294 33282 33346 33294
rect 35086 33346 35138 33358
rect 35086 33282 35138 33294
rect 36990 33346 37042 33358
rect 42142 33346 42194 33358
rect 38210 33294 38222 33346
rect 38274 33294 38286 33346
rect 39554 33294 39566 33346
rect 39618 33294 39630 33346
rect 36990 33282 37042 33294
rect 42142 33282 42194 33294
rect 42590 33346 42642 33358
rect 42590 33282 42642 33294
rect 43374 33346 43426 33358
rect 43810 33294 43822 33346
rect 43874 33294 43886 33346
rect 45266 33294 45278 33346
rect 45330 33294 45342 33346
rect 45938 33294 45950 33346
rect 46002 33294 46014 33346
rect 43374 33282 43426 33294
rect 10222 33234 10274 33246
rect 4610 33182 4622 33234
rect 4674 33182 4686 33234
rect 10222 33170 10274 33182
rect 10670 33234 10722 33246
rect 15486 33234 15538 33246
rect 12114 33182 12126 33234
rect 12178 33182 12190 33234
rect 13794 33182 13806 33234
rect 13858 33182 13870 33234
rect 10670 33170 10722 33182
rect 15486 33170 15538 33182
rect 16046 33234 16098 33246
rect 16046 33170 16098 33182
rect 16494 33234 16546 33246
rect 27134 33234 27186 33246
rect 23202 33182 23214 33234
rect 23266 33182 23278 33234
rect 23650 33182 23662 33234
rect 23714 33182 23726 33234
rect 16494 33170 16546 33182
rect 27134 33170 27186 33182
rect 28366 33234 28418 33246
rect 28366 33170 28418 33182
rect 28478 33234 28530 33246
rect 32846 33234 32898 33246
rect 41918 33234 41970 33246
rect 29698 33182 29710 33234
rect 29762 33182 29774 33234
rect 30706 33182 30718 33234
rect 30770 33182 30782 33234
rect 35298 33182 35310 33234
rect 35362 33182 35374 33234
rect 35858 33182 35870 33234
rect 35922 33182 35934 33234
rect 43922 33182 43934 33234
rect 43986 33182 43998 33234
rect 28478 33170 28530 33182
rect 32846 33170 32898 33182
rect 41918 33170 41970 33182
rect 3502 33122 3554 33134
rect 3502 33058 3554 33070
rect 10894 33122 10946 33134
rect 10894 33058 10946 33070
rect 11006 33122 11058 33134
rect 11006 33058 11058 33070
rect 11790 33122 11842 33134
rect 11790 33058 11842 33070
rect 12462 33122 12514 33134
rect 12462 33058 12514 33070
rect 12910 33122 12962 33134
rect 12910 33058 12962 33070
rect 13470 33122 13522 33134
rect 13470 33058 13522 33070
rect 14366 33122 14418 33134
rect 14366 33058 14418 33070
rect 18174 33122 18226 33134
rect 18174 33058 18226 33070
rect 18622 33122 18674 33134
rect 18622 33058 18674 33070
rect 19294 33122 19346 33134
rect 19294 33058 19346 33070
rect 20414 33122 20466 33134
rect 20414 33058 20466 33070
rect 20862 33122 20914 33134
rect 20862 33058 20914 33070
rect 26798 33122 26850 33134
rect 26798 33058 26850 33070
rect 27582 33122 27634 33134
rect 27582 33058 27634 33070
rect 28142 33122 28194 33134
rect 28142 33058 28194 33070
rect 31502 33122 31554 33134
rect 31502 33058 31554 33070
rect 32398 33122 32450 33134
rect 32398 33058 32450 33070
rect 32958 33122 33010 33134
rect 32958 33058 33010 33070
rect 37326 33122 37378 33134
rect 37326 33058 37378 33070
rect 37774 33122 37826 33134
rect 37774 33058 37826 33070
rect 42254 33122 42306 33134
rect 48290 33070 48302 33122
rect 48354 33070 48366 33122
rect 42254 33058 42306 33070
rect 1344 32954 48720 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48720 32954
rect 1344 32868 48720 32902
rect 6974 32786 7026 32798
rect 4722 32734 4734 32786
rect 4786 32734 4798 32786
rect 6974 32722 7026 32734
rect 9662 32786 9714 32798
rect 9662 32722 9714 32734
rect 11006 32786 11058 32798
rect 11006 32722 11058 32734
rect 11230 32786 11282 32798
rect 11230 32722 11282 32734
rect 12126 32786 12178 32798
rect 12126 32722 12178 32734
rect 12574 32786 12626 32798
rect 12574 32722 12626 32734
rect 14254 32786 14306 32798
rect 14254 32722 14306 32734
rect 15150 32786 15202 32798
rect 39342 32786 39394 32798
rect 29138 32734 29150 32786
rect 29202 32734 29214 32786
rect 30594 32734 30606 32786
rect 30658 32734 30670 32786
rect 35410 32734 35422 32786
rect 35474 32734 35486 32786
rect 15150 32722 15202 32734
rect 39342 32722 39394 32734
rect 43038 32786 43090 32798
rect 43038 32722 43090 32734
rect 9998 32674 10050 32686
rect 8642 32622 8654 32674
rect 8706 32622 8718 32674
rect 9998 32610 10050 32622
rect 10110 32674 10162 32686
rect 10110 32610 10162 32622
rect 12910 32674 12962 32686
rect 12910 32610 12962 32622
rect 13806 32674 13858 32686
rect 20526 32674 20578 32686
rect 15474 32622 15486 32674
rect 15538 32622 15550 32674
rect 13806 32610 13858 32622
rect 20526 32610 20578 32622
rect 29934 32674 29986 32686
rect 29934 32610 29986 32622
rect 31614 32674 31666 32686
rect 31614 32610 31666 32622
rect 31950 32674 32002 32686
rect 33742 32674 33794 32686
rect 33394 32622 33406 32674
rect 33458 32622 33470 32674
rect 31950 32610 32002 32622
rect 33742 32610 33794 32622
rect 46286 32674 46338 32686
rect 46286 32610 46338 32622
rect 5742 32562 5794 32574
rect 1810 32510 1822 32562
rect 1874 32510 1886 32562
rect 2258 32510 2270 32562
rect 2322 32510 2334 32562
rect 5742 32498 5794 32510
rect 7310 32562 7362 32574
rect 7310 32498 7362 32510
rect 7758 32562 7810 32574
rect 7758 32498 7810 32510
rect 8094 32562 8146 32574
rect 10334 32562 10386 32574
rect 8754 32510 8766 32562
rect 8818 32510 8830 32562
rect 8094 32498 8146 32510
rect 10334 32498 10386 32510
rect 10782 32562 10834 32574
rect 10782 32498 10834 32510
rect 11454 32562 11506 32574
rect 11454 32498 11506 32510
rect 11566 32562 11618 32574
rect 11566 32498 11618 32510
rect 12238 32562 12290 32574
rect 12238 32498 12290 32510
rect 12574 32562 12626 32574
rect 12574 32498 12626 32510
rect 13134 32562 13186 32574
rect 13134 32498 13186 32510
rect 13470 32562 13522 32574
rect 13470 32498 13522 32510
rect 17950 32562 18002 32574
rect 17950 32498 18002 32510
rect 20862 32562 20914 32574
rect 30942 32562 30994 32574
rect 33966 32562 34018 32574
rect 39790 32562 39842 32574
rect 26226 32510 26238 32562
rect 26290 32510 26302 32562
rect 26786 32510 26798 32562
rect 26850 32510 26862 32562
rect 30146 32510 30158 32562
rect 30210 32510 30222 32562
rect 33506 32510 33518 32562
rect 33570 32510 33582 32562
rect 37762 32510 37774 32562
rect 37826 32510 37838 32562
rect 38546 32510 38558 32562
rect 38610 32510 38622 32562
rect 20862 32498 20914 32510
rect 30942 32498 30994 32510
rect 33966 32498 34018 32510
rect 39790 32498 39842 32510
rect 40910 32562 40962 32574
rect 46622 32562 46674 32574
rect 41234 32510 41246 32562
rect 41298 32510 41310 32562
rect 42130 32510 42142 32562
rect 42194 32510 42206 32562
rect 40910 32498 40962 32510
rect 46622 32498 46674 32510
rect 5182 32450 5234 32462
rect 5182 32386 5234 32398
rect 6190 32450 6242 32462
rect 6190 32386 6242 32398
rect 13358 32450 13410 32462
rect 13358 32386 13410 32398
rect 17390 32450 17442 32462
rect 17390 32386 17442 32398
rect 18398 32450 18450 32462
rect 18398 32386 18450 32398
rect 18846 32450 18898 32462
rect 18846 32386 18898 32398
rect 19742 32450 19794 32462
rect 19742 32386 19794 32398
rect 20302 32450 20354 32462
rect 20302 32386 20354 32398
rect 21310 32450 21362 32462
rect 21310 32386 21362 32398
rect 29598 32450 29650 32462
rect 29598 32386 29650 32398
rect 32510 32450 32562 32462
rect 39566 32450 39618 32462
rect 33618 32398 33630 32450
rect 33682 32398 33694 32450
rect 32510 32386 32562 32398
rect 39566 32386 39618 32398
rect 40126 32450 40178 32462
rect 41122 32398 41134 32450
rect 41186 32398 41198 32450
rect 42466 32398 42478 32450
rect 42530 32398 42542 32450
rect 40126 32386 40178 32398
rect 5954 32286 5966 32338
rect 6018 32335 6030 32338
rect 6178 32335 6190 32338
rect 6018 32289 6190 32335
rect 6018 32286 6030 32289
rect 6178 32286 6190 32289
rect 6242 32286 6254 32338
rect 18162 32286 18174 32338
rect 18226 32335 18238 32338
rect 18386 32335 18398 32338
rect 18226 32289 18398 32335
rect 18226 32286 18238 32289
rect 18386 32286 18398 32289
rect 18450 32286 18462 32338
rect 19506 32286 19518 32338
rect 19570 32335 19582 32338
rect 19730 32335 19742 32338
rect 19570 32289 19742 32335
rect 19570 32286 19582 32289
rect 19730 32286 19742 32289
rect 19794 32335 19806 32338
rect 20066 32335 20078 32338
rect 19794 32289 20078 32335
rect 19794 32286 19806 32289
rect 20066 32286 20078 32289
rect 20130 32286 20142 32338
rect 1344 32170 48720 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48720 32170
rect 1344 32084 48720 32118
rect 3950 32002 4002 32014
rect 3950 31938 4002 31950
rect 21534 32002 21586 32014
rect 21534 31938 21586 31950
rect 33518 32002 33570 32014
rect 33518 31938 33570 31950
rect 11678 31890 11730 31902
rect 11678 31826 11730 31838
rect 18510 31890 18562 31902
rect 23662 31890 23714 31902
rect 18834 31838 18846 31890
rect 18898 31838 18910 31890
rect 18510 31826 18562 31838
rect 23662 31826 23714 31838
rect 32062 31890 32114 31902
rect 43038 31890 43090 31902
rect 40114 31838 40126 31890
rect 40178 31838 40190 31890
rect 32062 31826 32114 31838
rect 43038 31826 43090 31838
rect 2494 31778 2546 31790
rect 19630 31778 19682 31790
rect 21870 31778 21922 31790
rect 30270 31778 30322 31790
rect 4722 31726 4734 31778
rect 4786 31726 4798 31778
rect 15250 31726 15262 31778
rect 15314 31726 15326 31778
rect 15810 31726 15822 31778
rect 15874 31726 15886 31778
rect 19954 31726 19966 31778
rect 20018 31726 20030 31778
rect 22530 31726 22542 31778
rect 22594 31726 22606 31778
rect 26002 31726 26014 31778
rect 26066 31726 26078 31778
rect 27010 31726 27022 31778
rect 27074 31726 27086 31778
rect 27458 31726 27470 31778
rect 27522 31726 27534 31778
rect 2494 31714 2546 31726
rect 19630 31714 19682 31726
rect 21870 31714 21922 31726
rect 30270 31714 30322 31726
rect 31166 31778 31218 31790
rect 31166 31714 31218 31726
rect 32622 31778 32674 31790
rect 32622 31714 32674 31726
rect 32958 31778 33010 31790
rect 32958 31714 33010 31726
rect 33854 31778 33906 31790
rect 33854 31714 33906 31726
rect 34078 31778 34130 31790
rect 37202 31726 37214 31778
rect 37266 31726 37278 31778
rect 40562 31726 40574 31778
rect 40626 31726 40638 31778
rect 41010 31726 41022 31778
rect 41074 31726 41086 31778
rect 42242 31726 42254 31778
rect 42306 31726 42318 31778
rect 45266 31726 45278 31778
rect 45330 31726 45342 31778
rect 45938 31726 45950 31778
rect 46002 31726 46014 31778
rect 34078 31714 34130 31726
rect 2158 31666 2210 31678
rect 11566 31666 11618 31678
rect 4498 31614 4510 31666
rect 4562 31614 4574 31666
rect 2158 31602 2210 31614
rect 11566 31602 11618 31614
rect 11902 31666 11954 31678
rect 11902 31602 11954 31614
rect 12126 31666 12178 31678
rect 12126 31602 12178 31614
rect 18734 31666 18786 31678
rect 18734 31602 18786 31614
rect 20414 31666 20466 31678
rect 20414 31602 20466 31614
rect 20638 31666 20690 31678
rect 33182 31666 33234 31678
rect 43262 31666 43314 31678
rect 22642 31614 22654 31666
rect 22706 31614 22718 31666
rect 23874 31614 23886 31666
rect 23938 31614 23950 31666
rect 24210 31614 24222 31666
rect 24274 31614 24286 31666
rect 26114 31614 26126 31666
rect 26178 31614 26190 31666
rect 26674 31614 26686 31666
rect 26738 31614 26750 31666
rect 29922 31614 29934 31666
rect 29986 31614 29998 31666
rect 40450 31614 40462 31666
rect 40514 31614 40526 31666
rect 40898 31614 40910 31666
rect 40962 31614 40974 31666
rect 20638 31602 20690 31614
rect 33182 31602 33234 31614
rect 43262 31602 43314 31614
rect 43598 31666 43650 31678
rect 43598 31602 43650 31614
rect 3614 31554 3666 31566
rect 3614 31490 3666 31502
rect 12686 31554 12738 31566
rect 19406 31554 19458 31566
rect 18162 31502 18174 31554
rect 18226 31502 18238 31554
rect 12686 31490 12738 31502
rect 19406 31490 19458 31502
rect 19518 31554 19570 31566
rect 19518 31490 19570 31502
rect 20526 31554 20578 31566
rect 20526 31490 20578 31502
rect 23326 31554 23378 31566
rect 23326 31490 23378 31502
rect 25118 31554 25170 31566
rect 25118 31490 25170 31502
rect 25454 31554 25506 31566
rect 25454 31490 25506 31502
rect 27918 31554 27970 31566
rect 27918 31490 27970 31502
rect 30606 31554 30658 31566
rect 30606 31490 30658 31502
rect 31502 31554 31554 31566
rect 31502 31490 31554 31502
rect 32846 31554 32898 31566
rect 32846 31490 32898 31502
rect 34526 31554 34578 31566
rect 34526 31490 34578 31502
rect 35982 31554 36034 31566
rect 35982 31490 36034 31502
rect 37438 31554 37490 31566
rect 37438 31490 37490 31502
rect 39902 31554 39954 31566
rect 43934 31554 43986 31566
rect 42690 31502 42702 31554
rect 42754 31502 42766 31554
rect 48290 31502 48302 31554
rect 48354 31502 48366 31554
rect 39902 31490 39954 31502
rect 43934 31490 43986 31502
rect 1344 31386 48720 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48720 31386
rect 1344 31300 48720 31334
rect 5406 31218 5458 31230
rect 17502 31218 17554 31230
rect 24670 31218 24722 31230
rect 8866 31166 8878 31218
rect 8930 31166 8942 31218
rect 19058 31166 19070 31218
rect 19122 31166 19134 31218
rect 22754 31166 22766 31218
rect 22818 31166 22830 31218
rect 5406 31154 5458 31166
rect 17502 31154 17554 31166
rect 24670 31154 24722 31166
rect 26126 31218 26178 31230
rect 26126 31154 26178 31166
rect 27134 31218 27186 31230
rect 27134 31154 27186 31166
rect 30046 31218 30098 31230
rect 30046 31154 30098 31166
rect 30830 31218 30882 31230
rect 30830 31154 30882 31166
rect 31726 31218 31778 31230
rect 31726 31154 31778 31166
rect 35646 31218 35698 31230
rect 35646 31154 35698 31166
rect 41022 31218 41074 31230
rect 41022 31154 41074 31166
rect 41134 31218 41186 31230
rect 41134 31154 41186 31166
rect 46622 31218 46674 31230
rect 46622 31154 46674 31166
rect 48302 31218 48354 31230
rect 48302 31154 48354 31166
rect 2158 31106 2210 31118
rect 2158 31042 2210 31054
rect 2494 31106 2546 31118
rect 17390 31106 17442 31118
rect 4386 31054 4398 31106
rect 4450 31054 4462 31106
rect 4834 31054 4846 31106
rect 4898 31054 4910 31106
rect 14578 31054 14590 31106
rect 14642 31054 14654 31106
rect 2494 31042 2546 31054
rect 17390 31042 17442 31054
rect 17726 31106 17778 31118
rect 17726 31042 17778 31054
rect 17950 31106 18002 31118
rect 17950 31042 18002 31054
rect 23886 31106 23938 31118
rect 23886 31042 23938 31054
rect 26462 31106 26514 31118
rect 35086 31106 35138 31118
rect 28242 31054 28254 31106
rect 28306 31054 28318 31106
rect 26462 31042 26514 31054
rect 35086 31042 35138 31054
rect 40910 31106 40962 31118
rect 41458 31054 41470 31106
rect 41522 31054 41534 31106
rect 47170 31054 47182 31106
rect 47234 31054 47246 31106
rect 47506 31054 47518 31106
rect 47570 31054 47582 31106
rect 40910 31042 40962 31054
rect 5070 30994 5122 31006
rect 18622 30994 18674 31006
rect 5954 30942 5966 30994
rect 6018 30942 6030 30994
rect 6514 30942 6526 30994
rect 6578 30942 6590 30994
rect 9650 30942 9662 30994
rect 9714 30942 9726 30994
rect 10210 30942 10222 30994
rect 10274 30942 10286 30994
rect 14802 30942 14814 30994
rect 14866 30942 14878 30994
rect 5070 30930 5122 30942
rect 18622 30930 18674 30942
rect 18958 30994 19010 31006
rect 25230 30994 25282 31006
rect 19394 30942 19406 30994
rect 19458 30942 19470 30994
rect 19730 30942 19742 30994
rect 19794 30942 19806 30994
rect 20290 30942 20302 30994
rect 20354 30942 20366 30994
rect 24098 30942 24110 30994
rect 24162 30942 24174 30994
rect 24434 30942 24446 30994
rect 24498 30942 24510 30994
rect 18958 30930 19010 30942
rect 25230 30930 25282 30942
rect 25454 30994 25506 31006
rect 46958 30994 47010 31006
rect 28018 30942 28030 30994
rect 28082 30942 28094 30994
rect 30258 30942 30270 30994
rect 30322 30942 30334 30994
rect 38658 30942 38670 30994
rect 38722 30942 38734 30994
rect 39442 30942 39454 30994
rect 39506 30942 39518 30994
rect 41346 30942 41358 30994
rect 41410 30942 41422 30994
rect 44706 30942 44718 30994
rect 44770 30942 44782 30994
rect 45266 30942 45278 30994
rect 45330 30942 45342 30994
rect 25454 30930 25506 30942
rect 46958 30930 47010 30942
rect 15374 30882 15426 30894
rect 12562 30830 12574 30882
rect 12626 30830 12638 30882
rect 15374 30818 15426 30830
rect 23550 30882 23602 30894
rect 33182 30882 33234 30894
rect 40350 30882 40402 30894
rect 31266 30830 31278 30882
rect 31330 30830 31342 30882
rect 32162 30830 32174 30882
rect 32226 30830 32238 30882
rect 36306 30830 36318 30882
rect 36370 30830 36382 30882
rect 42354 30830 42366 30882
rect 42418 30830 42430 30882
rect 23550 30818 23602 30830
rect 33182 30818 33234 30830
rect 40350 30818 40402 30830
rect 13694 30770 13746 30782
rect 13694 30706 13746 30718
rect 14030 30770 14082 30782
rect 24334 30770 24386 30782
rect 19170 30718 19182 30770
rect 19234 30718 19246 30770
rect 14030 30706 14082 30718
rect 24334 30706 24386 30718
rect 25678 30770 25730 30782
rect 25678 30706 25730 30718
rect 27470 30770 27522 30782
rect 27470 30706 27522 30718
rect 1344 30602 48720 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48720 30602
rect 1344 30516 48720 30550
rect 12014 30434 12066 30446
rect 37774 30434 37826 30446
rect 20066 30382 20078 30434
rect 20130 30382 20142 30434
rect 22082 30382 22094 30434
rect 22146 30431 22158 30434
rect 22642 30431 22654 30434
rect 22146 30385 22654 30431
rect 22146 30382 22158 30385
rect 22642 30382 22654 30385
rect 22706 30382 22718 30434
rect 12014 30370 12066 30382
rect 37774 30370 37826 30382
rect 8430 30322 8482 30334
rect 8430 30258 8482 30270
rect 19630 30322 19682 30334
rect 40798 30322 40850 30334
rect 26562 30270 26574 30322
rect 26626 30270 26638 30322
rect 29922 30270 29934 30322
rect 29986 30270 29998 30322
rect 35074 30270 35086 30322
rect 35138 30270 35150 30322
rect 19630 30258 19682 30270
rect 40798 30258 40850 30270
rect 43374 30322 43426 30334
rect 47170 30270 47182 30322
rect 47234 30270 47246 30322
rect 43374 30258 43426 30270
rect 5742 30210 5794 30222
rect 1810 30158 1822 30210
rect 1874 30158 1886 30210
rect 2258 30158 2270 30210
rect 2322 30158 2334 30210
rect 5742 30146 5794 30158
rect 10670 30210 10722 30222
rect 10670 30146 10722 30158
rect 11678 30210 11730 30222
rect 11678 30146 11730 30158
rect 19854 30210 19906 30222
rect 30382 30210 30434 30222
rect 35534 30210 35586 30222
rect 20066 30158 20078 30210
rect 20130 30158 20142 30210
rect 23090 30158 23102 30210
rect 23154 30158 23166 30210
rect 26674 30158 26686 30210
rect 26738 30158 26750 30210
rect 27010 30158 27022 30210
rect 27074 30158 27086 30210
rect 32274 30158 32286 30210
rect 32338 30158 32350 30210
rect 19854 30146 19906 30158
rect 30382 30146 30434 30158
rect 35534 30146 35586 30158
rect 38110 30210 38162 30222
rect 38110 30146 38162 30158
rect 40686 30210 40738 30222
rect 40686 30146 40738 30158
rect 40910 30210 40962 30222
rect 40910 30146 40962 30158
rect 43038 30210 43090 30222
rect 44146 30158 44158 30210
rect 44210 30158 44222 30210
rect 46050 30158 46062 30210
rect 46114 30158 46126 30210
rect 43038 30146 43090 30158
rect 6862 30098 6914 30110
rect 6862 30034 6914 30046
rect 7198 30098 7250 30110
rect 7198 30034 7250 30046
rect 8094 30098 8146 30110
rect 10334 30098 10386 30110
rect 19518 30098 19570 30110
rect 41246 30098 41298 30110
rect 8754 30046 8766 30098
rect 8818 30046 8830 30098
rect 8978 30046 8990 30098
rect 9042 30046 9054 30098
rect 12226 30046 12238 30098
rect 12290 30046 12302 30098
rect 12562 30046 12574 30098
rect 12626 30046 12638 30098
rect 16034 30046 16046 30098
rect 16098 30046 16110 30098
rect 17714 30046 17726 30098
rect 17778 30046 17790 30098
rect 22866 30046 22878 30098
rect 22930 30046 22942 30098
rect 32946 30046 32958 30098
rect 33010 30046 33022 30098
rect 38434 30046 38446 30098
rect 38498 30046 38510 30098
rect 38658 30046 38670 30098
rect 38722 30046 38734 30098
rect 8094 30034 8146 30046
rect 10334 30034 10386 30046
rect 19518 30034 19570 30046
rect 41246 30034 41298 30046
rect 41582 30098 41634 30110
rect 41582 30034 41634 30046
rect 41918 30098 41970 30110
rect 43922 30046 43934 30098
rect 43986 30046 43998 30098
rect 41918 30034 41970 30046
rect 16382 29986 16434 29998
rect 4722 29934 4734 29986
rect 4786 29934 4798 29986
rect 16382 29922 16434 29934
rect 18062 29986 18114 29998
rect 18062 29922 18114 29934
rect 18510 29986 18562 29998
rect 18510 29922 18562 29934
rect 20862 29986 20914 29998
rect 20862 29922 20914 29934
rect 22430 29986 22482 29998
rect 22430 29922 22482 29934
rect 23662 29986 23714 29998
rect 23662 29922 23714 29934
rect 24894 29986 24946 29998
rect 24894 29922 24946 29934
rect 26238 29986 26290 29998
rect 26238 29922 26290 29934
rect 30942 29986 30994 29998
rect 30942 29922 30994 29934
rect 39454 29986 39506 29998
rect 39454 29922 39506 29934
rect 45614 29986 45666 29998
rect 45614 29922 45666 29934
rect 45838 29986 45890 29998
rect 45838 29922 45890 29934
rect 46734 29986 46786 29998
rect 46734 29922 46786 29934
rect 1344 29818 48720 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48720 29818
rect 1344 29732 48720 29766
rect 30270 29650 30322 29662
rect 23202 29598 23214 29650
rect 23266 29598 23278 29650
rect 24322 29598 24334 29650
rect 24386 29598 24398 29650
rect 28130 29598 28142 29650
rect 28194 29598 28206 29650
rect 36754 29598 36766 29650
rect 36818 29598 36830 29650
rect 44930 29598 44942 29650
rect 44994 29598 45006 29650
rect 30270 29586 30322 29598
rect 18622 29538 18674 29550
rect 13906 29486 13918 29538
rect 13970 29486 13982 29538
rect 14466 29486 14478 29538
rect 14530 29486 14542 29538
rect 18622 29474 18674 29486
rect 19182 29538 19234 29550
rect 19182 29474 19234 29486
rect 22542 29538 22594 29550
rect 22542 29474 22594 29486
rect 29374 29538 29426 29550
rect 29374 29474 29426 29486
rect 31838 29538 31890 29550
rect 31838 29474 31890 29486
rect 33182 29538 33234 29550
rect 39566 29538 39618 29550
rect 34514 29486 34526 29538
rect 34578 29486 34590 29538
rect 33182 29474 33234 29486
rect 39566 29474 39618 29486
rect 41246 29538 41298 29550
rect 41246 29474 41298 29486
rect 22878 29426 22930 29438
rect 24334 29426 24386 29438
rect 15698 29374 15710 29426
rect 15762 29374 15774 29426
rect 18162 29374 18174 29426
rect 18226 29374 18238 29426
rect 21746 29374 21758 29426
rect 21810 29374 21822 29426
rect 23426 29374 23438 29426
rect 23490 29374 23502 29426
rect 23874 29374 23886 29426
rect 23938 29374 23950 29426
rect 22878 29362 22930 29374
rect 24334 29362 24386 29374
rect 24670 29426 24722 29438
rect 26014 29426 26066 29438
rect 28814 29426 28866 29438
rect 25218 29374 25230 29426
rect 25282 29374 25294 29426
rect 28354 29374 28366 29426
rect 28418 29374 28430 29426
rect 24670 29362 24722 29374
rect 26014 29362 26066 29374
rect 28814 29362 28866 29374
rect 30606 29426 30658 29438
rect 34974 29426 35026 29438
rect 37102 29426 37154 29438
rect 31378 29374 31390 29426
rect 31442 29374 31454 29426
rect 34290 29374 34302 29426
rect 34354 29374 34366 29426
rect 35970 29374 35982 29426
rect 36034 29374 36046 29426
rect 30606 29362 30658 29374
rect 34974 29362 35026 29374
rect 37102 29362 37154 29374
rect 38670 29426 38722 29438
rect 38670 29362 38722 29374
rect 39790 29426 39842 29438
rect 41794 29374 41806 29426
rect 41858 29374 41870 29426
rect 42578 29374 42590 29426
rect 42642 29374 42654 29426
rect 45266 29374 45278 29426
rect 45330 29374 45342 29426
rect 45826 29374 45838 29426
rect 45890 29374 45902 29426
rect 48290 29374 48302 29426
rect 48354 29374 48366 29426
rect 39790 29362 39842 29374
rect 16158 29314 16210 29326
rect 32510 29314 32562 29326
rect 33406 29314 33458 29326
rect 17826 29262 17838 29314
rect 17890 29262 17902 29314
rect 22082 29262 22094 29314
rect 22146 29262 22158 29314
rect 33058 29262 33070 29314
rect 33122 29262 33134 29314
rect 16158 29250 16210 29262
rect 32510 29250 32562 29262
rect 33406 29250 33458 29262
rect 33966 29314 34018 29326
rect 33966 29250 34018 29262
rect 35534 29314 35586 29326
rect 35534 29250 35586 29262
rect 36430 29314 36482 29326
rect 36430 29250 36482 29262
rect 38334 29314 38386 29326
rect 38334 29250 38386 29262
rect 39230 29314 39282 29326
rect 39230 29250 39282 29262
rect 13358 29202 13410 29214
rect 13358 29138 13410 29150
rect 13694 29202 13746 29214
rect 13694 29138 13746 29150
rect 24222 29202 24274 29214
rect 24222 29138 24274 29150
rect 25230 29202 25282 29214
rect 25230 29138 25282 29150
rect 25566 29202 25618 29214
rect 25566 29138 25618 29150
rect 40126 29202 40178 29214
rect 40126 29138 40178 29150
rect 1344 29034 48720 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48720 29034
rect 1344 28948 48720 28982
rect 16606 28866 16658 28878
rect 16606 28802 16658 28814
rect 45950 28866 46002 28878
rect 45950 28802 46002 28814
rect 9886 28754 9938 28766
rect 9886 28690 9938 28702
rect 14254 28754 14306 28766
rect 14254 28690 14306 28702
rect 17390 28754 17442 28766
rect 30718 28754 30770 28766
rect 36094 28754 36146 28766
rect 20402 28702 20414 28754
rect 20466 28702 20478 28754
rect 27458 28702 27470 28754
rect 27522 28702 27534 28754
rect 34178 28702 34190 28754
rect 34242 28702 34254 28754
rect 17390 28690 17442 28702
rect 30718 28690 30770 28702
rect 36094 28690 36146 28702
rect 37438 28754 37490 28766
rect 37438 28690 37490 28702
rect 8206 28642 8258 28654
rect 1810 28590 1822 28642
rect 1874 28590 1886 28642
rect 2482 28590 2494 28642
rect 2546 28590 2558 28642
rect 4834 28590 4846 28642
rect 4898 28590 4910 28642
rect 8206 28578 8258 28590
rect 8318 28642 8370 28654
rect 8318 28578 8370 28590
rect 8766 28642 8818 28654
rect 8766 28578 8818 28590
rect 9774 28642 9826 28654
rect 9774 28578 9826 28590
rect 11006 28642 11058 28654
rect 11006 28578 11058 28590
rect 11902 28642 11954 28654
rect 14030 28642 14082 28654
rect 13570 28590 13582 28642
rect 13634 28590 13646 28642
rect 13794 28590 13806 28642
rect 13858 28590 13870 28642
rect 11902 28578 11954 28590
rect 14030 28578 14082 28590
rect 14926 28642 14978 28654
rect 19518 28642 19570 28654
rect 16930 28590 16942 28642
rect 16994 28590 17006 28642
rect 18386 28590 18398 28642
rect 18450 28590 18462 28642
rect 14926 28578 14978 28590
rect 19518 28578 19570 28590
rect 19742 28642 19794 28654
rect 19742 28578 19794 28590
rect 20078 28642 20130 28654
rect 23550 28642 23602 28654
rect 22418 28590 22430 28642
rect 22482 28590 22494 28642
rect 20078 28578 20130 28590
rect 23550 28578 23602 28590
rect 23662 28642 23714 28654
rect 29486 28642 29538 28654
rect 24322 28590 24334 28642
rect 24386 28590 24398 28642
rect 24994 28590 25006 28642
rect 25058 28590 25070 28642
rect 23662 28578 23714 28590
rect 29486 28578 29538 28590
rect 30158 28642 30210 28654
rect 34862 28642 34914 28654
rect 32610 28590 32622 28642
rect 32674 28590 32686 28642
rect 30158 28578 30210 28590
rect 34862 28578 34914 28590
rect 38558 28642 38610 28654
rect 38558 28578 38610 28590
rect 38894 28642 38946 28654
rect 39902 28642 39954 28654
rect 45502 28642 45554 28654
rect 39106 28590 39118 28642
rect 39170 28590 39182 28642
rect 40226 28590 40238 28642
rect 40290 28590 40302 28642
rect 40898 28590 40910 28642
rect 40962 28590 40974 28642
rect 41682 28590 41694 28642
rect 41746 28590 41758 28642
rect 38894 28578 38946 28590
rect 39902 28578 39954 28590
rect 45502 28578 45554 28590
rect 46286 28642 46338 28654
rect 47518 28642 47570 28654
rect 47058 28590 47070 28642
rect 47122 28590 47134 28642
rect 47954 28590 47966 28642
rect 48018 28590 48030 28642
rect 46286 28578 46338 28590
rect 47518 28578 47570 28590
rect 10670 28530 10722 28542
rect 10670 28466 10722 28478
rect 14478 28530 14530 28542
rect 14478 28466 14530 28478
rect 18174 28530 18226 28542
rect 18174 28466 18226 28478
rect 20526 28530 20578 28542
rect 20526 28466 20578 28478
rect 20750 28530 20802 28542
rect 23886 28530 23938 28542
rect 22642 28478 22654 28530
rect 22706 28478 22718 28530
rect 20750 28466 20802 28478
rect 23886 28466 23938 28478
rect 24110 28530 24162 28542
rect 24110 28466 24162 28478
rect 29822 28530 29874 28542
rect 34526 28530 34578 28542
rect 42702 28530 42754 28542
rect 31602 28478 31614 28530
rect 31666 28478 31678 28530
rect 39218 28478 39230 28530
rect 39282 28478 39294 28530
rect 41906 28478 41918 28530
rect 41970 28478 41982 28530
rect 29822 28466 29874 28478
rect 34526 28466 34578 28478
rect 42702 28466 42754 28478
rect 43038 28530 43090 28542
rect 46834 28478 46846 28530
rect 46898 28478 46910 28530
rect 43038 28466 43090 28478
rect 8094 28418 8146 28430
rect 8094 28354 8146 28366
rect 10446 28418 10498 28430
rect 10446 28354 10498 28366
rect 10782 28418 10834 28430
rect 10782 28354 10834 28366
rect 11566 28418 11618 28430
rect 11566 28354 11618 28366
rect 14590 28418 14642 28430
rect 14590 28354 14642 28366
rect 16718 28418 16770 28430
rect 16718 28354 16770 28366
rect 19630 28418 19682 28430
rect 35422 28418 35474 28430
rect 31714 28366 31726 28418
rect 31778 28366 31790 28418
rect 19630 28354 19682 28366
rect 35422 28354 35474 28366
rect 35982 28418 36034 28430
rect 35982 28354 36034 28366
rect 37998 28418 38050 28430
rect 41010 28366 41022 28418
rect 41074 28366 41086 28418
rect 37998 28354 38050 28366
rect 1344 28250 48720 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48720 28250
rect 1344 28164 48720 28198
rect 2494 28082 2546 28094
rect 9662 28082 9714 28094
rect 16494 28082 16546 28094
rect 8978 28030 8990 28082
rect 9042 28030 9054 28082
rect 13794 28030 13806 28082
rect 13858 28030 13870 28082
rect 2494 28018 2546 28030
rect 9662 28018 9714 28030
rect 16494 28018 16546 28030
rect 18622 28082 18674 28094
rect 22430 28082 22482 28094
rect 21970 28030 21982 28082
rect 22034 28030 22046 28082
rect 18622 28018 18674 28030
rect 22430 28018 22482 28030
rect 24110 28082 24162 28094
rect 24110 28018 24162 28030
rect 25342 28082 25394 28094
rect 25342 28018 25394 28030
rect 25454 28082 25506 28094
rect 31950 28082 32002 28094
rect 29922 28030 29934 28082
rect 29986 28030 29998 28082
rect 30258 28030 30270 28082
rect 30322 28030 30334 28082
rect 25454 28018 25506 28030
rect 31950 28018 32002 28030
rect 42478 28082 42530 28094
rect 42478 28018 42530 28030
rect 45502 28082 45554 28094
rect 45502 28018 45554 28030
rect 47182 28082 47234 28094
rect 47182 28018 47234 28030
rect 9774 27970 9826 27982
rect 14478 27970 14530 27982
rect 5170 27918 5182 27970
rect 5234 27918 5246 27970
rect 10098 27918 10110 27970
rect 10162 27918 10174 27970
rect 14130 27918 14142 27970
rect 14194 27918 14206 27970
rect 9774 27906 9826 27918
rect 14478 27906 14530 27918
rect 14814 27970 14866 27982
rect 26014 27970 26066 27982
rect 16818 27918 16830 27970
rect 16882 27918 16894 27970
rect 14814 27906 14866 27918
rect 26014 27906 26066 27918
rect 30606 27970 30658 27982
rect 33506 27918 33518 27970
rect 33570 27918 33582 27970
rect 44482 27918 44494 27970
rect 44546 27918 44558 27970
rect 46050 27918 46062 27970
rect 46114 27918 46126 27970
rect 46386 27918 46398 27970
rect 46450 27918 46462 27970
rect 30606 27906 30658 27918
rect 2830 27858 2882 27870
rect 2830 27794 2882 27806
rect 4062 27858 4114 27870
rect 4062 27794 4114 27806
rect 4398 27858 4450 27870
rect 9438 27858 9490 27870
rect 17390 27858 17442 27870
rect 4834 27806 4846 27858
rect 4898 27806 4910 27858
rect 6066 27806 6078 27858
rect 6130 27806 6142 27858
rect 6626 27806 6638 27858
rect 6690 27806 6702 27858
rect 10322 27806 10334 27858
rect 10386 27806 10398 27858
rect 10882 27806 10894 27858
rect 10946 27806 10958 27858
rect 11442 27806 11454 27858
rect 11506 27806 11518 27858
rect 15026 27806 15038 27858
rect 15090 27806 15102 27858
rect 4398 27794 4450 27806
rect 9438 27794 9490 27806
rect 17390 27794 17442 27806
rect 17726 27858 17778 27870
rect 26350 27858 26402 27870
rect 18162 27806 18174 27858
rect 18226 27806 18238 27858
rect 19058 27806 19070 27858
rect 19122 27806 19134 27858
rect 19618 27806 19630 27858
rect 19682 27806 19694 27858
rect 17726 27794 17778 27806
rect 26350 27794 26402 27806
rect 26574 27858 26626 27870
rect 34638 27858 34690 27870
rect 27010 27806 27022 27858
rect 27074 27806 27086 27858
rect 27458 27806 27470 27858
rect 27522 27806 27534 27858
rect 31378 27806 31390 27858
rect 31442 27806 31454 27858
rect 33618 27806 33630 27858
rect 33682 27806 33694 27858
rect 26574 27794 26626 27806
rect 34638 27794 34690 27806
rect 35198 27858 35250 27870
rect 42366 27858 42418 27870
rect 35634 27806 35646 27858
rect 35698 27806 35710 27858
rect 38882 27806 38894 27858
rect 38946 27806 38958 27858
rect 41122 27806 41134 27858
rect 41186 27806 41198 27858
rect 42690 27806 42702 27858
rect 42754 27806 42766 27858
rect 44706 27806 44718 27858
rect 44770 27806 44782 27858
rect 35198 27794 35250 27806
rect 42366 27794 42418 27806
rect 17502 27746 17554 27758
rect 17502 27682 17554 27694
rect 17838 27746 17890 27758
rect 17838 27682 17890 27694
rect 26126 27746 26178 27758
rect 26126 27682 26178 27694
rect 30942 27746 30994 27758
rect 39566 27746 39618 27758
rect 33170 27694 33182 27746
rect 33234 27694 33246 27746
rect 34178 27694 34190 27746
rect 34242 27694 34254 27746
rect 36082 27694 36094 27746
rect 36146 27694 36158 27746
rect 38210 27694 38222 27746
rect 38274 27694 38286 27746
rect 30942 27682 30994 27694
rect 39566 27682 39618 27694
rect 40350 27746 40402 27758
rect 40350 27682 40402 27694
rect 48302 27746 48354 27758
rect 48302 27682 48354 27694
rect 25566 27634 25618 27646
rect 25566 27570 25618 27582
rect 45838 27634 45890 27646
rect 45838 27570 45890 27582
rect 1344 27466 48720 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48720 27466
rect 1344 27380 48720 27414
rect 21646 27298 21698 27310
rect 17490 27246 17502 27298
rect 17554 27246 17566 27298
rect 21646 27234 21698 27246
rect 24446 27298 24498 27310
rect 24446 27234 24498 27246
rect 26574 27298 26626 27310
rect 26574 27234 26626 27246
rect 36990 27298 37042 27310
rect 36990 27234 37042 27246
rect 37326 27298 37378 27310
rect 37326 27234 37378 27246
rect 43038 27298 43090 27310
rect 43038 27234 43090 27246
rect 9998 27186 10050 27198
rect 20638 27186 20690 27198
rect 11106 27134 11118 27186
rect 11170 27134 11182 27186
rect 11666 27134 11678 27186
rect 11730 27134 11742 27186
rect 16594 27134 16606 27186
rect 16658 27134 16670 27186
rect 9998 27122 10050 27134
rect 20638 27122 20690 27134
rect 26686 27186 26738 27198
rect 26686 27122 26738 27134
rect 27358 27186 27410 27198
rect 38446 27186 38498 27198
rect 30482 27134 30494 27186
rect 30546 27134 30558 27186
rect 32610 27134 32622 27186
rect 32674 27134 32686 27186
rect 27358 27122 27410 27134
rect 38446 27122 38498 27134
rect 38894 27186 38946 27198
rect 38894 27122 38946 27134
rect 42702 27186 42754 27198
rect 42702 27122 42754 27134
rect 4174 27074 4226 27086
rect 9326 27074 9378 27086
rect 4834 27022 4846 27074
rect 4898 27022 4910 27074
rect 5618 27022 5630 27074
rect 5682 27022 5694 27074
rect 8082 27022 8094 27074
rect 8146 27022 8158 27074
rect 8754 27022 8766 27074
rect 8818 27022 8830 27074
rect 4174 27010 4226 27022
rect 9326 27010 9378 27022
rect 9438 27074 9490 27086
rect 11566 27074 11618 27086
rect 10770 27022 10782 27074
rect 10834 27022 10846 27074
rect 12002 27022 12014 27074
rect 12066 27022 12078 27074
rect 13682 27022 13694 27074
rect 13746 27022 13758 27074
rect 14130 27034 14142 27086
rect 14194 27034 14206 27086
rect 19630 27074 19682 27086
rect 17714 27022 17726 27074
rect 17778 27022 17790 27074
rect 9438 27010 9490 27022
rect 11566 27010 11618 27022
rect 19630 27010 19682 27022
rect 19742 27074 19794 27086
rect 19742 27010 19794 27022
rect 20302 27074 20354 27086
rect 33966 27074 34018 27086
rect 35086 27074 35138 27086
rect 39230 27074 39282 27086
rect 21298 27022 21310 27074
rect 21362 27022 21374 27074
rect 26898 27022 26910 27074
rect 26962 27022 26974 27074
rect 30818 27022 30830 27074
rect 30882 27022 30894 27074
rect 31266 27022 31278 27074
rect 31330 27022 31342 27074
rect 32946 27022 32958 27074
rect 33010 27022 33022 27074
rect 34850 27022 34862 27074
rect 34914 27022 34926 27074
rect 37874 27022 37886 27074
rect 37938 27022 37950 27074
rect 20302 27010 20354 27022
rect 33966 27010 34018 27022
rect 35086 27010 35138 27022
rect 39230 27010 39282 27022
rect 39454 27074 39506 27086
rect 39454 27010 39506 27022
rect 39902 27074 39954 27086
rect 41582 27074 41634 27086
rect 40674 27022 40686 27074
rect 40738 27022 40750 27074
rect 41234 27022 41246 27074
rect 41298 27022 41310 27074
rect 39902 27010 39954 27022
rect 41582 27010 41634 27022
rect 41918 27074 41970 27086
rect 41918 27010 41970 27022
rect 42254 27074 42306 27086
rect 42254 27010 42306 27022
rect 43374 27074 43426 27086
rect 47182 27074 47234 27086
rect 44146 27022 44158 27074
rect 44210 27022 44222 27074
rect 43374 27010 43426 27022
rect 47182 27010 47234 27022
rect 2606 26962 2658 26974
rect 2606 26898 2658 26910
rect 3838 26962 3890 26974
rect 8990 26962 9042 26974
rect 4722 26910 4734 26962
rect 4786 26910 4798 26962
rect 3838 26898 3890 26910
rect 8990 26898 9042 26910
rect 9550 26962 9602 26974
rect 9550 26898 9602 26910
rect 12686 26962 12738 26974
rect 12686 26898 12738 26910
rect 16942 26962 16994 26974
rect 23662 26962 23714 26974
rect 17154 26910 17166 26962
rect 17218 26910 17230 26962
rect 16942 26898 16994 26910
rect 23662 26898 23714 26910
rect 23774 26962 23826 26974
rect 23774 26898 23826 26910
rect 24558 26962 24610 26974
rect 24558 26898 24610 26910
rect 25118 26962 25170 26974
rect 29486 26962 29538 26974
rect 35198 26962 35250 26974
rect 29138 26910 29150 26962
rect 29202 26910 29214 26962
rect 31602 26910 31614 26962
rect 31666 26910 31678 26962
rect 31826 26910 31838 26962
rect 31890 26910 31902 26962
rect 25118 26898 25170 26910
rect 29486 26898 29538 26910
rect 35198 26898 35250 26910
rect 37214 26962 37266 26974
rect 46398 26962 46450 26974
rect 37650 26910 37662 26962
rect 37714 26910 37726 26962
rect 40114 26910 40126 26962
rect 40178 26910 40190 26962
rect 44034 26910 44046 26962
rect 44098 26910 44110 26962
rect 37214 26898 37266 26910
rect 46398 26898 46450 26910
rect 46846 26962 46898 26974
rect 47394 26910 47406 26962
rect 47458 26910 47470 26962
rect 47954 26910 47966 26962
rect 48018 26910 48030 26962
rect 46846 26898 46898 26910
rect 2270 26850 2322 26862
rect 2270 26786 2322 26798
rect 17726 26850 17778 26862
rect 17726 26786 17778 26798
rect 19854 26850 19906 26862
rect 19854 26786 19906 26798
rect 21534 26850 21586 26862
rect 21534 26786 21586 26798
rect 23438 26850 23490 26862
rect 23438 26786 23490 26798
rect 30046 26850 30098 26862
rect 39678 26850 39730 26862
rect 42030 26850 42082 26862
rect 35634 26798 35646 26850
rect 35698 26798 35710 26850
rect 41122 26798 41134 26850
rect 41186 26798 41198 26850
rect 30046 26786 30098 26798
rect 39678 26786 39730 26798
rect 42030 26786 42082 26798
rect 46062 26850 46114 26862
rect 46062 26786 46114 26798
rect 1344 26682 48720 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48720 26682
rect 1344 26596 48720 26630
rect 8878 26514 8930 26526
rect 8878 26450 8930 26462
rect 12462 26514 12514 26526
rect 12462 26450 12514 26462
rect 14142 26514 14194 26526
rect 14142 26450 14194 26462
rect 18510 26514 18562 26526
rect 18510 26450 18562 26462
rect 19854 26514 19906 26526
rect 19854 26450 19906 26462
rect 20750 26514 20802 26526
rect 32398 26514 32450 26526
rect 24658 26462 24670 26514
rect 24722 26462 24734 26514
rect 30818 26462 30830 26514
rect 30882 26462 30894 26514
rect 20750 26450 20802 26462
rect 32398 26450 32450 26462
rect 35310 26514 35362 26526
rect 35310 26450 35362 26462
rect 39902 26514 39954 26526
rect 39902 26450 39954 26462
rect 40350 26514 40402 26526
rect 40350 26450 40402 26462
rect 40798 26514 40850 26526
rect 48290 26462 48302 26514
rect 48354 26462 48366 26514
rect 40798 26450 40850 26462
rect 9998 26402 10050 26414
rect 9998 26338 10050 26350
rect 10110 26402 10162 26414
rect 10110 26338 10162 26350
rect 10670 26402 10722 26414
rect 20190 26402 20242 26414
rect 18834 26350 18846 26402
rect 18898 26350 18910 26402
rect 10670 26338 10722 26350
rect 20190 26338 20242 26350
rect 31502 26402 31554 26414
rect 31502 26338 31554 26350
rect 33630 26402 33682 26414
rect 33630 26338 33682 26350
rect 33966 26402 34018 26414
rect 33966 26338 34018 26350
rect 37326 26402 37378 26414
rect 42018 26350 42030 26402
rect 42082 26350 42094 26402
rect 42690 26350 42702 26402
rect 42754 26350 42766 26402
rect 37326 26338 37378 26350
rect 5182 26290 5234 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 2258 26238 2270 26290
rect 2322 26238 2334 26290
rect 5182 26226 5234 26238
rect 10334 26290 10386 26302
rect 10334 26226 10386 26238
rect 13806 26290 13858 26302
rect 13806 26226 13858 26238
rect 14254 26290 14306 26302
rect 14254 26226 14306 26238
rect 14478 26290 14530 26302
rect 14478 26226 14530 26238
rect 14926 26290 14978 26302
rect 17614 26290 17666 26302
rect 15138 26238 15150 26290
rect 15202 26238 15214 26290
rect 14926 26226 14978 26238
rect 17614 26226 17666 26238
rect 17838 26290 17890 26302
rect 17838 26226 17890 26238
rect 19518 26290 19570 26302
rect 19518 26226 19570 26238
rect 19854 26290 19906 26302
rect 31166 26290 31218 26302
rect 21634 26238 21646 26290
rect 21698 26238 21710 26290
rect 22194 26238 22206 26290
rect 22258 26238 22270 26290
rect 25218 26238 25230 26290
rect 25282 26238 25294 26290
rect 19854 26226 19906 26238
rect 31166 26226 31218 26238
rect 31838 26290 31890 26302
rect 31838 26226 31890 26238
rect 33406 26290 33458 26302
rect 40898 26238 40910 26290
rect 40962 26238 40974 26290
rect 41906 26238 41918 26290
rect 41970 26238 41982 26290
rect 43026 26238 43038 26290
rect 43090 26238 43102 26290
rect 45154 26238 45166 26290
rect 45218 26238 45230 26290
rect 45938 26238 45950 26290
rect 46002 26238 46014 26290
rect 33406 26226 33458 26238
rect 9662 26178 9714 26190
rect 4722 26126 4734 26178
rect 4786 26126 4798 26178
rect 8978 26126 8990 26178
rect 9042 26126 9054 26178
rect 9662 26114 9714 26126
rect 11118 26178 11170 26190
rect 11118 26114 11170 26126
rect 16606 26178 16658 26190
rect 16606 26114 16658 26126
rect 17390 26178 17442 26190
rect 17390 26114 17442 26126
rect 19294 26178 19346 26190
rect 44942 26178 44994 26190
rect 28690 26126 28702 26178
rect 28754 26126 28766 26178
rect 34402 26126 34414 26178
rect 34466 26126 34478 26178
rect 35746 26126 35758 26178
rect 35810 26126 35822 26178
rect 19294 26114 19346 26126
rect 44942 26114 44994 26126
rect 8654 26066 8706 26078
rect 14814 26066 14866 26078
rect 10434 26014 10446 26066
rect 10498 26063 10510 26066
rect 10882 26063 10894 26066
rect 10498 26017 10894 26063
rect 10498 26014 10510 26017
rect 10882 26014 10894 26017
rect 10946 26014 10958 26066
rect 8654 26002 8706 26014
rect 14814 26002 14866 26014
rect 18286 26066 18338 26078
rect 18286 26002 18338 26014
rect 33070 26066 33122 26078
rect 33070 26002 33122 26014
rect 37438 26066 37490 26078
rect 37438 26002 37490 26014
rect 1344 25898 48720 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48720 25898
rect 1344 25812 48720 25846
rect 8654 25730 8706 25742
rect 8654 25666 8706 25678
rect 18286 25730 18338 25742
rect 31502 25730 31554 25742
rect 25890 25678 25902 25730
rect 25954 25678 25966 25730
rect 18286 25666 18338 25678
rect 31502 25666 31554 25678
rect 42702 25730 42754 25742
rect 42702 25666 42754 25678
rect 45838 25730 45890 25742
rect 45838 25666 45890 25678
rect 12014 25618 12066 25630
rect 23102 25618 23154 25630
rect 9650 25566 9662 25618
rect 9714 25566 9726 25618
rect 13570 25566 13582 25618
rect 13634 25566 13646 25618
rect 12014 25554 12066 25566
rect 23102 25554 23154 25566
rect 24222 25618 24274 25630
rect 28030 25618 28082 25630
rect 30830 25618 30882 25630
rect 45390 25618 45442 25630
rect 26898 25566 26910 25618
rect 26962 25566 26974 25618
rect 29810 25566 29822 25618
rect 29874 25566 29886 25618
rect 36978 25566 36990 25618
rect 37042 25566 37054 25618
rect 24222 25554 24274 25566
rect 28030 25554 28082 25566
rect 30830 25554 30882 25566
rect 45390 25554 45442 25566
rect 10894 25506 10946 25518
rect 8306 25454 8318 25506
rect 8370 25454 8382 25506
rect 9202 25454 9214 25506
rect 9266 25454 9278 25506
rect 10322 25454 10334 25506
rect 10386 25454 10398 25506
rect 10894 25442 10946 25454
rect 12350 25506 12402 25518
rect 12350 25442 12402 25454
rect 12910 25506 12962 25518
rect 18398 25506 18450 25518
rect 13458 25454 13470 25506
rect 13522 25454 13534 25506
rect 12910 25442 12962 25454
rect 18398 25442 18450 25454
rect 18622 25506 18674 25518
rect 22430 25506 22482 25518
rect 19730 25454 19742 25506
rect 19794 25454 19806 25506
rect 18622 25442 18674 25454
rect 22430 25442 22482 25454
rect 23214 25506 23266 25518
rect 25342 25506 25394 25518
rect 26574 25506 26626 25518
rect 28142 25506 28194 25518
rect 23538 25454 23550 25506
rect 23602 25454 23614 25506
rect 25554 25454 25566 25506
rect 25618 25454 25630 25506
rect 26114 25454 26126 25506
rect 26178 25454 26190 25506
rect 27010 25454 27022 25506
rect 27074 25454 27086 25506
rect 27794 25454 27806 25506
rect 27858 25454 27870 25506
rect 23214 25442 23266 25454
rect 25342 25442 25394 25454
rect 26574 25442 26626 25454
rect 28142 25442 28194 25454
rect 28478 25506 28530 25518
rect 28478 25442 28530 25454
rect 29374 25506 29426 25518
rect 29374 25442 29426 25454
rect 30270 25506 30322 25518
rect 30270 25442 30322 25454
rect 31838 25506 31890 25518
rect 41918 25506 41970 25518
rect 39890 25454 39902 25506
rect 39954 25454 39966 25506
rect 31838 25442 31890 25454
rect 41918 25442 41970 25454
rect 43038 25506 43090 25518
rect 46174 25506 46226 25518
rect 43586 25454 43598 25506
rect 43650 25454 43662 25506
rect 43038 25442 43090 25454
rect 46174 25442 46226 25454
rect 9886 25394 9938 25406
rect 9886 25330 9938 25342
rect 9998 25394 10050 25406
rect 9998 25330 10050 25342
rect 11342 25394 11394 25406
rect 11342 25330 11394 25342
rect 11566 25394 11618 25406
rect 11566 25330 11618 25342
rect 12686 25394 12738 25406
rect 12686 25330 12738 25342
rect 13806 25394 13858 25406
rect 13806 25330 13858 25342
rect 18286 25394 18338 25406
rect 18286 25330 18338 25342
rect 19294 25394 19346 25406
rect 21310 25394 21362 25406
rect 19954 25342 19966 25394
rect 20018 25342 20030 25394
rect 19294 25330 19346 25342
rect 21310 25330 21362 25342
rect 22318 25394 22370 25406
rect 22318 25330 22370 25342
rect 22990 25394 23042 25406
rect 22990 25330 23042 25342
rect 24446 25394 24498 25406
rect 24446 25330 24498 25342
rect 24558 25394 24610 25406
rect 31278 25394 31330 25406
rect 27122 25342 27134 25394
rect 27186 25342 27198 25394
rect 24558 25330 24610 25342
rect 31278 25330 31330 25342
rect 32734 25394 32786 25406
rect 39106 25342 39118 25394
rect 39170 25342 39182 25394
rect 43810 25342 43822 25394
rect 43874 25342 43886 25394
rect 46498 25342 46510 25394
rect 46562 25342 46574 25394
rect 46946 25342 46958 25394
rect 47010 25342 47022 25394
rect 32734 25330 32786 25342
rect 8542 25282 8594 25294
rect 8542 25218 8594 25230
rect 11230 25282 11282 25294
rect 11230 25218 11282 25230
rect 12462 25282 12514 25294
rect 12462 25218 12514 25230
rect 19070 25282 19122 25294
rect 19070 25218 19122 25230
rect 19182 25282 19234 25294
rect 19182 25218 19234 25230
rect 20414 25282 20466 25294
rect 20414 25218 20466 25230
rect 21422 25282 21474 25294
rect 21422 25218 21474 25230
rect 21534 25282 21586 25294
rect 21534 25218 21586 25230
rect 21758 25282 21810 25294
rect 21758 25218 21810 25230
rect 22094 25282 22146 25294
rect 22094 25218 22146 25230
rect 24782 25282 24834 25294
rect 24782 25218 24834 25230
rect 25454 25282 25506 25294
rect 25454 25218 25506 25230
rect 26798 25282 26850 25294
rect 26798 25218 26850 25230
rect 27694 25282 27746 25294
rect 27694 25218 27746 25230
rect 31390 25282 31442 25294
rect 31390 25218 31442 25230
rect 32174 25282 32226 25294
rect 32174 25218 32226 25230
rect 32398 25282 32450 25294
rect 32398 25218 32450 25230
rect 32622 25282 32674 25294
rect 32622 25218 32674 25230
rect 40350 25282 40402 25294
rect 40350 25218 40402 25230
rect 42254 25282 42306 25294
rect 42254 25218 42306 25230
rect 1344 25114 48720 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48720 25114
rect 1344 25028 48720 25062
rect 10894 24946 10946 24958
rect 20750 24946 20802 24958
rect 9426 24894 9438 24946
rect 9490 24894 9502 24946
rect 14242 24894 14254 24946
rect 14306 24894 14318 24946
rect 8990 24722 9042 24734
rect 1922 24670 1934 24722
rect 1986 24670 1998 24722
rect 2594 24670 2606 24722
rect 2658 24670 2670 24722
rect 7970 24670 7982 24722
rect 8034 24670 8046 24722
rect 8530 24670 8542 24722
rect 8594 24670 8606 24722
rect 8990 24658 9042 24670
rect 4946 24558 4958 24610
rect 5010 24558 5022 24610
rect 5506 24558 5518 24610
rect 5570 24558 5582 24610
rect 9441 24495 9487 24894
rect 10894 24882 10946 24894
rect 20750 24882 20802 24894
rect 23998 24946 24050 24958
rect 23998 24882 24050 24894
rect 27134 24946 27186 24958
rect 27134 24882 27186 24894
rect 28814 24946 28866 24958
rect 28814 24882 28866 24894
rect 29710 24946 29762 24958
rect 29710 24882 29762 24894
rect 31054 24946 31106 24958
rect 31054 24882 31106 24894
rect 40350 24946 40402 24958
rect 45154 24894 45166 24946
rect 45218 24894 45230 24946
rect 40350 24882 40402 24894
rect 9886 24834 9938 24846
rect 9886 24770 9938 24782
rect 24222 24834 24274 24846
rect 24222 24770 24274 24782
rect 26350 24834 26402 24846
rect 26350 24770 26402 24782
rect 26798 24834 26850 24846
rect 26798 24770 26850 24782
rect 30046 24834 30098 24846
rect 40910 24834 40962 24846
rect 35746 24782 35758 24834
rect 35810 24782 35822 24834
rect 36754 24782 36766 24834
rect 36818 24782 36830 24834
rect 38546 24782 38558 24834
rect 38610 24782 38622 24834
rect 30046 24770 30098 24782
rect 40910 24770 40962 24782
rect 9774 24722 9826 24734
rect 14702 24722 14754 24734
rect 20862 24722 20914 24734
rect 11330 24670 11342 24722
rect 11394 24670 11406 24722
rect 11890 24670 11902 24722
rect 11954 24670 11966 24722
rect 17490 24670 17502 24722
rect 17554 24670 17566 24722
rect 18050 24670 18062 24722
rect 18114 24670 18126 24722
rect 20402 24670 20414 24722
rect 20466 24670 20478 24722
rect 9774 24658 9826 24670
rect 14702 24658 14754 24670
rect 20862 24658 20914 24670
rect 24670 24722 24722 24734
rect 24670 24658 24722 24670
rect 27134 24722 27186 24734
rect 27134 24658 27186 24670
rect 27470 24722 27522 24734
rect 27470 24658 27522 24670
rect 29150 24722 29202 24734
rect 29150 24658 29202 24670
rect 30382 24722 30434 24734
rect 30382 24658 30434 24670
rect 30494 24722 30546 24734
rect 30494 24658 30546 24670
rect 32286 24722 32338 24734
rect 41134 24722 41186 24734
rect 35970 24670 35982 24722
rect 36034 24670 36046 24722
rect 36530 24670 36542 24722
rect 36594 24670 36606 24722
rect 38770 24670 38782 24722
rect 38834 24670 38846 24722
rect 42018 24670 42030 24722
rect 42082 24670 42094 24722
rect 42690 24670 42702 24722
rect 42754 24670 42766 24722
rect 32286 24658 32338 24670
rect 41134 24658 41186 24670
rect 10446 24610 10498 24622
rect 10446 24546 10498 24558
rect 15150 24610 15202 24622
rect 15150 24546 15202 24558
rect 24110 24610 24162 24622
rect 24110 24546 24162 24558
rect 26462 24610 26514 24622
rect 26462 24546 26514 24558
rect 27806 24610 27858 24622
rect 27806 24546 27858 24558
rect 28254 24610 28306 24622
rect 28254 24546 28306 24558
rect 30158 24610 30210 24622
rect 30158 24546 30210 24558
rect 31614 24610 31666 24622
rect 31614 24546 31666 24558
rect 32510 24610 32562 24622
rect 32510 24546 32562 24558
rect 45614 24610 45666 24622
rect 45614 24546 45666 24558
rect 9886 24498 9938 24510
rect 36318 24498 36370 24510
rect 9538 24495 9550 24498
rect 9441 24449 9550 24495
rect 9538 24446 9550 24449
rect 9602 24446 9614 24498
rect 10322 24446 10334 24498
rect 10386 24495 10398 24498
rect 10994 24495 11006 24498
rect 10386 24449 11006 24495
rect 10386 24446 10398 24449
rect 10994 24446 11006 24449
rect 11058 24446 11070 24498
rect 31938 24446 31950 24498
rect 32002 24446 32014 24498
rect 9886 24434 9938 24446
rect 36318 24434 36370 24446
rect 41470 24498 41522 24510
rect 41470 24434 41522 24446
rect 1344 24330 48720 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48720 24330
rect 1344 24244 48720 24278
rect 15486 24162 15538 24174
rect 12114 24110 12126 24162
rect 12178 24110 12190 24162
rect 15486 24098 15538 24110
rect 22094 24162 22146 24174
rect 22094 24098 22146 24110
rect 38334 24162 38386 24174
rect 38334 24098 38386 24110
rect 38670 24162 38722 24174
rect 41346 24110 41358 24162
rect 41410 24110 41422 24162
rect 38670 24098 38722 24110
rect 5742 24050 5794 24062
rect 5742 23986 5794 23998
rect 7758 24050 7810 24062
rect 7758 23986 7810 23998
rect 8094 24050 8146 24062
rect 8094 23986 8146 23998
rect 13582 24050 13634 24062
rect 26798 24050 26850 24062
rect 26450 23998 26462 24050
rect 26514 23998 26526 24050
rect 13582 23986 13634 23998
rect 26798 23986 26850 23998
rect 28366 24050 28418 24062
rect 28366 23986 28418 23998
rect 30942 24050 30994 24062
rect 30942 23986 30994 23998
rect 31278 24050 31330 24062
rect 36430 24050 36482 24062
rect 32610 23998 32622 24050
rect 32674 23998 32686 24050
rect 33842 23998 33854 24050
rect 33906 23998 33918 24050
rect 35970 23998 35982 24050
rect 36034 23998 36046 24050
rect 31278 23986 31330 23998
rect 36430 23986 36482 23998
rect 4174 23938 4226 23950
rect 7870 23938 7922 23950
rect 4946 23886 4958 23938
rect 5010 23886 5022 23938
rect 4174 23874 4226 23886
rect 7870 23874 7922 23886
rect 8206 23938 8258 23950
rect 8206 23874 8258 23886
rect 8430 23938 8482 23950
rect 8430 23874 8482 23886
rect 9438 23938 9490 23950
rect 9438 23874 9490 23886
rect 9998 23938 10050 23950
rect 9998 23874 10050 23886
rect 10334 23938 10386 23950
rect 10334 23874 10386 23886
rect 10558 23938 10610 23950
rect 12126 23938 12178 23950
rect 14142 23938 14194 23950
rect 10770 23886 10782 23938
rect 10834 23886 10846 23938
rect 11666 23886 11678 23938
rect 11730 23886 11742 23938
rect 12226 23886 12238 23938
rect 12290 23886 12302 23938
rect 10558 23874 10610 23886
rect 12126 23874 12178 23886
rect 14142 23874 14194 23886
rect 14478 23938 14530 23950
rect 14478 23874 14530 23886
rect 14702 23938 14754 23950
rect 14702 23874 14754 23886
rect 15150 23938 15202 23950
rect 15150 23874 15202 23886
rect 16046 23938 16098 23950
rect 16046 23874 16098 23886
rect 16382 23938 16434 23950
rect 29150 23938 29202 23950
rect 37102 23938 37154 23950
rect 40686 23938 40738 23950
rect 23314 23886 23326 23938
rect 23378 23886 23390 23938
rect 24098 23886 24110 23938
rect 24162 23886 24174 23938
rect 29586 23886 29598 23938
rect 29650 23886 29662 23938
rect 33170 23886 33182 23938
rect 33234 23886 33246 23938
rect 37426 23886 37438 23938
rect 37490 23886 37502 23938
rect 39218 23886 39230 23938
rect 39282 23886 39294 23938
rect 40450 23886 40462 23938
rect 40514 23886 40526 23938
rect 41458 23886 41470 23938
rect 41522 23886 41534 23938
rect 16382 23874 16434 23886
rect 29150 23874 29202 23886
rect 37102 23874 37154 23886
rect 40686 23874 40738 23886
rect 2606 23826 2658 23838
rect 2606 23762 2658 23774
rect 2942 23826 2994 23838
rect 2942 23762 2994 23774
rect 3838 23826 3890 23838
rect 8990 23826 9042 23838
rect 4834 23774 4846 23826
rect 4898 23774 4910 23826
rect 3838 23762 3890 23774
rect 8990 23762 9042 23774
rect 9102 23826 9154 23838
rect 9102 23762 9154 23774
rect 9550 23826 9602 23838
rect 9550 23762 9602 23774
rect 14030 23826 14082 23838
rect 14030 23762 14082 23774
rect 15374 23826 15426 23838
rect 15374 23762 15426 23774
rect 15486 23826 15538 23838
rect 15486 23762 15538 23774
rect 16718 23826 16770 23838
rect 16718 23762 16770 23774
rect 17054 23826 17106 23838
rect 17054 23762 17106 23774
rect 22206 23826 22258 23838
rect 22206 23762 22258 23774
rect 30046 23826 30098 23838
rect 30046 23762 30098 23774
rect 30382 23826 30434 23838
rect 30382 23762 30434 23774
rect 32398 23826 32450 23838
rect 32398 23762 32450 23774
rect 37998 23826 38050 23838
rect 37998 23762 38050 23774
rect 38558 23826 38610 23838
rect 38558 23762 38610 23774
rect 39678 23826 39730 23838
rect 39678 23762 39730 23774
rect 41694 23826 41746 23838
rect 41694 23762 41746 23774
rect 46734 23826 46786 23838
rect 46734 23762 46786 23774
rect 8766 23714 8818 23726
rect 8766 23650 8818 23662
rect 9774 23714 9826 23726
rect 9774 23650 9826 23662
rect 10110 23714 10162 23726
rect 10110 23650 10162 23662
rect 13806 23714 13858 23726
rect 13806 23650 13858 23662
rect 14590 23714 14642 23726
rect 14590 23650 14642 23662
rect 16270 23714 16322 23726
rect 16270 23650 16322 23662
rect 17166 23714 17218 23726
rect 17166 23650 17218 23662
rect 17614 23714 17666 23726
rect 17614 23650 17666 23662
rect 27358 23714 27410 23726
rect 27358 23650 27410 23662
rect 27806 23714 27858 23726
rect 27806 23650 27858 23662
rect 32174 23714 32226 23726
rect 32174 23650 32226 23662
rect 32622 23714 32674 23726
rect 32622 23650 32674 23662
rect 46398 23714 46450 23726
rect 46398 23650 46450 23662
rect 1344 23546 48720 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48720 23546
rect 1344 23460 48720 23494
rect 7982 23378 8034 23390
rect 7982 23314 8034 23326
rect 9102 23378 9154 23390
rect 9102 23314 9154 23326
rect 10222 23378 10274 23390
rect 10222 23314 10274 23326
rect 10782 23378 10834 23390
rect 10782 23314 10834 23326
rect 11678 23378 11730 23390
rect 11678 23314 11730 23326
rect 12910 23378 12962 23390
rect 31054 23378 31106 23390
rect 16818 23326 16830 23378
rect 16882 23326 16894 23378
rect 23090 23326 23102 23378
rect 23154 23326 23166 23378
rect 12910 23314 12962 23326
rect 31054 23314 31106 23326
rect 34078 23378 34130 23390
rect 34078 23314 34130 23326
rect 38782 23378 38834 23390
rect 48290 23326 48302 23378
rect 48354 23326 48366 23378
rect 38782 23314 38834 23326
rect 10446 23266 10498 23278
rect 5842 23214 5854 23266
rect 5906 23214 5918 23266
rect 6402 23214 6414 23266
rect 6466 23214 6478 23266
rect 10446 23202 10498 23214
rect 11230 23266 11282 23278
rect 11230 23202 11282 23214
rect 27022 23266 27074 23278
rect 27022 23202 27074 23214
rect 27358 23266 27410 23278
rect 27358 23202 27410 23214
rect 30158 23266 30210 23278
rect 34526 23266 34578 23278
rect 36542 23266 36594 23278
rect 31714 23214 31726 23266
rect 31778 23214 31790 23266
rect 36082 23214 36094 23266
rect 36146 23214 36158 23266
rect 30158 23202 30210 23214
rect 34526 23202 34578 23214
rect 36542 23202 36594 23214
rect 36766 23266 36818 23278
rect 36766 23202 36818 23214
rect 40350 23266 40402 23278
rect 42130 23214 42142 23266
rect 42194 23214 42206 23266
rect 44146 23214 44158 23266
rect 44210 23214 44222 23266
rect 44706 23214 44718 23266
rect 44770 23214 44782 23266
rect 40350 23202 40402 23214
rect 5630 23154 5682 23166
rect 1810 23102 1822 23154
rect 1874 23102 1886 23154
rect 2258 23102 2270 23154
rect 2322 23102 2334 23154
rect 4722 23102 4734 23154
rect 4786 23102 4798 23154
rect 5630 23090 5682 23102
rect 8206 23154 8258 23166
rect 8206 23090 8258 23102
rect 8654 23154 8706 23166
rect 8654 23090 8706 23102
rect 10110 23154 10162 23166
rect 10110 23090 10162 23102
rect 10558 23154 10610 23166
rect 10558 23090 10610 23102
rect 10894 23154 10946 23166
rect 10894 23090 10946 23102
rect 12126 23154 12178 23166
rect 12126 23090 12178 23102
rect 13022 23154 13074 23166
rect 13022 23090 13074 23102
rect 13134 23154 13186 23166
rect 13134 23090 13186 23102
rect 13582 23154 13634 23166
rect 17390 23154 17442 23166
rect 13906 23102 13918 23154
rect 13970 23102 13982 23154
rect 14466 23102 14478 23154
rect 14530 23102 14542 23154
rect 13582 23090 13634 23102
rect 17390 23090 17442 23102
rect 17950 23154 18002 23166
rect 30270 23154 30322 23166
rect 41022 23154 41074 23166
rect 20178 23102 20190 23154
rect 20242 23102 20254 23154
rect 20738 23102 20750 23154
rect 20802 23102 20814 23154
rect 26562 23102 26574 23154
rect 26626 23102 26638 23154
rect 31826 23102 31838 23154
rect 31890 23102 31902 23154
rect 34738 23102 34750 23154
rect 34802 23102 34814 23154
rect 35746 23102 35758 23154
rect 35810 23102 35822 23154
rect 40114 23102 40126 23154
rect 40178 23102 40190 23154
rect 17950 23090 18002 23102
rect 30270 23090 30322 23102
rect 41022 23090 41074 23102
rect 41358 23154 41410 23166
rect 41906 23102 41918 23154
rect 41970 23102 41982 23154
rect 45154 23102 45166 23154
rect 45218 23102 45230 23154
rect 45938 23102 45950 23154
rect 46002 23102 46014 23154
rect 41358 23090 41410 23102
rect 8094 23042 8146 23054
rect 8094 22978 8146 22990
rect 9774 23042 9826 23054
rect 9774 22978 9826 22990
rect 12574 23042 12626 23054
rect 32510 23042 32562 23054
rect 26226 22990 26238 23042
rect 26290 22990 26302 23042
rect 31938 22990 31950 23042
rect 32002 22990 32014 23042
rect 12574 22978 12626 22990
rect 32510 22978 32562 22990
rect 34190 23042 34242 23054
rect 34190 22978 34242 22990
rect 37326 23042 37378 23054
rect 37326 22978 37378 22990
rect 37998 23042 38050 23054
rect 37998 22978 38050 22990
rect 39678 23042 39730 23054
rect 39678 22978 39730 22990
rect 5294 22930 5346 22942
rect 30718 22930 30770 22942
rect 12114 22878 12126 22930
rect 12178 22927 12190 22930
rect 12674 22927 12686 22930
rect 12178 22881 12686 22927
rect 12178 22878 12190 22881
rect 12674 22878 12686 22881
rect 12738 22878 12750 22930
rect 5294 22866 5346 22878
rect 30718 22866 30770 22878
rect 30942 22930 30994 22942
rect 36878 22930 36930 22942
rect 34962 22878 34974 22930
rect 35026 22878 35038 22930
rect 30942 22866 30994 22878
rect 36878 22866 36930 22878
rect 43598 22930 43650 22942
rect 43598 22866 43650 22878
rect 43934 22930 43986 22942
rect 43934 22866 43986 22878
rect 1344 22762 48720 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48720 22762
rect 1344 22676 48720 22710
rect 9998 22594 10050 22606
rect 9998 22530 10050 22542
rect 46846 22594 46898 22606
rect 46846 22530 46898 22542
rect 47182 22594 47234 22606
rect 47182 22530 47234 22542
rect 6302 22482 6354 22494
rect 6302 22418 6354 22430
rect 10670 22482 10722 22494
rect 12910 22482 12962 22494
rect 11666 22430 11678 22482
rect 11730 22430 11742 22482
rect 10670 22418 10722 22430
rect 12910 22418 12962 22430
rect 13582 22482 13634 22494
rect 13582 22418 13634 22430
rect 17390 22482 17442 22494
rect 23438 22482 23490 22494
rect 17714 22430 17726 22482
rect 17778 22430 17790 22482
rect 17390 22418 17442 22430
rect 23438 22418 23490 22430
rect 24222 22482 24274 22494
rect 24222 22418 24274 22430
rect 25230 22482 25282 22494
rect 37550 22482 37602 22494
rect 43262 22482 43314 22494
rect 27906 22430 27918 22482
rect 27970 22430 27982 22482
rect 35186 22430 35198 22482
rect 35250 22430 35262 22482
rect 36194 22430 36206 22482
rect 36258 22430 36270 22482
rect 42802 22430 42814 22482
rect 42866 22430 42878 22482
rect 25230 22418 25282 22430
rect 37550 22418 37602 22430
rect 43262 22418 43314 22430
rect 44942 22482 44994 22494
rect 44942 22418 44994 22430
rect 45390 22482 45442 22494
rect 45390 22418 45442 22430
rect 2606 22370 2658 22382
rect 2606 22306 2658 22318
rect 4958 22370 5010 22382
rect 12462 22370 12514 22382
rect 21982 22370 22034 22382
rect 24782 22370 24834 22382
rect 6514 22318 6526 22370
rect 6578 22318 6590 22370
rect 7298 22318 7310 22370
rect 7362 22318 7374 22370
rect 11554 22318 11566 22370
rect 11618 22318 11630 22370
rect 16930 22318 16942 22370
rect 16994 22318 17006 22370
rect 20066 22318 20078 22370
rect 20130 22318 20142 22370
rect 20850 22318 20862 22370
rect 20914 22318 20926 22370
rect 22978 22318 22990 22370
rect 23042 22318 23054 22370
rect 4958 22306 5010 22318
rect 12462 22306 12514 22318
rect 21982 22306 22034 22318
rect 24782 22306 24834 22318
rect 27470 22370 27522 22382
rect 29486 22370 29538 22382
rect 28242 22318 28254 22370
rect 28306 22318 28318 22370
rect 27470 22306 27522 22318
rect 29486 22306 29538 22318
rect 29710 22370 29762 22382
rect 29710 22306 29762 22318
rect 30158 22370 30210 22382
rect 37774 22370 37826 22382
rect 30594 22318 30606 22370
rect 30658 22318 30670 22370
rect 31490 22318 31502 22370
rect 31554 22318 31566 22370
rect 31826 22318 31838 22370
rect 31890 22318 31902 22370
rect 33954 22318 33966 22370
rect 34018 22318 34030 22370
rect 34850 22318 34862 22370
rect 34914 22318 34926 22370
rect 35858 22318 35870 22370
rect 35922 22318 35934 22370
rect 30158 22306 30210 22318
rect 37774 22306 37826 22318
rect 37998 22370 38050 22382
rect 43710 22370 43762 22382
rect 39666 22318 39678 22370
rect 39730 22318 39742 22370
rect 40338 22318 40350 22370
rect 40402 22318 40414 22370
rect 37998 22306 38050 22318
rect 43710 22306 43762 22318
rect 2270 22258 2322 22270
rect 10110 22258 10162 22270
rect 9650 22206 9662 22258
rect 9714 22206 9726 22258
rect 2270 22194 2322 22206
rect 10110 22194 10162 22206
rect 11006 22258 11058 22270
rect 29150 22258 29202 22270
rect 12114 22206 12126 22258
rect 12178 22206 12190 22258
rect 11006 22194 11058 22206
rect 29150 22194 29202 22206
rect 29598 22258 29650 22270
rect 32174 22258 32226 22270
rect 34414 22258 34466 22270
rect 30706 22206 30718 22258
rect 30770 22206 30782 22258
rect 33058 22206 33070 22258
rect 33122 22206 33134 22258
rect 33730 22206 33742 22258
rect 33794 22206 33806 22258
rect 29598 22194 29650 22206
rect 32174 22194 32226 22206
rect 34414 22194 34466 22206
rect 44046 22258 44098 22270
rect 47394 22206 47406 22258
rect 47458 22206 47470 22258
rect 47954 22206 47966 22258
rect 48018 22206 48030 22258
rect 44046 22194 44098 22206
rect 5742 22146 5794 22158
rect 5742 22082 5794 22094
rect 14030 22146 14082 22158
rect 14030 22082 14082 22094
rect 22542 22146 22594 22158
rect 22542 22082 22594 22094
rect 25790 22146 25842 22158
rect 32734 22146 32786 22158
rect 27122 22094 27134 22146
rect 27186 22094 27198 22146
rect 25790 22082 25842 22094
rect 32734 22082 32786 22094
rect 37102 22146 37154 22158
rect 37102 22082 37154 22094
rect 37214 22146 37266 22158
rect 37214 22082 37266 22094
rect 37326 22146 37378 22158
rect 37326 22082 37378 22094
rect 39006 22146 39058 22158
rect 39006 22082 39058 22094
rect 39454 22146 39506 22158
rect 39454 22082 39506 22094
rect 1344 21978 48720 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48720 21978
rect 1344 21892 48720 21926
rect 9102 21810 9154 21822
rect 23438 21810 23490 21822
rect 10658 21758 10670 21810
rect 10722 21758 10734 21810
rect 16482 21758 16494 21810
rect 16546 21758 16558 21810
rect 9102 21746 9154 21758
rect 23438 21746 23490 21758
rect 27806 21810 27858 21822
rect 27806 21746 27858 21758
rect 31726 21810 31778 21822
rect 31726 21746 31778 21758
rect 37102 21810 37154 21822
rect 47618 21758 47630 21810
rect 47682 21758 47694 21810
rect 37102 21746 37154 21758
rect 18174 21698 18226 21710
rect 6402 21646 6414 21698
rect 6466 21646 6478 21698
rect 9650 21646 9662 21698
rect 9714 21646 9726 21698
rect 10322 21646 10334 21698
rect 10386 21646 10398 21698
rect 18174 21634 18226 21646
rect 19070 21698 19122 21710
rect 19070 21634 19122 21646
rect 21086 21698 21138 21710
rect 21086 21634 21138 21646
rect 22206 21698 22258 21710
rect 22206 21634 22258 21646
rect 23774 21698 23826 21710
rect 23774 21634 23826 21646
rect 25454 21698 25506 21710
rect 25454 21634 25506 21646
rect 26014 21698 26066 21710
rect 27582 21698 27634 21710
rect 26786 21646 26798 21698
rect 26850 21646 26862 21698
rect 26014 21634 26066 21646
rect 27582 21634 27634 21646
rect 28254 21698 28306 21710
rect 28254 21634 28306 21646
rect 29710 21698 29762 21710
rect 29710 21634 29762 21646
rect 32286 21698 32338 21710
rect 37774 21698 37826 21710
rect 33170 21646 33182 21698
rect 33234 21646 33246 21698
rect 32286 21634 32338 21646
rect 37774 21634 37826 21646
rect 37998 21698 38050 21710
rect 37998 21634 38050 21646
rect 38334 21698 38386 21710
rect 38334 21634 38386 21646
rect 39454 21698 39506 21710
rect 39454 21634 39506 21646
rect 40126 21698 40178 21710
rect 40126 21634 40178 21646
rect 47966 21698 48018 21710
rect 47966 21634 48018 21646
rect 5630 21586 5682 21598
rect 16830 21586 16882 21598
rect 19630 21586 19682 21598
rect 1922 21534 1934 21586
rect 1986 21534 1998 21586
rect 2482 21534 2494 21586
rect 2546 21534 2558 21586
rect 4834 21534 4846 21586
rect 4898 21534 4910 21586
rect 6290 21534 6302 21586
rect 6354 21534 6366 21586
rect 9762 21534 9774 21586
rect 9826 21534 9838 21586
rect 10770 21534 10782 21586
rect 10834 21534 10846 21586
rect 11330 21534 11342 21586
rect 11394 21534 11406 21586
rect 12226 21534 12238 21586
rect 12290 21534 12302 21586
rect 13122 21534 13134 21586
rect 13186 21534 13198 21586
rect 13570 21534 13582 21586
rect 13634 21534 13646 21586
rect 17714 21534 17726 21586
rect 17778 21534 17790 21586
rect 5630 21522 5682 21534
rect 16830 21522 16882 21534
rect 19630 21522 19682 21534
rect 20190 21586 20242 21598
rect 20190 21522 20242 21534
rect 22542 21586 22594 21598
rect 22542 21522 22594 21534
rect 24334 21586 24386 21598
rect 28030 21586 28082 21598
rect 25778 21534 25790 21586
rect 25842 21534 25854 21586
rect 26674 21534 26686 21586
rect 26738 21534 26750 21586
rect 24334 21522 24386 21534
rect 28030 21522 28082 21534
rect 28702 21586 28754 21598
rect 28702 21522 28754 21534
rect 29262 21586 29314 21598
rect 29262 21522 29314 21534
rect 29598 21586 29650 21598
rect 29598 21522 29650 21534
rect 31838 21586 31890 21598
rect 31838 21522 31890 21534
rect 32174 21586 32226 21598
rect 36094 21586 36146 21598
rect 33282 21534 33294 21586
rect 33346 21534 33358 21586
rect 34066 21534 34078 21586
rect 34130 21534 34142 21586
rect 34514 21534 34526 21586
rect 34578 21534 34590 21586
rect 35746 21534 35758 21586
rect 35810 21534 35822 21586
rect 32174 21522 32226 21534
rect 36094 21522 36146 21534
rect 36318 21586 36370 21598
rect 36318 21522 36370 21534
rect 37438 21586 37490 21598
rect 37438 21522 37490 21534
rect 38446 21586 38498 21598
rect 38446 21522 38498 21534
rect 38670 21586 38722 21598
rect 42366 21586 42418 21598
rect 41122 21534 41134 21586
rect 41186 21534 41198 21586
rect 42802 21534 42814 21586
rect 42866 21534 42878 21586
rect 44482 21534 44494 21586
rect 44546 21534 44558 21586
rect 45154 21534 45166 21586
rect 45218 21534 45230 21586
rect 48178 21534 48190 21586
rect 48242 21534 48254 21586
rect 38670 21522 38722 21534
rect 42366 21522 42418 21534
rect 6974 21474 7026 21486
rect 6974 21410 7026 21422
rect 12686 21474 12738 21486
rect 18510 21474 18562 21486
rect 16034 21422 16046 21474
rect 16098 21422 16110 21474
rect 12686 21410 12738 21422
rect 18510 21410 18562 21422
rect 20526 21474 20578 21486
rect 20526 21410 20578 21422
rect 22878 21474 22930 21486
rect 28366 21474 28418 21486
rect 39342 21474 39394 21486
rect 26562 21422 26574 21474
rect 26626 21422 26638 21474
rect 33618 21422 33630 21474
rect 33682 21422 33694 21474
rect 40114 21422 40126 21474
rect 40178 21422 40190 21474
rect 43026 21422 43038 21474
rect 43090 21422 43102 21474
rect 22878 21410 22930 21422
rect 28366 21410 28418 21422
rect 39342 21410 39394 21422
rect 5294 21362 5346 21374
rect 5294 21298 5346 21310
rect 29710 21362 29762 21374
rect 29710 21298 29762 21310
rect 31726 21362 31778 21374
rect 31726 21298 31778 21310
rect 32286 21362 32338 21374
rect 32286 21298 32338 21310
rect 37214 21362 37266 21374
rect 37214 21298 37266 21310
rect 38782 21362 38834 21374
rect 38782 21298 38834 21310
rect 39230 21362 39282 21374
rect 39230 21298 39282 21310
rect 39902 21362 39954 21374
rect 43586 21310 43598 21362
rect 43650 21310 43662 21362
rect 39902 21298 39954 21310
rect 1344 21194 48720 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48720 21194
rect 1344 21108 48720 21142
rect 6414 21026 6466 21038
rect 6414 20962 6466 20974
rect 13582 21026 13634 21038
rect 13582 20962 13634 20974
rect 14254 21026 14306 21038
rect 14254 20962 14306 20974
rect 14366 21026 14418 21038
rect 14366 20962 14418 20974
rect 15150 21026 15202 21038
rect 25902 21026 25954 21038
rect 25330 20974 25342 21026
rect 25394 20974 25406 21026
rect 15150 20962 15202 20974
rect 25902 20962 25954 20974
rect 26126 21026 26178 21038
rect 26126 20962 26178 20974
rect 34190 21026 34242 21038
rect 34190 20962 34242 20974
rect 43486 21026 43538 21038
rect 43486 20962 43538 20974
rect 5070 20914 5122 20926
rect 5070 20850 5122 20862
rect 8990 20914 9042 20926
rect 8990 20850 9042 20862
rect 9326 20914 9378 20926
rect 9326 20850 9378 20862
rect 15262 20914 15314 20926
rect 20638 20914 20690 20926
rect 19506 20862 19518 20914
rect 19570 20862 19582 20914
rect 15262 20850 15314 20862
rect 20638 20850 20690 20862
rect 22094 20914 22146 20926
rect 28254 20914 28306 20926
rect 23986 20862 23998 20914
rect 24050 20862 24062 20914
rect 26674 20862 26686 20914
rect 26738 20862 26750 20914
rect 22094 20850 22146 20862
rect 28254 20850 28306 20862
rect 31054 20914 31106 20926
rect 31054 20850 31106 20862
rect 31950 20914 32002 20926
rect 31950 20850 32002 20862
rect 36990 20914 37042 20926
rect 44046 20914 44098 20926
rect 41570 20862 41582 20914
rect 41634 20862 41646 20914
rect 36990 20850 37042 20862
rect 44046 20850 44098 20862
rect 44942 20914 44994 20926
rect 48290 20862 48302 20914
rect 48354 20862 48366 20914
rect 44942 20850 44994 20862
rect 2942 20802 2994 20814
rect 2942 20738 2994 20750
rect 9998 20802 10050 20814
rect 13806 20802 13858 20814
rect 10546 20750 10558 20802
rect 10610 20750 10622 20802
rect 11554 20750 11566 20802
rect 11618 20750 11630 20802
rect 12114 20750 12126 20802
rect 12178 20750 12190 20802
rect 9998 20738 10050 20750
rect 13806 20738 13858 20750
rect 14814 20802 14866 20814
rect 22318 20802 22370 20814
rect 24782 20802 24834 20814
rect 26574 20802 26626 20814
rect 18050 20750 18062 20802
rect 18114 20750 18126 20802
rect 22978 20750 22990 20802
rect 23042 20750 23054 20802
rect 25554 20750 25566 20802
rect 25618 20750 25630 20802
rect 26450 20750 26462 20802
rect 26514 20750 26526 20802
rect 14814 20738 14866 20750
rect 22318 20738 22370 20750
rect 24782 20738 24834 20750
rect 26574 20738 26626 20750
rect 27246 20802 27298 20814
rect 27246 20738 27298 20750
rect 27806 20802 27858 20814
rect 27806 20738 27858 20750
rect 29822 20802 29874 20814
rect 30270 20802 30322 20814
rect 30830 20802 30882 20814
rect 30034 20750 30046 20802
rect 30098 20750 30110 20802
rect 30482 20750 30494 20802
rect 30546 20750 30558 20802
rect 29822 20738 29874 20750
rect 30270 20738 30322 20750
rect 30830 20738 30882 20750
rect 31166 20802 31218 20814
rect 31166 20738 31218 20750
rect 33406 20802 33458 20814
rect 33406 20738 33458 20750
rect 33742 20802 33794 20814
rect 33742 20738 33794 20750
rect 34862 20802 34914 20814
rect 43822 20802 43874 20814
rect 37314 20750 37326 20802
rect 37378 20750 37390 20802
rect 37874 20750 37886 20802
rect 37938 20750 37950 20802
rect 39218 20750 39230 20802
rect 39282 20750 39294 20802
rect 40114 20750 40126 20802
rect 40178 20750 40190 20802
rect 42914 20750 42926 20802
rect 42978 20750 42990 20802
rect 45154 20750 45166 20802
rect 45218 20750 45230 20802
rect 45938 20750 45950 20802
rect 46002 20750 46014 20802
rect 34862 20738 34914 20750
rect 43822 20738 43874 20750
rect 2606 20690 2658 20702
rect 9662 20690 9714 20702
rect 14142 20690 14194 20702
rect 6626 20638 6638 20690
rect 6690 20638 6702 20690
rect 6962 20638 6974 20690
rect 7026 20638 7038 20690
rect 10770 20638 10782 20690
rect 10834 20638 10846 20690
rect 11106 20638 11118 20690
rect 11170 20638 11182 20690
rect 2606 20626 2658 20638
rect 9662 20626 9714 20638
rect 14142 20626 14194 20638
rect 23438 20690 23490 20702
rect 31502 20690 31554 20702
rect 24994 20638 25006 20690
rect 25058 20638 25070 20690
rect 23438 20626 23490 20638
rect 31502 20626 31554 20638
rect 32286 20690 32338 20702
rect 32286 20626 32338 20638
rect 32398 20690 32450 20702
rect 32398 20626 32450 20638
rect 32622 20690 32674 20702
rect 32622 20626 32674 20638
rect 32846 20690 32898 20702
rect 32846 20626 32898 20638
rect 33518 20690 33570 20702
rect 33518 20626 33570 20638
rect 34526 20690 34578 20702
rect 34526 20626 34578 20638
rect 34974 20690 35026 20702
rect 34974 20626 35026 20638
rect 38446 20690 38498 20702
rect 38446 20626 38498 20638
rect 6078 20578 6130 20590
rect 6078 20514 6130 20526
rect 8094 20578 8146 20590
rect 8094 20514 8146 20526
rect 8430 20578 8482 20590
rect 17054 20578 17106 20590
rect 11442 20526 11454 20578
rect 11506 20526 11518 20578
rect 8430 20514 8482 20526
rect 17054 20514 17106 20526
rect 21534 20578 21586 20590
rect 21534 20514 21586 20526
rect 22430 20578 22482 20590
rect 22430 20514 22482 20526
rect 22654 20578 22706 20590
rect 22654 20514 22706 20526
rect 24446 20578 24498 20590
rect 26798 20578 26850 20590
rect 25218 20526 25230 20578
rect 25282 20526 25294 20578
rect 24446 20514 24498 20526
rect 26798 20514 26850 20526
rect 30606 20578 30658 20590
rect 30606 20514 30658 20526
rect 32958 20578 33010 20590
rect 32958 20514 33010 20526
rect 33182 20578 33234 20590
rect 33182 20514 33234 20526
rect 34302 20578 34354 20590
rect 34302 20514 34354 20526
rect 35198 20578 35250 20590
rect 37986 20526 37998 20578
rect 38050 20526 38062 20578
rect 35198 20514 35250 20526
rect 1344 20410 48720 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48720 20410
rect 1344 20324 48720 20358
rect 27246 20242 27298 20254
rect 39118 20242 39170 20254
rect 25890 20190 25902 20242
rect 25954 20190 25966 20242
rect 28690 20190 28702 20242
rect 28754 20190 28766 20242
rect 43810 20190 43822 20242
rect 43874 20239 43886 20242
rect 43874 20193 43983 20239
rect 43874 20190 43886 20193
rect 27246 20178 27298 20190
rect 39118 20178 39170 20190
rect 5630 20130 5682 20142
rect 13918 20130 13970 20142
rect 8978 20078 8990 20130
rect 9042 20078 9054 20130
rect 5630 20066 5682 20078
rect 13918 20066 13970 20078
rect 14366 20130 14418 20142
rect 14366 20066 14418 20078
rect 15150 20130 15202 20142
rect 27806 20130 27858 20142
rect 23874 20078 23886 20130
rect 23938 20078 23950 20130
rect 25330 20078 25342 20130
rect 25394 20078 25406 20130
rect 26786 20078 26798 20130
rect 26850 20078 26862 20130
rect 15150 20066 15202 20078
rect 27806 20066 27858 20078
rect 29710 20130 29762 20142
rect 29710 20066 29762 20078
rect 29822 20130 29874 20142
rect 29822 20066 29874 20078
rect 29934 20130 29986 20142
rect 29934 20066 29986 20078
rect 30382 20130 30434 20142
rect 30382 20066 30434 20078
rect 32174 20130 32226 20142
rect 32174 20066 32226 20078
rect 32398 20130 32450 20142
rect 35522 20078 35534 20130
rect 35586 20078 35598 20130
rect 36418 20078 36430 20130
rect 36482 20078 36494 20130
rect 39666 20078 39678 20130
rect 39730 20078 39742 20130
rect 40002 20078 40014 20130
rect 40066 20078 40078 20130
rect 43937 20127 43983 20193
rect 44146 20127 44158 20130
rect 43937 20081 44158 20127
rect 44146 20078 44158 20081
rect 44210 20078 44222 20130
rect 32398 20066 32450 20078
rect 10446 20018 10498 20030
rect 14702 20018 14754 20030
rect 5394 19966 5406 20018
rect 5458 19966 5470 20018
rect 5842 19966 5854 20018
rect 5906 19966 5918 20018
rect 6514 19966 6526 20018
rect 6578 19966 6590 20018
rect 9986 19966 9998 20018
rect 10050 19966 10062 20018
rect 13346 19966 13358 20018
rect 13410 19966 13422 20018
rect 10446 19954 10498 19966
rect 14702 19954 14754 19966
rect 16830 20018 16882 20030
rect 27358 20018 27410 20030
rect 18162 19966 18174 20018
rect 18226 19966 18238 20018
rect 21298 19966 21310 20018
rect 21362 19966 21374 20018
rect 22530 19966 22542 20018
rect 22594 19966 22606 20018
rect 23426 19966 23438 20018
rect 23490 19966 23502 20018
rect 25890 19966 25902 20018
rect 25954 19966 25966 20018
rect 26898 19966 26910 20018
rect 26962 19966 26974 20018
rect 16830 19954 16882 19966
rect 27358 19954 27410 19966
rect 28254 20018 28306 20030
rect 28254 19954 28306 19966
rect 29038 20018 29090 20030
rect 29038 19954 29090 19966
rect 29262 20018 29314 20030
rect 29262 19954 29314 19966
rect 30270 20018 30322 20030
rect 30270 19954 30322 19966
rect 32510 20018 32562 20030
rect 34414 20018 34466 20030
rect 46062 20018 46114 20030
rect 33394 19966 33406 20018
rect 33458 19966 33470 20018
rect 32510 19954 32562 19966
rect 33730 19965 33742 20017
rect 33794 19965 33806 20017
rect 36194 19966 36206 20018
rect 36258 19966 36270 20018
rect 38098 19966 38110 20018
rect 38162 19966 38174 20018
rect 42914 19966 42926 20018
rect 42978 19966 42990 20018
rect 44258 19966 44270 20018
rect 44322 19966 44334 20018
rect 45378 19966 45390 20018
rect 45442 19966 45454 20018
rect 46274 19966 46286 20018
rect 46338 19966 46350 20018
rect 34414 19954 34466 19966
rect 46062 19954 46114 19966
rect 16270 19906 16322 19918
rect 10994 19854 11006 19906
rect 11058 19854 11070 19906
rect 16270 19842 16322 19854
rect 17614 19906 17666 19918
rect 38558 19906 38610 19918
rect 18834 19854 18846 19906
rect 18898 19854 18910 19906
rect 20962 19854 20974 19906
rect 21026 19854 21038 19906
rect 33618 19854 33630 19906
rect 33682 19854 33694 19906
rect 36418 19854 36430 19906
rect 36482 19854 36494 19906
rect 41906 19854 41918 19906
rect 41970 19854 41982 19906
rect 17614 19842 17666 19854
rect 38558 19842 38610 19854
rect 39454 19794 39506 19806
rect 24546 19742 24558 19794
rect 24610 19742 24622 19794
rect 44594 19742 44606 19794
rect 44658 19742 44670 19794
rect 39454 19730 39506 19742
rect 1344 19626 48720 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48720 19626
rect 1344 19540 48720 19574
rect 43150 19458 43202 19470
rect 48078 19458 48130 19470
rect 28018 19406 28030 19458
rect 28082 19406 28094 19458
rect 37202 19406 37214 19458
rect 37266 19406 37278 19458
rect 45490 19406 45502 19458
rect 45554 19406 45566 19458
rect 43150 19394 43202 19406
rect 48078 19394 48130 19406
rect 5742 19346 5794 19358
rect 5742 19282 5794 19294
rect 7310 19346 7362 19358
rect 7310 19282 7362 19294
rect 8430 19346 8482 19358
rect 8430 19282 8482 19294
rect 8990 19346 9042 19358
rect 20750 19346 20802 19358
rect 26014 19346 26066 19358
rect 28590 19346 28642 19358
rect 37662 19346 37714 19358
rect 42590 19346 42642 19358
rect 10546 19294 10558 19346
rect 10610 19294 10622 19346
rect 17266 19294 17278 19346
rect 17330 19294 17342 19346
rect 19954 19294 19966 19346
rect 20018 19294 20030 19346
rect 23986 19294 23998 19346
rect 24050 19294 24062 19346
rect 26786 19294 26798 19346
rect 26850 19294 26862 19346
rect 29586 19294 29598 19346
rect 29650 19294 29662 19346
rect 33394 19294 33406 19346
rect 33458 19294 33470 19346
rect 35970 19294 35982 19346
rect 36034 19294 36046 19346
rect 39330 19294 39342 19346
rect 39394 19294 39406 19346
rect 41794 19294 41806 19346
rect 41858 19294 41870 19346
rect 8990 19282 9042 19294
rect 20750 19282 20802 19294
rect 26014 19282 26066 19294
rect 28590 19282 28642 19294
rect 37662 19282 37714 19294
rect 42590 19282 42642 19294
rect 43486 19346 43538 19358
rect 45266 19294 45278 19346
rect 45330 19294 45342 19346
rect 43486 19282 43538 19294
rect 6862 19234 6914 19246
rect 21422 19234 21474 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 2258 19182 2270 19234
rect 2322 19182 2334 19234
rect 9986 19182 9998 19234
rect 10050 19182 10062 19234
rect 12786 19182 12798 19234
rect 12850 19182 12862 19234
rect 13682 19182 13694 19234
rect 13746 19182 13758 19234
rect 14354 19182 14366 19234
rect 14418 19182 14430 19234
rect 18050 19182 18062 19234
rect 18114 19182 18126 19234
rect 6862 19170 6914 19182
rect 21422 19170 21474 19182
rect 21982 19234 22034 19246
rect 28366 19234 28418 19246
rect 34526 19234 34578 19246
rect 22418 19182 22430 19234
rect 22482 19182 22494 19234
rect 24098 19182 24110 19234
rect 24162 19182 24174 19234
rect 26674 19182 26686 19234
rect 26738 19182 26750 19234
rect 29138 19182 29150 19234
rect 29202 19182 29214 19234
rect 30818 19182 30830 19234
rect 30882 19182 30894 19234
rect 21982 19170 22034 19182
rect 28366 19170 28418 19182
rect 34526 19170 34578 19182
rect 36430 19234 36482 19246
rect 42814 19234 42866 19246
rect 37090 19182 37102 19234
rect 37154 19182 37166 19234
rect 37538 19182 37550 19234
rect 37602 19182 37614 19234
rect 40338 19182 40350 19234
rect 40402 19182 40414 19234
rect 41010 19182 41022 19234
rect 41074 19182 41086 19234
rect 36430 19170 36482 19182
rect 42814 19170 42866 19182
rect 43710 19234 43762 19246
rect 47742 19234 47794 19246
rect 45042 19182 45054 19234
rect 45106 19182 45118 19234
rect 46274 19182 46286 19234
rect 46338 19182 46350 19234
rect 43710 19170 43762 19182
rect 47742 19170 47794 19182
rect 6302 19122 6354 19134
rect 6302 19058 6354 19070
rect 9438 19122 9490 19134
rect 9438 19058 9490 19070
rect 9550 19122 9602 19134
rect 27358 19122 27410 19134
rect 15138 19070 15150 19122
rect 15202 19070 15214 19122
rect 22978 19070 22990 19122
rect 23042 19070 23054 19122
rect 24210 19070 24222 19122
rect 24274 19070 24286 19122
rect 9550 19058 9602 19070
rect 27358 19058 27410 19070
rect 27694 19122 27746 19134
rect 31950 19122 32002 19134
rect 29362 19070 29374 19122
rect 29426 19070 29438 19122
rect 27694 19058 27746 19070
rect 31950 19058 32002 19070
rect 33966 19122 34018 19134
rect 33966 19058 34018 19070
rect 37774 19122 37826 19134
rect 37774 19058 37826 19070
rect 45838 19122 45890 19134
rect 47170 19070 47182 19122
rect 47234 19070 47246 19122
rect 47394 19070 47406 19122
rect 47458 19070 47470 19122
rect 45838 19058 45890 19070
rect 9214 19010 9266 19022
rect 4722 18958 4734 19010
rect 4786 18958 4798 19010
rect 9214 18946 9266 18958
rect 9326 19010 9378 19022
rect 34974 19010 35026 19022
rect 13458 18958 13470 19010
rect 13522 18958 13534 19010
rect 35298 18958 35310 19010
rect 35362 18958 35374 19010
rect 44034 18958 44046 19010
rect 44098 18958 44110 19010
rect 9326 18946 9378 18958
rect 34974 18946 35026 18958
rect 1344 18842 48720 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48720 18842
rect 1344 18756 48720 18790
rect 2270 18674 2322 18686
rect 2270 18610 2322 18622
rect 14926 18674 14978 18686
rect 14926 18610 14978 18622
rect 25566 18674 25618 18686
rect 25566 18610 25618 18622
rect 27694 18674 27746 18686
rect 27694 18610 27746 18622
rect 29262 18674 29314 18686
rect 29262 18610 29314 18622
rect 29486 18674 29538 18686
rect 29486 18610 29538 18622
rect 32510 18674 32562 18686
rect 43598 18674 43650 18686
rect 34066 18622 34078 18674
rect 34130 18622 34142 18674
rect 37426 18622 37438 18674
rect 37490 18622 37502 18674
rect 32510 18610 32562 18622
rect 43598 18610 43650 18622
rect 6750 18562 6802 18574
rect 5170 18510 5182 18562
rect 5234 18510 5246 18562
rect 6750 18498 6802 18510
rect 19294 18562 19346 18574
rect 28590 18562 28642 18574
rect 25218 18510 25230 18562
rect 25282 18510 25294 18562
rect 19294 18498 19346 18510
rect 28590 18498 28642 18510
rect 29038 18562 29090 18574
rect 29038 18498 29090 18510
rect 29598 18562 29650 18574
rect 36990 18562 37042 18574
rect 42814 18562 42866 18574
rect 34290 18510 34302 18562
rect 34354 18510 34366 18562
rect 36642 18510 36654 18562
rect 36706 18510 36718 18562
rect 41010 18510 41022 18562
rect 41074 18510 41086 18562
rect 29598 18498 29650 18510
rect 36990 18498 37042 18510
rect 42814 18498 42866 18510
rect 44942 18562 44994 18574
rect 44942 18498 44994 18510
rect 2606 18450 2658 18462
rect 2606 18386 2658 18398
rect 4062 18450 4114 18462
rect 4062 18386 4114 18398
rect 4398 18450 4450 18462
rect 6414 18450 6466 18462
rect 10334 18450 10386 18462
rect 4834 18398 4846 18450
rect 4898 18398 4910 18450
rect 9986 18398 9998 18450
rect 10050 18398 10062 18450
rect 4398 18386 4450 18398
rect 6414 18386 6466 18398
rect 10334 18386 10386 18398
rect 10670 18450 10722 18462
rect 10670 18386 10722 18398
rect 10894 18450 10946 18462
rect 10894 18386 10946 18398
rect 11454 18450 11506 18462
rect 12350 18450 12402 18462
rect 11778 18398 11790 18450
rect 11842 18398 11854 18450
rect 11454 18386 11506 18398
rect 12350 18386 12402 18398
rect 12462 18450 12514 18462
rect 12462 18386 12514 18398
rect 14254 18450 14306 18462
rect 14254 18386 14306 18398
rect 14702 18450 14754 18462
rect 14702 18386 14754 18398
rect 15262 18450 15314 18462
rect 15262 18386 15314 18398
rect 15710 18450 15762 18462
rect 19630 18450 19682 18462
rect 17938 18398 17950 18450
rect 18002 18398 18014 18450
rect 18274 18398 18286 18450
rect 18338 18398 18350 18450
rect 15710 18386 15762 18398
rect 19630 18386 19682 18398
rect 20414 18450 20466 18462
rect 20414 18386 20466 18398
rect 24558 18450 24610 18462
rect 26910 18450 26962 18462
rect 30494 18450 30546 18462
rect 31950 18450 32002 18462
rect 35534 18450 35586 18462
rect 37998 18450 38050 18462
rect 26450 18398 26462 18450
rect 26514 18398 26526 18450
rect 26674 18398 26686 18450
rect 26738 18398 26750 18450
rect 28802 18398 28814 18450
rect 28866 18398 28878 18450
rect 30930 18398 30942 18450
rect 30994 18398 31006 18450
rect 33170 18398 33182 18450
rect 33234 18398 33246 18450
rect 33394 18398 33406 18450
rect 33458 18398 33470 18450
rect 34178 18398 34190 18450
rect 34242 18398 34254 18450
rect 36418 18398 36430 18450
rect 36482 18398 36494 18450
rect 37202 18398 37214 18450
rect 37266 18398 37278 18450
rect 37538 18398 37550 18450
rect 37602 18398 37614 18450
rect 24558 18386 24610 18398
rect 26910 18386 26962 18398
rect 30494 18386 30546 18398
rect 31950 18386 32002 18398
rect 35534 18386 35586 18398
rect 37998 18386 38050 18398
rect 38222 18450 38274 18462
rect 38222 18386 38274 18398
rect 38334 18450 38386 18462
rect 38334 18386 38386 18398
rect 38670 18450 38722 18462
rect 38670 18386 38722 18398
rect 39006 18450 39058 18462
rect 39006 18386 39058 18398
rect 39230 18450 39282 18462
rect 39230 18386 39282 18398
rect 39454 18450 39506 18462
rect 39454 18386 39506 18398
rect 39678 18450 39730 18462
rect 41918 18450 41970 18462
rect 40898 18398 40910 18450
rect 40962 18398 40974 18450
rect 43026 18398 43038 18450
rect 43090 18398 43102 18450
rect 44706 18398 44718 18450
rect 44770 18398 44782 18450
rect 45154 18398 45166 18450
rect 45218 18398 45230 18450
rect 45826 18398 45838 18450
rect 45890 18398 45902 18450
rect 39678 18386 39730 18398
rect 41918 18386 41970 18398
rect 9774 18338 9826 18350
rect 9774 18274 9826 18286
rect 10782 18338 10834 18350
rect 10782 18274 10834 18286
rect 12238 18338 12290 18350
rect 12238 18274 12290 18286
rect 13134 18338 13186 18350
rect 13134 18274 13186 18286
rect 13806 18338 13858 18350
rect 20862 18338 20914 18350
rect 18386 18286 18398 18338
rect 18450 18286 18462 18338
rect 13806 18274 13858 18286
rect 20862 18274 20914 18286
rect 22094 18338 22146 18350
rect 22094 18274 22146 18286
rect 23774 18338 23826 18350
rect 35086 18338 35138 18350
rect 24098 18286 24110 18338
rect 24162 18286 24174 18338
rect 31266 18286 31278 18338
rect 31330 18286 31342 18338
rect 23774 18274 23826 18286
rect 35086 18274 35138 18286
rect 35982 18338 36034 18350
rect 35982 18274 36034 18286
rect 40014 18338 40066 18350
rect 44046 18338 44098 18350
rect 42354 18286 42366 18338
rect 42418 18286 42430 18338
rect 48290 18286 48302 18338
rect 48354 18286 48366 18338
rect 40014 18274 40066 18286
rect 44046 18274 44098 18286
rect 10446 18226 10498 18238
rect 10446 18162 10498 18174
rect 12014 18226 12066 18238
rect 12014 18162 12066 18174
rect 14030 18226 14082 18238
rect 14030 18162 14082 18174
rect 17726 18226 17778 18238
rect 17726 18162 17778 18174
rect 28702 18226 28754 18238
rect 28702 18162 28754 18174
rect 37438 18226 37490 18238
rect 37438 18162 37490 18174
rect 41022 18226 41074 18238
rect 41022 18162 41074 18174
rect 1344 18058 48720 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48720 18058
rect 1344 17972 48720 18006
rect 4174 17890 4226 17902
rect 4174 17826 4226 17838
rect 6190 17890 6242 17902
rect 6190 17826 6242 17838
rect 9102 17890 9154 17902
rect 9102 17826 9154 17838
rect 11790 17890 11842 17902
rect 11790 17826 11842 17838
rect 16046 17890 16098 17902
rect 16046 17826 16098 17838
rect 17950 17890 18002 17902
rect 17950 17826 18002 17838
rect 18958 17890 19010 17902
rect 18958 17826 19010 17838
rect 45726 17890 45778 17902
rect 45726 17826 45778 17838
rect 46062 17890 46114 17902
rect 46062 17826 46114 17838
rect 8542 17778 8594 17790
rect 8542 17714 8594 17726
rect 11118 17778 11170 17790
rect 11118 17714 11170 17726
rect 12126 17778 12178 17790
rect 12126 17714 12178 17726
rect 12910 17778 12962 17790
rect 12910 17714 12962 17726
rect 13582 17778 13634 17790
rect 13582 17714 13634 17726
rect 14702 17778 14754 17790
rect 14702 17714 14754 17726
rect 19182 17778 19234 17790
rect 19182 17714 19234 17726
rect 19406 17778 19458 17790
rect 32734 17778 32786 17790
rect 23650 17726 23662 17778
rect 23714 17726 23726 17778
rect 29922 17726 29934 17778
rect 29986 17726 29998 17778
rect 32162 17726 32174 17778
rect 32226 17726 32238 17778
rect 19406 17714 19458 17726
rect 32734 17714 32786 17726
rect 34750 17778 34802 17790
rect 34750 17714 34802 17726
rect 35534 17778 35586 17790
rect 39902 17778 39954 17790
rect 45054 17778 45106 17790
rect 37202 17726 37214 17778
rect 37266 17726 37278 17778
rect 40786 17726 40798 17778
rect 40850 17726 40862 17778
rect 44258 17726 44270 17778
rect 44322 17726 44334 17778
rect 35534 17714 35586 17726
rect 39902 17714 39954 17726
rect 45054 17714 45106 17726
rect 6526 17666 6578 17678
rect 4610 17614 4622 17666
rect 4674 17614 4686 17666
rect 6526 17602 6578 17614
rect 8766 17666 8818 17678
rect 8766 17602 8818 17614
rect 9326 17666 9378 17678
rect 9886 17666 9938 17678
rect 9650 17614 9662 17666
rect 9714 17614 9726 17666
rect 9326 17602 9378 17614
rect 9886 17602 9938 17614
rect 10110 17666 10162 17678
rect 10110 17602 10162 17614
rect 11230 17666 11282 17678
rect 12014 17666 12066 17678
rect 11554 17614 11566 17666
rect 11618 17614 11630 17666
rect 11230 17602 11282 17614
rect 12014 17602 12066 17614
rect 15822 17666 15874 17678
rect 15822 17602 15874 17614
rect 16158 17666 16210 17678
rect 16158 17602 16210 17614
rect 17054 17666 17106 17678
rect 17054 17602 17106 17614
rect 17390 17666 17442 17678
rect 17390 17602 17442 17614
rect 17614 17666 17666 17678
rect 17614 17602 17666 17614
rect 18734 17666 18786 17678
rect 18734 17602 18786 17614
rect 20414 17666 20466 17678
rect 20414 17602 20466 17614
rect 21198 17666 21250 17678
rect 28254 17666 28306 17678
rect 30830 17666 30882 17678
rect 21522 17614 21534 17666
rect 21586 17614 21598 17666
rect 23202 17614 23214 17666
rect 23266 17614 23278 17666
rect 27010 17614 27022 17666
rect 27074 17614 27086 17666
rect 27458 17614 27470 17666
rect 27522 17614 27534 17666
rect 29474 17614 29486 17666
rect 29538 17614 29550 17666
rect 30594 17614 30606 17666
rect 30658 17614 30670 17666
rect 21198 17602 21250 17614
rect 28254 17602 28306 17614
rect 30830 17602 30882 17614
rect 31054 17666 31106 17678
rect 35422 17666 35474 17678
rect 33170 17614 33182 17666
rect 33234 17614 33246 17666
rect 33506 17614 33518 17666
rect 33570 17614 33582 17666
rect 38994 17614 39006 17666
rect 39058 17614 39070 17666
rect 40562 17614 40574 17666
rect 40626 17614 40638 17666
rect 41122 17614 41134 17666
rect 41186 17614 41198 17666
rect 41794 17614 41806 17666
rect 41858 17614 41870 17666
rect 46722 17614 46734 17666
rect 46786 17614 46798 17666
rect 31054 17602 31106 17614
rect 35422 17602 35474 17614
rect 2494 17554 2546 17566
rect 2494 17490 2546 17502
rect 3838 17554 3890 17566
rect 10334 17554 10386 17566
rect 4946 17502 4958 17554
rect 5010 17502 5022 17554
rect 6738 17502 6750 17554
rect 6802 17502 6814 17554
rect 7074 17502 7086 17554
rect 7138 17502 7150 17554
rect 3838 17490 3890 17502
rect 10334 17490 10386 17502
rect 12238 17554 12290 17566
rect 12238 17490 12290 17502
rect 13694 17554 13746 17566
rect 13694 17490 13746 17502
rect 13806 17554 13858 17566
rect 20078 17554 20130 17566
rect 13906 17502 13918 17554
rect 13970 17502 13982 17554
rect 13806 17490 13858 17502
rect 20078 17490 20130 17502
rect 21758 17554 21810 17566
rect 21758 17490 21810 17502
rect 21870 17554 21922 17566
rect 21870 17490 21922 17502
rect 22094 17554 22146 17566
rect 22094 17490 22146 17502
rect 24446 17554 24498 17566
rect 28478 17554 28530 17566
rect 26898 17502 26910 17554
rect 26962 17502 26974 17554
rect 27682 17502 27694 17554
rect 27746 17502 27758 17554
rect 24446 17490 24498 17502
rect 28478 17490 28530 17502
rect 28590 17554 28642 17566
rect 33070 17554 33122 17566
rect 29138 17502 29150 17554
rect 29202 17502 29214 17554
rect 28590 17490 28642 17502
rect 33070 17490 33122 17502
rect 35646 17554 35698 17566
rect 46610 17502 46622 17554
rect 46674 17502 46686 17554
rect 35646 17490 35698 17502
rect 2158 17442 2210 17454
rect 2158 17378 2210 17390
rect 9886 17442 9938 17454
rect 9886 17378 9938 17390
rect 13470 17442 13522 17454
rect 13470 17378 13522 17390
rect 16158 17442 16210 17454
rect 18286 17442 18338 17454
rect 16706 17390 16718 17442
rect 16770 17390 16782 17442
rect 16158 17378 16210 17390
rect 18286 17378 18338 17390
rect 20190 17442 20242 17454
rect 20190 17378 20242 17390
rect 22206 17442 22258 17454
rect 22206 17378 22258 17390
rect 22430 17442 22482 17454
rect 22430 17378 22482 17390
rect 22878 17442 22930 17454
rect 30942 17442 30994 17454
rect 27458 17390 27470 17442
rect 27522 17390 27534 17442
rect 22878 17378 22930 17390
rect 30942 17378 30994 17390
rect 31278 17442 31330 17454
rect 31278 17378 31330 17390
rect 31726 17442 31778 17454
rect 31726 17378 31778 17390
rect 34190 17442 34242 17454
rect 34190 17378 34242 17390
rect 35198 17442 35250 17454
rect 35198 17378 35250 17390
rect 36094 17442 36146 17454
rect 36094 17378 36146 17390
rect 1344 17274 48720 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48720 17274
rect 1344 17188 48720 17222
rect 9662 17106 9714 17118
rect 4722 17054 4734 17106
rect 4786 17054 4798 17106
rect 9662 17042 9714 17054
rect 10894 17106 10946 17118
rect 10894 17042 10946 17054
rect 11342 17106 11394 17118
rect 13022 17106 13074 17118
rect 12450 17054 12462 17106
rect 12514 17054 12526 17106
rect 11342 17042 11394 17054
rect 13022 17042 13074 17054
rect 13470 17106 13522 17118
rect 13470 17042 13522 17054
rect 14030 17106 14082 17118
rect 14030 17042 14082 17054
rect 14254 17106 14306 17118
rect 14254 17042 14306 17054
rect 15374 17106 15426 17118
rect 19070 17106 19122 17118
rect 18274 17054 18286 17106
rect 18338 17054 18350 17106
rect 15374 17042 15426 17054
rect 19070 17042 19122 17054
rect 19854 17106 19906 17118
rect 19854 17042 19906 17054
rect 27358 17106 27410 17118
rect 27358 17042 27410 17054
rect 28254 17106 28306 17118
rect 28254 17042 28306 17054
rect 29934 17106 29986 17118
rect 36990 17106 37042 17118
rect 35186 17054 35198 17106
rect 35250 17054 35262 17106
rect 36082 17054 36094 17106
rect 36146 17054 36158 17106
rect 29934 17042 29986 17054
rect 36990 17042 37042 17054
rect 37438 17106 37490 17118
rect 37438 17042 37490 17054
rect 37662 17106 37714 17118
rect 37662 17042 37714 17054
rect 37774 17106 37826 17118
rect 37774 17042 37826 17054
rect 38222 17106 38274 17118
rect 38222 17042 38274 17054
rect 40014 17106 40066 17118
rect 40014 17042 40066 17054
rect 40910 17106 40962 17118
rect 40910 17042 40962 17054
rect 41358 17106 41410 17118
rect 41358 17042 41410 17054
rect 41918 17106 41970 17118
rect 41918 17042 41970 17054
rect 42366 17106 42418 17118
rect 42366 17042 42418 17054
rect 42814 17106 42866 17118
rect 42814 17042 42866 17054
rect 47294 17106 47346 17118
rect 47294 17042 47346 17054
rect 11902 16994 11954 17006
rect 15486 16994 15538 17006
rect 8978 16942 8990 16994
rect 9042 16942 9054 16994
rect 14578 16942 14590 16994
rect 14642 16942 14654 16994
rect 11902 16930 11954 16942
rect 15486 16930 15538 16942
rect 16046 16994 16098 17006
rect 16046 16930 16098 16942
rect 16494 16994 16546 17006
rect 16494 16930 16546 16942
rect 16830 16994 16882 17006
rect 16830 16930 16882 16942
rect 17614 16994 17666 17006
rect 17614 16930 17666 16942
rect 20190 16994 20242 17006
rect 21310 16994 21362 17006
rect 20962 16942 20974 16994
rect 21026 16942 21038 16994
rect 20190 16930 20242 16942
rect 21310 16930 21362 16942
rect 21758 16994 21810 17006
rect 21758 16930 21810 16942
rect 25230 16994 25282 17006
rect 25230 16930 25282 16942
rect 27470 16994 27522 17006
rect 27470 16930 27522 16942
rect 27918 16994 27970 17006
rect 27918 16930 27970 16942
rect 28478 16994 28530 17006
rect 28478 16930 28530 16942
rect 30046 16994 30098 17006
rect 30046 16930 30098 16942
rect 30382 16994 30434 17006
rect 30382 16930 30434 16942
rect 31502 16994 31554 17006
rect 34190 16994 34242 17006
rect 33730 16942 33742 16994
rect 33794 16942 33806 16994
rect 31502 16930 31554 16942
rect 34190 16930 34242 16942
rect 34302 16994 34354 17006
rect 39454 16994 39506 17006
rect 38546 16942 38558 16994
rect 38610 16942 38622 16994
rect 34302 16930 34354 16942
rect 39454 16930 39506 16942
rect 41470 16994 41522 17006
rect 43810 16942 43822 16994
rect 43874 16942 43886 16994
rect 45714 16942 45726 16994
rect 45778 16942 45790 16994
rect 46050 16942 46062 16994
rect 46114 16942 46126 16994
rect 41470 16930 41522 16942
rect 17838 16882 17890 16894
rect 1698 16830 1710 16882
rect 1762 16830 1774 16882
rect 2258 16830 2270 16882
rect 2322 16830 2334 16882
rect 5842 16830 5854 16882
rect 5906 16830 5918 16882
rect 6626 16830 6638 16882
rect 6690 16830 6702 16882
rect 17838 16818 17890 16830
rect 18062 16882 18114 16894
rect 18062 16818 18114 16830
rect 18286 16882 18338 16894
rect 18286 16818 18338 16830
rect 19294 16882 19346 16894
rect 20750 16882 20802 16894
rect 20402 16830 20414 16882
rect 20466 16830 20478 16882
rect 19294 16818 19346 16830
rect 20750 16818 20802 16830
rect 22430 16882 22482 16894
rect 23774 16882 23826 16894
rect 23314 16830 23326 16882
rect 23378 16830 23390 16882
rect 22430 16818 22482 16830
rect 23774 16818 23826 16830
rect 24334 16882 24386 16894
rect 24334 16818 24386 16830
rect 27694 16882 27746 16894
rect 27694 16818 27746 16830
rect 28030 16882 28082 16894
rect 28030 16818 28082 16830
rect 28590 16882 28642 16894
rect 31166 16882 31218 16894
rect 30930 16830 30942 16882
rect 30994 16830 31006 16882
rect 28590 16818 28642 16830
rect 31166 16818 31218 16830
rect 31726 16882 31778 16894
rect 35534 16882 35586 16894
rect 33170 16830 33182 16882
rect 33234 16830 33246 16882
rect 31726 16818 31778 16830
rect 35534 16818 35586 16830
rect 36318 16882 36370 16894
rect 36318 16818 36370 16830
rect 36766 16882 36818 16894
rect 36766 16818 36818 16830
rect 37886 16882 37938 16894
rect 37886 16818 37938 16830
rect 38894 16882 38946 16894
rect 38894 16818 38946 16830
rect 41022 16882 41074 16894
rect 46734 16882 46786 16894
rect 43586 16830 43598 16882
rect 43650 16830 43662 16882
rect 41022 16818 41074 16830
rect 46734 16818 46786 16830
rect 5182 16770 5234 16782
rect 5182 16706 5234 16718
rect 10222 16770 10274 16782
rect 10222 16706 10274 16718
rect 18846 16770 18898 16782
rect 18846 16706 18898 16718
rect 19182 16770 19234 16782
rect 19182 16706 19234 16718
rect 20078 16770 20130 16782
rect 21982 16770 22034 16782
rect 21634 16718 21646 16770
rect 21698 16718 21710 16770
rect 20078 16706 20130 16718
rect 21982 16706 22034 16718
rect 22766 16770 22818 16782
rect 34638 16770 34690 16782
rect 25442 16718 25454 16770
rect 25506 16718 25518 16770
rect 33506 16718 33518 16770
rect 33570 16718 33582 16770
rect 22766 16706 22818 16718
rect 34638 16706 34690 16718
rect 34862 16770 34914 16782
rect 34862 16706 34914 16718
rect 35758 16770 35810 16782
rect 35758 16706 35810 16718
rect 36878 16770 36930 16782
rect 36878 16706 36930 16718
rect 39902 16770 39954 16782
rect 39902 16706 39954 16718
rect 44718 16770 44770 16782
rect 44718 16706 44770 16718
rect 47742 16770 47794 16782
rect 47742 16706 47794 16718
rect 12126 16658 12178 16670
rect 10210 16606 10222 16658
rect 10274 16655 10286 16658
rect 11554 16655 11566 16658
rect 10274 16609 11566 16655
rect 10274 16606 10286 16609
rect 11554 16606 11566 16609
rect 11618 16606 11630 16658
rect 12126 16594 12178 16606
rect 15374 16658 15426 16670
rect 15374 16594 15426 16606
rect 15822 16658 15874 16670
rect 15822 16594 15874 16606
rect 16158 16658 16210 16670
rect 16158 16594 16210 16606
rect 18622 16658 18674 16670
rect 18622 16594 18674 16606
rect 22990 16658 23042 16670
rect 22990 16594 23042 16606
rect 27358 16658 27410 16670
rect 27358 16594 27410 16606
rect 29934 16658 29986 16670
rect 29934 16594 29986 16606
rect 31950 16658 32002 16670
rect 31950 16594 32002 16606
rect 32174 16658 32226 16670
rect 32174 16594 32226 16606
rect 32622 16658 32674 16670
rect 32622 16594 32674 16606
rect 34190 16658 34242 16670
rect 34190 16594 34242 16606
rect 39790 16658 39842 16670
rect 39790 16594 39842 16606
rect 43150 16658 43202 16670
rect 43150 16594 43202 16606
rect 45166 16658 45218 16670
rect 45166 16594 45218 16606
rect 45502 16658 45554 16670
rect 45502 16594 45554 16606
rect 1344 16490 48720 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48720 16490
rect 1344 16404 48720 16438
rect 4174 16322 4226 16334
rect 4174 16258 4226 16270
rect 27134 16322 27186 16334
rect 27134 16258 27186 16270
rect 37326 16322 37378 16334
rect 37326 16258 37378 16270
rect 43262 16322 43314 16334
rect 43262 16258 43314 16270
rect 8318 16210 8370 16222
rect 8318 16146 8370 16158
rect 8878 16210 8930 16222
rect 11566 16210 11618 16222
rect 9986 16158 9998 16210
rect 10050 16158 10062 16210
rect 11106 16158 11118 16210
rect 11170 16158 11182 16210
rect 8878 16146 8930 16158
rect 11566 16146 11618 16158
rect 12798 16210 12850 16222
rect 30494 16210 30546 16222
rect 28354 16158 28366 16210
rect 28418 16158 28430 16210
rect 29362 16158 29374 16210
rect 29426 16158 29438 16210
rect 12798 16146 12850 16158
rect 30494 16146 30546 16158
rect 31278 16210 31330 16222
rect 31278 16146 31330 16158
rect 35982 16210 36034 16222
rect 35982 16146 36034 16158
rect 36990 16210 37042 16222
rect 36990 16146 37042 16158
rect 38110 16210 38162 16222
rect 41694 16210 41746 16222
rect 39106 16158 39118 16210
rect 39170 16158 39182 16210
rect 41234 16158 41246 16210
rect 41298 16158 41310 16210
rect 48290 16158 48302 16210
rect 48354 16158 48366 16210
rect 38110 16146 38162 16158
rect 41694 16146 41746 16158
rect 8542 16098 8594 16110
rect 15822 16098 15874 16110
rect 17614 16098 17666 16110
rect 4834 16046 4846 16098
rect 4898 16046 4910 16098
rect 14690 16046 14702 16098
rect 14754 16046 14766 16098
rect 16258 16046 16270 16098
rect 16322 16046 16334 16098
rect 8542 16034 8594 16046
rect 15822 16034 15874 16046
rect 17614 16034 17666 16046
rect 19406 16098 19458 16110
rect 27022 16098 27074 16110
rect 33406 16098 33458 16110
rect 35870 16098 35922 16110
rect 22418 16046 22430 16098
rect 22482 16046 22494 16098
rect 23986 16046 23998 16098
rect 24050 16046 24062 16098
rect 26450 16046 26462 16098
rect 26514 16046 26526 16098
rect 28242 16046 28254 16098
rect 28306 16046 28318 16098
rect 29474 16046 29486 16098
rect 29538 16046 29550 16098
rect 33730 16046 33742 16098
rect 33794 16046 33806 16098
rect 19406 16034 19458 16046
rect 27022 16034 27074 16046
rect 33406 16034 33458 16046
rect 35870 16034 35922 16046
rect 36542 16098 36594 16110
rect 38434 16046 38446 16098
rect 38498 16046 38510 16098
rect 43698 16046 43710 16098
rect 43762 16046 43774 16098
rect 45154 16046 45166 16098
rect 45218 16046 45230 16098
rect 45826 16046 45838 16098
rect 45890 16046 45902 16098
rect 36542 16034 36594 16046
rect 9550 15986 9602 15998
rect 10670 15986 10722 15998
rect 30158 15986 30210 15998
rect 34302 15986 34354 15998
rect 4946 15934 4958 15986
rect 5010 15934 5022 15986
rect 9650 15934 9662 15986
rect 9714 15934 9726 15986
rect 10770 15934 10782 15986
rect 10834 15934 10846 15986
rect 15362 15934 15374 15986
rect 15426 15934 15438 15986
rect 16818 15934 16830 15986
rect 16882 15934 16894 15986
rect 17938 15934 17950 15986
rect 18002 15934 18014 15986
rect 18498 15934 18510 15986
rect 18562 15934 18574 15986
rect 18946 15934 18958 15986
rect 19010 15934 19022 15986
rect 22306 15934 22318 15986
rect 22370 15934 22382 15986
rect 25666 15934 25678 15986
rect 25730 15934 25742 15986
rect 31826 15934 31838 15986
rect 31890 15934 31902 15986
rect 9550 15922 9602 15934
rect 10670 15922 10722 15934
rect 30158 15922 30210 15934
rect 34302 15922 34354 15934
rect 36094 15986 36146 15998
rect 36094 15922 36146 15934
rect 37550 15986 37602 15998
rect 43810 15934 43822 15986
rect 43874 15934 43886 15986
rect 37550 15922 37602 15934
rect 3838 15874 3890 15886
rect 3838 15810 3890 15822
rect 9214 15874 9266 15886
rect 9214 15810 9266 15822
rect 9438 15874 9490 15886
rect 9438 15810 9490 15822
rect 10334 15874 10386 15886
rect 10334 15810 10386 15822
rect 10558 15874 10610 15886
rect 20414 15874 20466 15886
rect 14914 15822 14926 15874
rect 14978 15822 14990 15874
rect 16258 15822 16270 15874
rect 16322 15822 16334 15874
rect 19282 15822 19294 15874
rect 19346 15822 19358 15874
rect 10558 15810 10610 15822
rect 20414 15810 20466 15822
rect 20862 15874 20914 15886
rect 20862 15810 20914 15822
rect 21646 15874 21698 15886
rect 24894 15874 24946 15886
rect 21970 15822 21982 15874
rect 22034 15822 22046 15874
rect 21646 15810 21698 15822
rect 24894 15810 24946 15822
rect 27134 15874 27186 15886
rect 27134 15810 27186 15822
rect 27806 15874 27858 15886
rect 27806 15810 27858 15822
rect 30606 15874 30658 15886
rect 42926 15874 42978 15886
rect 33170 15822 33182 15874
rect 33234 15822 33246 15874
rect 30606 15810 30658 15822
rect 42926 15810 42978 15822
rect 45054 15874 45106 15886
rect 45054 15810 45106 15822
rect 1344 15706 48720 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48720 15706
rect 1344 15620 48720 15654
rect 5070 15538 5122 15550
rect 20078 15538 20130 15550
rect 10210 15486 10222 15538
rect 10274 15486 10286 15538
rect 5070 15474 5122 15486
rect 20078 15474 20130 15486
rect 26910 15538 26962 15550
rect 26910 15474 26962 15486
rect 36206 15538 36258 15550
rect 36206 15474 36258 15486
rect 36318 15538 36370 15550
rect 36318 15474 36370 15486
rect 39006 15538 39058 15550
rect 45838 15538 45890 15550
rect 44818 15486 44830 15538
rect 44882 15486 44894 15538
rect 39006 15474 39058 15486
rect 45838 15474 45890 15486
rect 46622 15538 46674 15550
rect 46622 15474 46674 15486
rect 2158 15426 2210 15438
rect 2158 15362 2210 15374
rect 2494 15426 2546 15438
rect 2494 15362 2546 15374
rect 4286 15426 4338 15438
rect 4286 15362 4338 15374
rect 9662 15426 9714 15438
rect 9662 15362 9714 15374
rect 16494 15426 16546 15438
rect 16494 15362 16546 15374
rect 20414 15426 20466 15438
rect 20414 15362 20466 15374
rect 21422 15426 21474 15438
rect 21422 15362 21474 15374
rect 25902 15426 25954 15438
rect 38782 15426 38834 15438
rect 27010 15374 27022 15426
rect 27074 15374 27086 15426
rect 34962 15374 34974 15426
rect 35026 15374 35038 15426
rect 25902 15362 25954 15374
rect 38782 15362 38834 15374
rect 45502 15426 45554 15438
rect 45502 15362 45554 15374
rect 4622 15314 4674 15326
rect 14926 15314 14978 15326
rect 11666 15262 11678 15314
rect 11730 15262 11742 15314
rect 4622 15250 4674 15262
rect 14926 15250 14978 15262
rect 15374 15314 15426 15326
rect 15374 15250 15426 15262
rect 15598 15314 15650 15326
rect 15598 15250 15650 15262
rect 15822 15314 15874 15326
rect 25342 15314 25394 15326
rect 16034 15262 16046 15314
rect 16098 15262 16110 15314
rect 19618 15262 19630 15314
rect 19682 15262 19694 15314
rect 19842 15262 19854 15314
rect 19906 15262 19918 15314
rect 20626 15262 20638 15314
rect 20690 15262 20702 15314
rect 21970 15262 21982 15314
rect 22034 15262 22046 15314
rect 22194 15262 22206 15314
rect 22258 15262 22270 15314
rect 23538 15262 23550 15314
rect 23602 15262 23614 15314
rect 15822 15250 15874 15262
rect 25342 15250 25394 15262
rect 25566 15314 25618 15326
rect 34414 15314 34466 15326
rect 36094 15314 36146 15326
rect 36990 15314 37042 15326
rect 27794 15262 27806 15314
rect 27858 15262 27870 15314
rect 29922 15262 29934 15314
rect 29986 15262 29998 15314
rect 30482 15262 30494 15314
rect 30546 15262 30558 15314
rect 30930 15262 30942 15314
rect 30994 15262 31006 15314
rect 31490 15262 31502 15314
rect 31554 15262 31566 15314
rect 32274 15262 32286 15314
rect 32338 15262 32350 15314
rect 33170 15262 33182 15314
rect 33234 15262 33246 15314
rect 33394 15262 33406 15314
rect 33458 15262 33470 15314
rect 33730 15262 33742 15314
rect 33794 15262 33806 15314
rect 34626 15262 34638 15314
rect 34690 15262 34702 15314
rect 35746 15262 35758 15314
rect 35810 15262 35822 15314
rect 36642 15262 36654 15314
rect 36706 15262 36718 15314
rect 37538 15262 37550 15314
rect 37602 15262 37614 15314
rect 37874 15262 37886 15314
rect 37938 15262 37950 15314
rect 41682 15262 41694 15314
rect 41746 15262 41758 15314
rect 42466 15262 42478 15314
rect 42530 15262 42542 15314
rect 47282 15262 47294 15314
rect 47346 15262 47358 15314
rect 25566 15250 25618 15262
rect 34414 15250 34466 15262
rect 36094 15250 36146 15262
rect 36990 15250 37042 15262
rect 19742 15202 19794 15214
rect 24670 15202 24722 15214
rect 38110 15202 38162 15214
rect 12338 15150 12350 15202
rect 12402 15150 12414 15202
rect 14466 15150 14478 15202
rect 14530 15150 14542 15202
rect 21858 15150 21870 15202
rect 21922 15150 21934 15202
rect 23202 15150 23214 15202
rect 23266 15150 23278 15202
rect 35298 15150 35310 15202
rect 35362 15150 35374 15202
rect 19742 15138 19794 15150
rect 24670 15138 24722 15150
rect 38110 15138 38162 15150
rect 38334 15202 38386 15214
rect 38334 15138 38386 15150
rect 38446 15202 38498 15214
rect 38446 15138 38498 15150
rect 38894 15202 38946 15214
rect 38894 15138 38946 15150
rect 39566 15202 39618 15214
rect 46946 15150 46958 15202
rect 47010 15150 47022 15202
rect 39566 15138 39618 15150
rect 9886 15090 9938 15102
rect 9886 15026 9938 15038
rect 15262 15090 15314 15102
rect 15262 15026 15314 15038
rect 16382 15090 16434 15102
rect 26014 15090 26066 15102
rect 23426 15038 23438 15090
rect 23490 15038 23502 15090
rect 16382 15026 16434 15038
rect 26014 15026 26066 15038
rect 26126 15090 26178 15102
rect 26126 15026 26178 15038
rect 31726 15090 31778 15102
rect 31726 15026 31778 15038
rect 37214 15090 37266 15102
rect 37214 15026 37266 15038
rect 1344 14922 48720 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48720 14922
rect 1344 14836 48720 14870
rect 5742 14754 5794 14766
rect 5742 14690 5794 14702
rect 6078 14754 6130 14766
rect 6078 14690 6130 14702
rect 12574 14754 12626 14766
rect 20638 14754 20690 14766
rect 19730 14702 19742 14754
rect 19794 14702 19806 14754
rect 12574 14690 12626 14702
rect 20638 14690 20690 14702
rect 21198 14754 21250 14766
rect 47182 14754 47234 14766
rect 44930 14702 44942 14754
rect 44994 14751 45006 14754
rect 45378 14751 45390 14754
rect 44994 14705 45390 14751
rect 44994 14702 45006 14705
rect 45378 14702 45390 14705
rect 45442 14702 45454 14754
rect 21198 14690 21250 14702
rect 47182 14690 47234 14702
rect 11566 14642 11618 14654
rect 27470 14642 27522 14654
rect 10994 14590 11006 14642
rect 11058 14590 11070 14642
rect 25330 14590 25342 14642
rect 25394 14590 25406 14642
rect 26450 14590 26462 14642
rect 26514 14590 26526 14642
rect 11566 14578 11618 14590
rect 27470 14578 27522 14590
rect 35646 14642 35698 14654
rect 35646 14578 35698 14590
rect 36206 14642 36258 14654
rect 36206 14578 36258 14590
rect 37886 14642 37938 14654
rect 44942 14642 44994 14654
rect 39106 14590 39118 14642
rect 39170 14590 39182 14642
rect 41234 14590 41246 14642
rect 41298 14590 41310 14642
rect 37886 14578 37938 14590
rect 44942 14578 44994 14590
rect 45390 14642 45442 14654
rect 45390 14578 45442 14590
rect 17166 14530 17218 14542
rect 1698 14478 1710 14530
rect 1762 14478 1774 14530
rect 2258 14478 2270 14530
rect 2322 14478 2334 14530
rect 7410 14478 7422 14530
rect 7474 14478 7486 14530
rect 7858 14478 7870 14530
rect 7922 14478 7934 14530
rect 8530 14478 8542 14530
rect 8594 14478 8606 14530
rect 17166 14466 17218 14478
rect 17278 14530 17330 14542
rect 17278 14466 17330 14478
rect 17726 14530 17778 14542
rect 17726 14466 17778 14478
rect 19406 14530 19458 14542
rect 19406 14466 19458 14478
rect 20078 14530 20130 14542
rect 20078 14466 20130 14478
rect 20302 14530 20354 14542
rect 22430 14530 22482 14542
rect 26014 14530 26066 14542
rect 27582 14530 27634 14542
rect 42814 14530 42866 14542
rect 21522 14478 21534 14530
rect 21586 14478 21598 14530
rect 22978 14478 22990 14530
rect 23042 14478 23054 14530
rect 23538 14478 23550 14530
rect 23602 14478 23614 14530
rect 24322 14478 24334 14530
rect 24386 14478 24398 14530
rect 25218 14478 25230 14530
rect 25282 14478 25294 14530
rect 26226 14478 26238 14530
rect 26290 14478 26302 14530
rect 27906 14478 27918 14530
rect 27970 14478 27982 14530
rect 29810 14478 29822 14530
rect 29874 14478 29886 14530
rect 30370 14478 30382 14530
rect 30434 14478 30446 14530
rect 31378 14478 31390 14530
rect 31442 14478 31454 14530
rect 33394 14478 33406 14530
rect 33458 14478 33470 14530
rect 37426 14478 37438 14530
rect 37490 14478 37502 14530
rect 38434 14478 38446 14530
rect 38498 14478 38510 14530
rect 20302 14466 20354 14478
rect 22430 14466 22482 14478
rect 26014 14466 26066 14478
rect 27582 14466 27634 14478
rect 42814 14466 42866 14478
rect 7646 14418 7698 14430
rect 6290 14366 6302 14418
rect 6354 14366 6366 14418
rect 6850 14366 6862 14418
rect 6914 14366 6926 14418
rect 7646 14354 7698 14366
rect 12910 14418 12962 14430
rect 12910 14354 12962 14366
rect 17054 14418 17106 14430
rect 17054 14354 17106 14366
rect 18734 14418 18786 14430
rect 18734 14354 18786 14366
rect 20750 14418 20802 14430
rect 20750 14354 20802 14366
rect 21310 14418 21362 14430
rect 21310 14354 21362 14366
rect 21758 14418 21810 14430
rect 23998 14418 24050 14430
rect 22754 14366 22766 14418
rect 22818 14366 22830 14418
rect 21758 14354 21810 14366
rect 23998 14354 24050 14366
rect 24110 14418 24162 14430
rect 24110 14354 24162 14366
rect 28366 14418 28418 14430
rect 33966 14418 34018 14430
rect 31042 14366 31054 14418
rect 31106 14366 31118 14418
rect 31490 14366 31502 14418
rect 31554 14366 31566 14418
rect 28366 14354 28418 14366
rect 33966 14354 34018 14366
rect 35534 14418 35586 14430
rect 35534 14354 35586 14366
rect 36990 14418 37042 14430
rect 36990 14354 37042 14366
rect 42478 14418 42530 14430
rect 47394 14366 47406 14418
rect 47458 14366 47470 14418
rect 47730 14366 47742 14418
rect 47794 14366 47806 14418
rect 42478 14354 42530 14366
rect 12686 14306 12738 14318
rect 4722 14254 4734 14306
rect 4786 14254 4798 14306
rect 12686 14242 12738 14254
rect 14366 14306 14418 14318
rect 18622 14306 18674 14318
rect 16594 14254 16606 14306
rect 16658 14254 16670 14306
rect 18050 14254 18062 14306
rect 18114 14254 18126 14306
rect 14366 14242 14418 14254
rect 18622 14242 18674 14254
rect 18958 14306 19010 14318
rect 18958 14242 19010 14254
rect 19182 14306 19234 14318
rect 27358 14306 27410 14318
rect 22082 14254 22094 14306
rect 22146 14254 22158 14306
rect 19182 14242 19234 14254
rect 27358 14242 27410 14254
rect 28478 14306 28530 14318
rect 28478 14242 28530 14254
rect 28702 14306 28754 14318
rect 36878 14306 36930 14318
rect 32386 14254 32398 14306
rect 32450 14254 32462 14306
rect 28702 14242 28754 14254
rect 36878 14242 36930 14254
rect 37214 14306 37266 14318
rect 37214 14242 37266 14254
rect 41694 14306 41746 14318
rect 41694 14242 41746 14254
rect 46846 14306 46898 14318
rect 46846 14242 46898 14254
rect 1344 14138 48720 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48720 14138
rect 1344 14052 48720 14086
rect 6974 13970 7026 13982
rect 6514 13918 6526 13970
rect 6578 13918 6590 13970
rect 6974 13906 7026 13918
rect 7422 13970 7474 13982
rect 7422 13906 7474 13918
rect 15710 13970 15762 13982
rect 15710 13906 15762 13918
rect 21310 13970 21362 13982
rect 21310 13906 21362 13918
rect 25230 13970 25282 13982
rect 34526 13970 34578 13982
rect 28242 13918 28254 13970
rect 28306 13918 28318 13970
rect 25230 13906 25282 13918
rect 34526 13906 34578 13918
rect 36094 13970 36146 13982
rect 37886 13970 37938 13982
rect 36978 13918 36990 13970
rect 37042 13918 37054 13970
rect 36094 13906 36146 13918
rect 37886 13906 37938 13918
rect 41134 13970 41186 13982
rect 41134 13906 41186 13918
rect 45166 13970 45218 13982
rect 45166 13906 45218 13918
rect 45502 13970 45554 13982
rect 45502 13906 45554 13918
rect 48302 13970 48354 13982
rect 48302 13906 48354 13918
rect 15262 13858 15314 13870
rect 17390 13858 17442 13870
rect 7970 13806 7982 13858
rect 8034 13806 8046 13858
rect 8418 13806 8430 13858
rect 8482 13806 8494 13858
rect 12002 13806 12014 13858
rect 12066 13806 12078 13858
rect 15922 13806 15934 13858
rect 15986 13806 15998 13858
rect 15262 13794 15314 13806
rect 17390 13794 17442 13806
rect 17838 13858 17890 13870
rect 21198 13858 21250 13870
rect 19058 13806 19070 13858
rect 19122 13806 19134 13858
rect 20514 13806 20526 13858
rect 20578 13806 20590 13858
rect 17838 13794 17890 13806
rect 21198 13794 21250 13806
rect 25566 13858 25618 13870
rect 25566 13794 25618 13806
rect 26686 13858 26738 13870
rect 31838 13858 31890 13870
rect 29250 13806 29262 13858
rect 29314 13806 29326 13858
rect 26686 13794 26738 13806
rect 31838 13794 31890 13806
rect 34078 13858 34130 13870
rect 35198 13858 35250 13870
rect 34850 13806 34862 13858
rect 34914 13806 34926 13858
rect 46386 13806 46398 13858
rect 46450 13806 46462 13858
rect 34078 13794 34130 13806
rect 35198 13794 35250 13806
rect 7758 13746 7810 13758
rect 19518 13746 19570 13758
rect 21422 13746 21474 13758
rect 28590 13746 28642 13758
rect 30830 13746 30882 13758
rect 35758 13746 35810 13758
rect 3602 13694 3614 13746
rect 3666 13694 3678 13746
rect 4162 13694 4174 13746
rect 4226 13694 4238 13746
rect 11330 13694 11342 13746
rect 11394 13694 11406 13746
rect 16146 13694 16158 13746
rect 16210 13694 16222 13746
rect 17602 13694 17614 13746
rect 17666 13694 17678 13746
rect 20066 13694 20078 13746
rect 20130 13694 20142 13746
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 26450 13694 26462 13746
rect 26514 13694 26526 13746
rect 27234 13694 27246 13746
rect 27298 13694 27310 13746
rect 27682 13694 27694 13746
rect 27746 13694 27758 13746
rect 29138 13694 29150 13746
rect 29202 13694 29214 13746
rect 31042 13694 31054 13746
rect 31106 13694 31118 13746
rect 33618 13694 33630 13746
rect 33682 13694 33694 13746
rect 7758 13682 7810 13694
rect 19518 13682 19570 13694
rect 21422 13682 21474 13694
rect 28590 13682 28642 13694
rect 30830 13682 30882 13694
rect 35758 13682 35810 13694
rect 37326 13746 37378 13758
rect 37326 13682 37378 13694
rect 38222 13746 38274 13758
rect 38222 13682 38274 13694
rect 45838 13746 45890 13758
rect 46498 13694 46510 13746
rect 46562 13694 46574 13746
rect 45838 13682 45890 13694
rect 15038 13634 15090 13646
rect 14130 13582 14142 13634
rect 14194 13582 14206 13634
rect 15038 13570 15090 13582
rect 15486 13634 15538 13646
rect 15486 13570 15538 13582
rect 17502 13634 17554 13646
rect 26126 13634 26178 13646
rect 38670 13634 38722 13646
rect 19618 13582 19630 13634
rect 19682 13582 19694 13634
rect 22530 13582 22542 13634
rect 22594 13582 22606 13634
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 33170 13582 33182 13634
rect 33234 13582 33246 13634
rect 36530 13582 36542 13634
rect 36594 13582 36606 13634
rect 17502 13570 17554 13582
rect 26126 13570 26178 13582
rect 38670 13570 38722 13582
rect 15710 13522 15762 13534
rect 27570 13470 27582 13522
rect 27634 13470 27646 13522
rect 15710 13458 15762 13470
rect 1344 13354 48720 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48720 13354
rect 1344 13268 48720 13302
rect 7982 13186 8034 13198
rect 28254 13186 28306 13198
rect 15362 13134 15374 13186
rect 15426 13134 15438 13186
rect 7982 13122 8034 13134
rect 28254 13122 28306 13134
rect 28590 13186 28642 13198
rect 28590 13122 28642 13134
rect 6750 13074 6802 13086
rect 13470 13074 13522 13086
rect 14814 13074 14866 13086
rect 6178 13022 6190 13074
rect 6242 13022 6254 13074
rect 12786 13022 12798 13074
rect 12850 13022 12862 13074
rect 14354 13022 14366 13074
rect 14418 13022 14430 13074
rect 6750 13010 6802 13022
rect 13470 13010 13522 13022
rect 14814 13010 14866 13022
rect 16382 13074 16434 13086
rect 16382 13010 16434 13022
rect 21646 13074 21698 13086
rect 21646 13010 21698 13022
rect 24558 13074 24610 13086
rect 30270 13074 30322 13086
rect 32734 13074 32786 13086
rect 29586 13022 29598 13074
rect 29650 13022 29662 13074
rect 31154 13022 31166 13074
rect 31218 13022 31230 13074
rect 32274 13022 32286 13074
rect 32338 13022 32350 13074
rect 24558 13010 24610 13022
rect 30270 13010 30322 13022
rect 32734 13010 32786 13022
rect 33182 13074 33234 13086
rect 33182 13010 33234 13022
rect 33742 13074 33794 13086
rect 33742 13010 33794 13022
rect 34078 13074 34130 13086
rect 35198 13074 35250 13086
rect 34962 13022 34974 13074
rect 35026 13022 35038 13074
rect 34078 13010 34130 13022
rect 35198 13010 35250 13022
rect 36318 13074 36370 13086
rect 37986 13022 37998 13074
rect 38050 13022 38062 13074
rect 44258 13022 44270 13074
rect 44322 13022 44334 13074
rect 48290 13022 48302 13074
rect 48354 13022 48366 13074
rect 36318 13010 36370 13022
rect 4174 12962 4226 12974
rect 5742 12962 5794 12974
rect 15038 12962 15090 12974
rect 17390 12962 17442 12974
rect 4946 12910 4958 12962
rect 5010 12910 5022 12962
rect 8418 12910 8430 12962
rect 8482 12910 8494 12962
rect 14130 12910 14142 12962
rect 14194 12910 14206 12962
rect 15698 12910 15710 12962
rect 15762 12910 15774 12962
rect 16930 12910 16942 12962
rect 16994 12910 17006 12962
rect 4174 12898 4226 12910
rect 5742 12898 5794 12910
rect 15038 12898 15090 12910
rect 17390 12898 17442 12910
rect 17838 12962 17890 12974
rect 25678 12962 25730 12974
rect 27918 12962 27970 12974
rect 33854 12962 33906 12974
rect 24994 12910 25006 12962
rect 25058 12910 25070 12962
rect 26450 12910 26462 12962
rect 26514 12910 26526 12962
rect 27346 12910 27358 12962
rect 27410 12910 27422 12962
rect 29250 12910 29262 12962
rect 29314 12910 29326 12962
rect 30706 12910 30718 12962
rect 30770 12910 30782 12962
rect 31938 12910 31950 12962
rect 32002 12910 32014 12962
rect 17838 12898 17890 12910
rect 25678 12898 25730 12910
rect 27918 12898 27970 12910
rect 33854 12898 33906 12910
rect 35534 12962 35586 12974
rect 40786 12910 40798 12962
rect 40850 12910 40862 12962
rect 41122 12910 41134 12962
rect 41186 12910 41198 12962
rect 41906 12910 41918 12962
rect 41970 12910 41982 12962
rect 45154 12910 45166 12962
rect 45218 12910 45230 12962
rect 45938 12910 45950 12962
rect 46002 12910 46014 12962
rect 35534 12898 35586 12910
rect 2606 12850 2658 12862
rect 2606 12786 2658 12798
rect 3838 12850 3890 12862
rect 15934 12850 15986 12862
rect 4834 12798 4846 12850
rect 4898 12798 4910 12850
rect 8754 12798 8766 12850
rect 8818 12798 8830 12850
rect 3838 12786 3890 12798
rect 15934 12786 15986 12798
rect 16494 12850 16546 12862
rect 16494 12786 16546 12798
rect 17726 12850 17778 12862
rect 17726 12786 17778 12798
rect 25454 12850 25506 12862
rect 25454 12786 25506 12798
rect 26126 12850 26178 12862
rect 34190 12850 34242 12862
rect 27682 12798 27694 12850
rect 27746 12798 27758 12850
rect 31714 12798 31726 12850
rect 31778 12798 31790 12850
rect 26126 12786 26178 12798
rect 34190 12786 34242 12798
rect 34414 12850 34466 12862
rect 37326 12850 37378 12862
rect 35858 12798 35870 12850
rect 35922 12798 35934 12850
rect 40114 12798 40126 12850
rect 40178 12798 40190 12850
rect 34414 12786 34466 12798
rect 37326 12786 37378 12798
rect 2270 12738 2322 12750
rect 2270 12674 2322 12686
rect 7646 12738 7698 12750
rect 7646 12674 7698 12686
rect 12126 12738 12178 12750
rect 12126 12674 12178 12686
rect 12350 12738 12402 12750
rect 12350 12674 12402 12686
rect 16158 12738 16210 12750
rect 16158 12674 16210 12686
rect 16270 12738 16322 12750
rect 16270 12674 16322 12686
rect 16718 12738 16770 12750
rect 16718 12674 16770 12686
rect 17614 12738 17666 12750
rect 17614 12674 17666 12686
rect 22094 12738 22146 12750
rect 22094 12674 22146 12686
rect 23886 12738 23938 12750
rect 23886 12674 23938 12686
rect 24222 12738 24274 12750
rect 24222 12674 24274 12686
rect 25902 12738 25954 12750
rect 25902 12674 25954 12686
rect 26238 12738 26290 12750
rect 26238 12674 26290 12686
rect 27806 12738 27858 12750
rect 27806 12674 27858 12686
rect 28366 12738 28418 12750
rect 28366 12674 28418 12686
rect 32622 12738 32674 12750
rect 32622 12674 32674 12686
rect 37662 12738 37714 12750
rect 37662 12674 37714 12686
rect 44942 12738 44994 12750
rect 44942 12674 44994 12686
rect 1344 12570 48720 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48720 12570
rect 1344 12484 48720 12518
rect 5294 12402 5346 12414
rect 4722 12350 4734 12402
rect 4786 12350 4798 12402
rect 5294 12338 5346 12350
rect 5742 12402 5794 12414
rect 5742 12338 5794 12350
rect 13134 12402 13186 12414
rect 13134 12338 13186 12350
rect 15934 12402 15986 12414
rect 15934 12338 15986 12350
rect 17726 12402 17778 12414
rect 17726 12338 17778 12350
rect 18510 12402 18562 12414
rect 25454 12402 25506 12414
rect 22530 12350 22542 12402
rect 22594 12350 22606 12402
rect 18510 12338 18562 12350
rect 25454 12338 25506 12350
rect 26238 12402 26290 12414
rect 26238 12338 26290 12350
rect 30494 12402 30546 12414
rect 38670 12402 38722 12414
rect 35410 12350 35422 12402
rect 35474 12350 35486 12402
rect 30494 12338 30546 12350
rect 38670 12338 38722 12350
rect 39230 12402 39282 12414
rect 39230 12338 39282 12350
rect 42254 12402 42306 12414
rect 42254 12338 42306 12350
rect 46286 12402 46338 12414
rect 46286 12338 46338 12350
rect 7870 12290 7922 12302
rect 7870 12226 7922 12238
rect 8206 12290 8258 12302
rect 8206 12226 8258 12238
rect 14590 12290 14642 12302
rect 17614 12290 17666 12302
rect 16258 12238 16270 12290
rect 16322 12238 16334 12290
rect 14590 12226 14642 12238
rect 17614 12226 17666 12238
rect 18622 12290 18674 12302
rect 18622 12226 18674 12238
rect 21086 12290 21138 12302
rect 21086 12226 21138 12238
rect 21422 12290 21474 12302
rect 21422 12226 21474 12238
rect 21982 12290 22034 12302
rect 21982 12226 22034 12238
rect 22318 12290 22370 12302
rect 28142 12290 28194 12302
rect 46622 12290 46674 12302
rect 27570 12238 27582 12290
rect 27634 12238 27646 12290
rect 31490 12238 31502 12290
rect 31554 12238 31566 12290
rect 32274 12238 32286 12290
rect 32338 12238 32350 12290
rect 44146 12238 44158 12290
rect 44210 12238 44222 12290
rect 22318 12226 22370 12238
rect 28142 12226 28194 12238
rect 46622 12226 46674 12238
rect 14366 12178 14418 12190
rect 1698 12126 1710 12178
rect 1762 12126 1774 12178
rect 2258 12126 2270 12178
rect 2322 12126 2334 12178
rect 14366 12114 14418 12126
rect 15038 12178 15090 12190
rect 21758 12178 21810 12190
rect 17938 12126 17950 12178
rect 18002 12126 18014 12178
rect 20850 12126 20862 12178
rect 20914 12126 20926 12178
rect 15038 12114 15090 12126
rect 21758 12114 21810 12126
rect 22654 12178 22706 12190
rect 25902 12178 25954 12190
rect 30270 12178 30322 12190
rect 32510 12178 32562 12190
rect 23090 12126 23102 12178
rect 23154 12126 23166 12178
rect 26562 12126 26574 12178
rect 26626 12126 26638 12178
rect 27682 12126 27694 12178
rect 27746 12126 27758 12178
rect 29138 12126 29150 12178
rect 29202 12126 29214 12178
rect 29922 12126 29934 12178
rect 29986 12126 29998 12178
rect 30706 12126 30718 12178
rect 30770 12126 30782 12178
rect 31042 12126 31054 12178
rect 31106 12126 31118 12178
rect 22654 12114 22706 12126
rect 25902 12114 25954 12126
rect 30270 12114 30322 12126
rect 32510 12114 32562 12126
rect 33070 12178 33122 12190
rect 34302 12178 34354 12190
rect 33506 12126 33518 12178
rect 33570 12126 33582 12178
rect 33070 12114 33122 12126
rect 34302 12114 34354 12126
rect 34526 12178 34578 12190
rect 35758 12178 35810 12190
rect 37998 12178 38050 12190
rect 34850 12126 34862 12178
rect 34914 12126 34926 12178
rect 36082 12126 36094 12178
rect 36146 12126 36158 12178
rect 37426 12126 37438 12178
rect 37490 12126 37502 12178
rect 34526 12114 34578 12126
rect 35758 12114 35810 12126
rect 37998 12114 38050 12126
rect 42590 12178 42642 12190
rect 42590 12114 42642 12126
rect 43262 12178 43314 12190
rect 44370 12126 44382 12178
rect 44434 12126 44446 12178
rect 43262 12114 43314 12126
rect 14478 12066 14530 12078
rect 14478 12002 14530 12014
rect 15598 12066 15650 12078
rect 15598 12002 15650 12014
rect 21870 12066 21922 12078
rect 21870 12002 21922 12014
rect 23550 12066 23602 12078
rect 32622 12066 32674 12078
rect 27010 12014 27022 12066
rect 27074 12014 27086 12066
rect 30482 12014 30494 12066
rect 30546 12014 30558 12066
rect 23550 12002 23602 12014
rect 32622 12002 32674 12014
rect 38110 12066 38162 12078
rect 38110 12002 38162 12014
rect 38446 12066 38498 12078
rect 41022 12066 41074 12078
rect 38770 12014 38782 12066
rect 38834 12014 38846 12066
rect 38446 12002 38498 12014
rect 41022 12002 41074 12014
rect 43598 12066 43650 12078
rect 43598 12002 43650 12014
rect 18398 11954 18450 11966
rect 29822 11954 29874 11966
rect 22866 11902 22878 11954
rect 22930 11902 22942 11954
rect 28578 11902 28590 11954
rect 28642 11902 28654 11954
rect 18398 11890 18450 11902
rect 29822 11890 29874 11902
rect 36094 11954 36146 11966
rect 36094 11890 36146 11902
rect 36430 11954 36482 11966
rect 36430 11890 36482 11902
rect 1344 11786 48720 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48720 11786
rect 1344 11700 48720 11734
rect 14926 11618 14978 11630
rect 14926 11554 14978 11566
rect 15374 11618 15426 11630
rect 15374 11554 15426 11566
rect 19182 11618 19234 11630
rect 19182 11554 19234 11566
rect 22878 11618 22930 11630
rect 22878 11554 22930 11566
rect 47406 11618 47458 11630
rect 47406 11554 47458 11566
rect 11454 11506 11506 11518
rect 10994 11454 11006 11506
rect 11058 11454 11070 11506
rect 11454 11442 11506 11454
rect 13918 11506 13970 11518
rect 13918 11442 13970 11454
rect 14702 11506 14754 11518
rect 14702 11442 14754 11454
rect 16046 11506 16098 11518
rect 18398 11506 18450 11518
rect 17602 11454 17614 11506
rect 17666 11454 17678 11506
rect 16046 11442 16098 11454
rect 18398 11442 18450 11454
rect 18958 11506 19010 11518
rect 27022 11506 27074 11518
rect 26450 11454 26462 11506
rect 26514 11454 26526 11506
rect 27794 11454 27806 11506
rect 27858 11454 27870 11506
rect 29922 11454 29934 11506
rect 29986 11454 29998 11506
rect 32162 11454 32174 11506
rect 32226 11454 32238 11506
rect 35410 11454 35422 11506
rect 35474 11454 35486 11506
rect 38994 11454 39006 11506
rect 39058 11454 39070 11506
rect 18958 11442 19010 11454
rect 27022 11442 27074 11454
rect 12910 11394 12962 11406
rect 7858 11342 7870 11394
rect 7922 11342 7934 11394
rect 8530 11342 8542 11394
rect 8594 11342 8606 11394
rect 12910 11330 12962 11342
rect 14254 11394 14306 11406
rect 14254 11330 14306 11342
rect 14478 11394 14530 11406
rect 14478 11330 14530 11342
rect 15934 11394 15986 11406
rect 20862 11394 20914 11406
rect 17826 11342 17838 11394
rect 17890 11342 17902 11394
rect 20290 11342 20302 11394
rect 20354 11342 20366 11394
rect 20514 11342 20526 11394
rect 20578 11342 20590 11394
rect 15934 11330 15986 11342
rect 20862 11330 20914 11342
rect 21422 11394 21474 11406
rect 21422 11330 21474 11342
rect 21534 11394 21586 11406
rect 23102 11394 23154 11406
rect 36990 11394 37042 11406
rect 38110 11394 38162 11406
rect 22082 11342 22094 11394
rect 22146 11342 22158 11394
rect 22642 11342 22654 11394
rect 22706 11342 22718 11394
rect 23650 11342 23662 11394
rect 23714 11342 23726 11394
rect 28466 11342 28478 11394
rect 28530 11342 28542 11394
rect 29586 11342 29598 11394
rect 29650 11342 29662 11394
rect 30594 11342 30606 11394
rect 30658 11342 30670 11394
rect 31602 11342 31614 11394
rect 31666 11342 31678 11394
rect 32610 11342 32622 11394
rect 32674 11342 32686 11394
rect 35074 11342 35086 11394
rect 35138 11342 35150 11394
rect 35522 11342 35534 11394
rect 35586 11342 35598 11394
rect 37202 11342 37214 11394
rect 37266 11342 37278 11394
rect 41906 11342 41918 11394
rect 41970 11342 41982 11394
rect 46946 11342 46958 11394
rect 47010 11342 47022 11394
rect 21534 11330 21586 11342
rect 23102 11330 23154 11342
rect 36990 11330 37042 11342
rect 38110 11330 38162 11342
rect 12350 11282 12402 11294
rect 12350 11218 12402 11230
rect 21646 11282 21698 11294
rect 21646 11218 21698 11230
rect 23214 11282 23266 11294
rect 29374 11282 29426 11294
rect 37774 11282 37826 11294
rect 24322 11230 24334 11282
rect 24386 11230 24398 11282
rect 30370 11230 30382 11282
rect 30434 11230 30446 11282
rect 31826 11230 31838 11282
rect 31890 11230 31902 11282
rect 32498 11230 32510 11282
rect 32562 11230 32574 11282
rect 34514 11230 34526 11282
rect 34578 11230 34590 11282
rect 36194 11230 36206 11282
rect 36258 11230 36270 11282
rect 23214 11218 23266 11230
rect 29374 11218 29426 11230
rect 37774 11218 37826 11230
rect 38222 11282 38274 11294
rect 41122 11230 41134 11282
rect 41186 11230 41198 11282
rect 46610 11230 46622 11282
rect 46674 11230 46686 11282
rect 38222 11218 38274 11230
rect 4958 11170 5010 11182
rect 4958 11106 5010 11118
rect 15710 11170 15762 11182
rect 15710 11106 15762 11118
rect 16158 11170 16210 11182
rect 20750 11170 20802 11182
rect 19506 11118 19518 11170
rect 19570 11118 19582 11170
rect 16158 11106 16210 11118
rect 20750 11106 20802 11118
rect 38446 11170 38498 11182
rect 38446 11106 38498 11118
rect 42366 11170 42418 11182
rect 42366 11106 42418 11118
rect 45502 11170 45554 11182
rect 45502 11106 45554 11118
rect 47742 11170 47794 11182
rect 47742 11106 47794 11118
rect 1344 11002 48720 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48720 11002
rect 1344 10916 48720 10950
rect 15150 10834 15202 10846
rect 4722 10782 4734 10834
rect 4786 10782 4798 10834
rect 8194 10782 8206 10834
rect 8258 10782 8270 10834
rect 15150 10770 15202 10782
rect 15262 10834 15314 10846
rect 15262 10770 15314 10782
rect 15374 10834 15426 10846
rect 15374 10770 15426 10782
rect 18062 10834 18114 10846
rect 18062 10770 18114 10782
rect 18958 10834 19010 10846
rect 18958 10770 19010 10782
rect 19070 10834 19122 10846
rect 19070 10770 19122 10782
rect 21198 10834 21250 10846
rect 21198 10770 21250 10782
rect 22318 10834 22370 10846
rect 22318 10770 22370 10782
rect 22542 10834 22594 10846
rect 22542 10770 22594 10782
rect 22990 10834 23042 10846
rect 38110 10834 38162 10846
rect 27010 10782 27022 10834
rect 27074 10782 27086 10834
rect 33282 10782 33294 10834
rect 33346 10782 33358 10834
rect 22990 10770 23042 10782
rect 38110 10770 38162 10782
rect 39454 10834 39506 10846
rect 45266 10782 45278 10834
rect 45330 10782 45342 10834
rect 39454 10770 39506 10782
rect 19966 10722 20018 10734
rect 14018 10670 14030 10722
rect 14082 10670 14094 10722
rect 19966 10658 20018 10670
rect 20078 10722 20130 10734
rect 20078 10658 20130 10670
rect 20414 10722 20466 10734
rect 35646 10722 35698 10734
rect 31826 10670 31838 10722
rect 31890 10670 31902 10722
rect 33170 10670 33182 10722
rect 33234 10670 33246 10722
rect 20414 10658 20466 10670
rect 35646 10658 35698 10670
rect 37326 10722 37378 10734
rect 38558 10722 38610 10734
rect 37538 10670 37550 10722
rect 37602 10670 37614 10722
rect 37326 10658 37378 10670
rect 38558 10658 38610 10670
rect 38670 10722 38722 10734
rect 38670 10658 38722 10670
rect 38782 10722 38834 10734
rect 38782 10658 38834 10670
rect 39678 10722 39730 10734
rect 47294 10722 47346 10734
rect 45714 10670 45726 10722
rect 45778 10670 45790 10722
rect 46274 10670 46286 10722
rect 46338 10670 46350 10722
rect 39678 10658 39730 10670
rect 47294 10658 47346 10670
rect 47630 10722 47682 10734
rect 47630 10658 47682 10670
rect 8654 10610 8706 10622
rect 19630 10610 19682 10622
rect 1698 10558 1710 10610
rect 1762 10558 1774 10610
rect 2258 10558 2270 10610
rect 2322 10558 2334 10610
rect 5170 10558 5182 10610
rect 5234 10558 5246 10610
rect 5842 10558 5854 10610
rect 5906 10558 5918 10610
rect 9650 10558 9662 10610
rect 9714 10558 9726 10610
rect 13906 10558 13918 10610
rect 13970 10558 13982 10610
rect 14802 10558 14814 10610
rect 14866 10558 14878 10610
rect 17826 10558 17838 10610
rect 17890 10558 17902 10610
rect 19282 10558 19294 10610
rect 19346 10558 19358 10610
rect 8654 10546 8706 10558
rect 19630 10546 19682 10558
rect 19742 10610 19794 10622
rect 21086 10610 21138 10622
rect 20738 10558 20750 10610
rect 20802 10558 20814 10610
rect 19742 10546 19794 10558
rect 21086 10546 21138 10558
rect 21422 10610 21474 10622
rect 21422 10546 21474 10558
rect 21870 10610 21922 10622
rect 27358 10610 27410 10622
rect 23202 10558 23214 10610
rect 23266 10558 23278 10610
rect 21870 10546 21922 10558
rect 27358 10546 27410 10558
rect 27694 10610 27746 10622
rect 29486 10610 29538 10622
rect 35198 10610 35250 10622
rect 28018 10558 28030 10610
rect 28082 10558 28094 10610
rect 30706 10558 30718 10610
rect 30770 10558 30782 10610
rect 31042 10558 31054 10610
rect 31106 10558 31118 10610
rect 34626 10558 34638 10610
rect 34690 10558 34702 10610
rect 27694 10546 27746 10558
rect 29486 10546 29538 10558
rect 35198 10546 35250 10558
rect 37774 10610 37826 10622
rect 39790 10610 39842 10622
rect 46510 10610 46562 10622
rect 37874 10558 37886 10610
rect 37938 10558 37950 10610
rect 42130 10558 42142 10610
rect 42194 10558 42206 10610
rect 42914 10558 42926 10610
rect 42978 10558 42990 10610
rect 37774 10546 37826 10558
rect 39790 10546 39842 10558
rect 46510 10546 46562 10558
rect 15822 10498 15874 10510
rect 10322 10446 10334 10498
rect 10386 10446 10398 10498
rect 12450 10446 12462 10498
rect 12514 10446 12526 10498
rect 14354 10446 14366 10498
rect 14418 10495 14430 10498
rect 14690 10495 14702 10498
rect 14418 10449 14702 10495
rect 14418 10446 14430 10449
rect 14690 10446 14702 10449
rect 14754 10446 14766 10498
rect 15822 10434 15874 10446
rect 22430 10498 22482 10510
rect 22430 10434 22482 10446
rect 22878 10498 22930 10510
rect 31938 10446 31950 10498
rect 32002 10446 32014 10498
rect 22878 10434 22930 10446
rect 12910 10386 12962 10398
rect 12910 10322 12962 10334
rect 13246 10386 13298 10398
rect 13246 10322 13298 10334
rect 20750 10386 20802 10398
rect 46846 10386 46898 10398
rect 39218 10334 39230 10386
rect 39282 10334 39294 10386
rect 20750 10322 20802 10334
rect 46846 10322 46898 10334
rect 1344 10218 48720 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48720 10218
rect 1344 10132 48720 10166
rect 3838 10050 3890 10062
rect 3838 9986 3890 9998
rect 7982 10050 8034 10062
rect 14030 10050 14082 10062
rect 12338 9998 12350 10050
rect 12402 10047 12414 10050
rect 12562 10047 12574 10050
rect 12402 10001 12574 10047
rect 12402 9998 12414 10001
rect 12562 9998 12574 10001
rect 12626 9998 12638 10050
rect 7982 9986 8034 9998
rect 14030 9986 14082 9998
rect 14366 10050 14418 10062
rect 14366 9986 14418 9998
rect 22430 10050 22482 10062
rect 29486 10050 29538 10062
rect 29138 9998 29150 10050
rect 29202 9998 29214 10050
rect 22430 9986 22482 9998
rect 29486 9986 29538 9998
rect 33630 10050 33682 10062
rect 33630 9986 33682 9998
rect 33854 10050 33906 10062
rect 33854 9986 33906 9998
rect 12686 9938 12738 9950
rect 29710 9938 29762 9950
rect 22642 9886 22654 9938
rect 22706 9886 22718 9938
rect 24882 9886 24894 9938
rect 24946 9886 24958 9938
rect 27010 9886 27022 9938
rect 27074 9886 27086 9938
rect 12686 9874 12738 9886
rect 29710 9874 29762 9886
rect 35086 9938 35138 9950
rect 37998 9938 38050 9950
rect 44942 9938 44994 9950
rect 35858 9886 35870 9938
rect 35922 9886 35934 9938
rect 39106 9886 39118 9938
rect 39170 9886 39182 9938
rect 48290 9886 48302 9938
rect 48354 9886 48366 9938
rect 35086 9874 35138 9886
rect 37998 9874 38050 9886
rect 44942 9874 44994 9886
rect 10894 9826 10946 9838
rect 4498 9774 4510 9826
rect 4562 9774 4574 9826
rect 10894 9762 10946 9774
rect 13582 9826 13634 9838
rect 21534 9826 21586 9838
rect 32398 9826 32450 9838
rect 21298 9774 21310 9826
rect 21362 9774 21374 9826
rect 21970 9774 21982 9826
rect 22034 9774 22046 9826
rect 24098 9774 24110 9826
rect 24162 9774 24174 9826
rect 27906 9774 27918 9826
rect 27970 9774 27982 9826
rect 31042 9774 31054 9826
rect 31106 9774 31118 9826
rect 31378 9774 31390 9826
rect 31442 9774 31454 9826
rect 13582 9762 13634 9774
rect 21534 9762 21586 9774
rect 32398 9762 32450 9774
rect 33070 9826 33122 9838
rect 33070 9762 33122 9774
rect 33182 9826 33234 9838
rect 37102 9826 37154 9838
rect 33394 9774 33406 9826
rect 33458 9774 33470 9826
rect 35522 9774 35534 9826
rect 35586 9774 35598 9826
rect 33182 9762 33234 9774
rect 37102 9762 37154 9774
rect 37662 9826 37714 9838
rect 43486 9826 43538 9838
rect 42018 9774 42030 9826
rect 42082 9774 42094 9826
rect 45154 9774 45166 9826
rect 45218 9774 45230 9826
rect 45938 9774 45950 9826
rect 46002 9774 46014 9826
rect 37662 9762 37714 9774
rect 43486 9762 43538 9774
rect 2158 9714 2210 9726
rect 2158 9650 2210 9662
rect 2494 9714 2546 9726
rect 2494 9650 2546 9662
rect 3502 9714 3554 9726
rect 6078 9714 6130 9726
rect 4610 9662 4622 9714
rect 4674 9662 4686 9714
rect 3502 9650 3554 9662
rect 6078 9650 6130 9662
rect 6414 9714 6466 9726
rect 6414 9650 6466 9662
rect 7646 9714 7698 9726
rect 10558 9714 10610 9726
rect 8306 9662 8318 9714
rect 8370 9662 8382 9714
rect 8530 9662 8542 9714
rect 8594 9662 8606 9714
rect 7646 9650 7698 9662
rect 10558 9650 10610 9662
rect 14142 9714 14194 9726
rect 14142 9650 14194 9662
rect 15486 9714 15538 9726
rect 15486 9650 15538 9662
rect 16606 9714 16658 9726
rect 16606 9650 16658 9662
rect 17166 9714 17218 9726
rect 17166 9650 17218 9662
rect 17502 9714 17554 9726
rect 17502 9650 17554 9662
rect 18398 9714 18450 9726
rect 18398 9650 18450 9662
rect 19294 9714 19346 9726
rect 19294 9650 19346 9662
rect 21758 9714 21810 9726
rect 32846 9714 32898 9726
rect 30370 9662 30382 9714
rect 30434 9662 30446 9714
rect 31938 9662 31950 9714
rect 32002 9662 32014 9714
rect 21758 9650 21810 9662
rect 32846 9650 32898 9662
rect 33966 9714 34018 9726
rect 37214 9714 37266 9726
rect 43150 9714 43202 9726
rect 36082 9662 36094 9714
rect 36146 9662 36158 9714
rect 41234 9662 41246 9714
rect 41298 9662 41310 9714
rect 33966 9650 34018 9662
rect 37214 9650 37266 9662
rect 43150 9650 43202 9662
rect 9438 9602 9490 9614
rect 9438 9538 9490 9550
rect 11902 9602 11954 9614
rect 11902 9538 11954 9550
rect 12350 9602 12402 9614
rect 12350 9538 12402 9550
rect 14926 9602 14978 9614
rect 14926 9538 14978 9550
rect 15262 9602 15314 9614
rect 15262 9538 15314 9550
rect 15374 9602 15426 9614
rect 15374 9538 15426 9550
rect 16046 9602 16098 9614
rect 16046 9538 16098 9550
rect 16718 9602 16770 9614
rect 16718 9538 16770 9550
rect 16942 9602 16994 9614
rect 16942 9538 16994 9550
rect 18062 9602 18114 9614
rect 18062 9538 18114 9550
rect 18286 9602 18338 9614
rect 18286 9538 18338 9550
rect 18846 9602 18898 9614
rect 18846 9538 18898 9550
rect 19406 9602 19458 9614
rect 19406 9538 19458 9550
rect 19854 9602 19906 9614
rect 19854 9538 19906 9550
rect 20638 9602 20690 9614
rect 20638 9538 20690 9550
rect 21646 9602 21698 9614
rect 21646 9538 21698 9550
rect 22654 9602 22706 9614
rect 22654 9538 22706 9550
rect 23774 9602 23826 9614
rect 28590 9602 28642 9614
rect 32622 9602 32674 9614
rect 28130 9550 28142 9602
rect 28194 9550 28206 9602
rect 31490 9550 31502 9602
rect 31554 9550 31566 9602
rect 23774 9538 23826 9550
rect 28590 9538 28642 9550
rect 32622 9538 32674 9550
rect 34302 9602 34354 9614
rect 37438 9602 37490 9614
rect 34626 9550 34638 9602
rect 34690 9550 34702 9602
rect 34302 9538 34354 9550
rect 37438 9538 37490 9550
rect 37886 9602 37938 9614
rect 37886 9538 37938 9550
rect 38110 9602 38162 9614
rect 38110 9538 38162 9550
rect 38334 9602 38386 9614
rect 38334 9538 38386 9550
rect 1344 9434 48720 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48720 9434
rect 1344 9348 48720 9382
rect 11006 9266 11058 9278
rect 11006 9202 11058 9214
rect 11342 9266 11394 9278
rect 11342 9202 11394 9214
rect 14478 9266 14530 9278
rect 14478 9202 14530 9214
rect 14702 9266 14754 9278
rect 14702 9202 14754 9214
rect 17614 9266 17666 9278
rect 17614 9202 17666 9214
rect 19070 9266 19122 9278
rect 19070 9202 19122 9214
rect 19294 9266 19346 9278
rect 19294 9202 19346 9214
rect 19406 9266 19458 9278
rect 19406 9202 19458 9214
rect 34302 9266 34354 9278
rect 34302 9202 34354 9214
rect 34862 9266 34914 9278
rect 34862 9202 34914 9214
rect 39454 9266 39506 9278
rect 39454 9202 39506 9214
rect 6302 9154 6354 9166
rect 17838 9154 17890 9166
rect 21534 9154 21586 9166
rect 4386 9102 4398 9154
rect 4450 9102 4462 9154
rect 8418 9102 8430 9154
rect 8482 9102 8494 9154
rect 15026 9102 15038 9154
rect 15090 9102 15102 9154
rect 18162 9102 18174 9154
rect 18226 9102 18238 9154
rect 19842 9102 19854 9154
rect 19906 9102 19918 9154
rect 6302 9090 6354 9102
rect 17838 9090 17890 9102
rect 21534 9090 21586 9102
rect 21646 9154 21698 9166
rect 21646 9090 21698 9102
rect 24670 9154 24722 9166
rect 24670 9090 24722 9102
rect 25230 9154 25282 9166
rect 25230 9090 25282 9102
rect 25678 9154 25730 9166
rect 33630 9154 33682 9166
rect 45950 9154 46002 9166
rect 32162 9102 32174 9154
rect 32226 9102 32238 9154
rect 37538 9102 37550 9154
rect 37602 9102 37614 9154
rect 25678 9090 25730 9102
rect 33630 9090 33682 9102
rect 45950 9090 46002 9102
rect 3726 9042 3778 9054
rect 6638 9042 6690 9054
rect 4498 8990 4510 9042
rect 4562 8990 4574 9042
rect 3726 8978 3778 8990
rect 6638 8978 6690 8990
rect 7422 9042 7474 9054
rect 7422 8978 7474 8990
rect 7758 9042 7810 9054
rect 17278 9042 17330 9054
rect 8306 8990 8318 9042
rect 8370 8990 8382 9042
rect 12562 8990 12574 9042
rect 12626 8990 12638 9042
rect 16146 8990 16158 9042
rect 16210 8990 16222 9042
rect 7758 8978 7810 8990
rect 17278 8978 17330 8990
rect 18510 9042 18562 9054
rect 19182 9042 19234 9054
rect 22990 9042 23042 9054
rect 27582 9042 27634 9054
rect 18834 8990 18846 9042
rect 18898 8990 18910 9042
rect 20178 8990 20190 9042
rect 20242 8990 20254 9042
rect 21186 8990 21198 9042
rect 21250 8990 21262 9042
rect 23314 8990 23326 9042
rect 23378 8990 23390 9042
rect 25442 8990 25454 9042
rect 25506 8990 25518 9042
rect 18510 8978 18562 8990
rect 19182 8978 19234 8990
rect 22990 8978 23042 8990
rect 27582 8978 27634 8990
rect 27918 9042 27970 9054
rect 27918 8978 27970 8990
rect 28478 9042 28530 9054
rect 33406 9042 33458 9054
rect 46286 9042 46338 9054
rect 28802 8990 28814 9042
rect 28866 8990 28878 9042
rect 29138 8990 29150 9042
rect 29202 8990 29214 9042
rect 32274 8990 32286 9042
rect 32338 8990 32350 9042
rect 34066 8990 34078 9042
rect 34130 8990 34142 9042
rect 38322 8990 38334 9042
rect 38386 8990 38398 9042
rect 39218 8990 39230 9042
rect 39282 8990 39294 9042
rect 28478 8978 28530 8990
rect 33406 8978 33458 8990
rect 46286 8978 46338 8990
rect 5070 8930 5122 8942
rect 5070 8866 5122 8878
rect 9662 8930 9714 8942
rect 9662 8866 9714 8878
rect 11902 8930 11954 8942
rect 11902 8866 11954 8878
rect 12126 8930 12178 8942
rect 13694 8930 13746 8942
rect 12450 8878 12462 8930
rect 12514 8878 12526 8930
rect 12126 8866 12178 8878
rect 13694 8866 13746 8878
rect 15374 8930 15426 8942
rect 16830 8930 16882 8942
rect 16482 8878 16494 8930
rect 16546 8878 16558 8930
rect 15374 8866 15426 8878
rect 16830 8866 16882 8878
rect 17502 8930 17554 8942
rect 22206 8930 22258 8942
rect 20290 8878 20302 8930
rect 20354 8878 20366 8930
rect 17502 8866 17554 8878
rect 22206 8866 22258 8878
rect 27134 8930 27186 8942
rect 33070 8930 33122 8942
rect 38782 8930 38834 8942
rect 31042 8878 31054 8930
rect 31106 8878 31118 8930
rect 35410 8878 35422 8930
rect 35474 8878 35486 8930
rect 27134 8866 27186 8878
rect 33070 8866 33122 8878
rect 38782 8866 38834 8878
rect 3390 8818 3442 8830
rect 3390 8754 3442 8766
rect 15486 8818 15538 8830
rect 15486 8754 15538 8766
rect 21646 8818 21698 8830
rect 21646 8754 21698 8766
rect 23326 8818 23378 8830
rect 23326 8754 23378 8766
rect 25790 8818 25842 8830
rect 25790 8754 25842 8766
rect 34414 8818 34466 8830
rect 34414 8754 34466 8766
rect 1344 8650 48720 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48720 8650
rect 1344 8564 48720 8598
rect 16158 8482 16210 8494
rect 16158 8418 16210 8430
rect 16494 8482 16546 8494
rect 16494 8418 16546 8430
rect 37326 8482 37378 8494
rect 37326 8418 37378 8430
rect 13694 8370 13746 8382
rect 4722 8318 4734 8370
rect 4786 8318 4798 8370
rect 8642 8318 8654 8370
rect 8706 8318 8718 8370
rect 11890 8318 11902 8370
rect 11954 8318 11966 8370
rect 13694 8306 13746 8318
rect 14590 8370 14642 8382
rect 28478 8370 28530 8382
rect 34078 8370 34130 8382
rect 37214 8370 37266 8382
rect 17378 8318 17390 8370
rect 17442 8318 17454 8370
rect 18722 8318 18734 8370
rect 18786 8318 18798 8370
rect 24210 8318 24222 8370
rect 24274 8318 24286 8370
rect 25666 8318 25678 8370
rect 25730 8318 25742 8370
rect 27906 8318 27918 8370
rect 27970 8318 27982 8370
rect 29474 8318 29486 8370
rect 29538 8318 29550 8370
rect 35186 8318 35198 8370
rect 35250 8318 35262 8370
rect 14590 8306 14642 8318
rect 28478 8306 28530 8318
rect 34078 8306 34130 8318
rect 37214 8306 37266 8318
rect 38558 8370 38610 8382
rect 38558 8306 38610 8318
rect 44942 8370 44994 8382
rect 44942 8306 44994 8318
rect 19294 8258 19346 8270
rect 34750 8258 34802 8270
rect 1698 8206 1710 8258
rect 1762 8206 1774 8258
rect 2258 8206 2270 8258
rect 2322 8206 2334 8258
rect 5730 8206 5742 8258
rect 5794 8206 5806 8258
rect 6290 8206 6302 8258
rect 6354 8206 6366 8258
rect 8978 8206 8990 8258
rect 9042 8206 9054 8258
rect 17714 8206 17726 8258
rect 17778 8206 17790 8258
rect 18834 8206 18846 8258
rect 18898 8206 18910 8258
rect 21298 8206 21310 8258
rect 21362 8206 21374 8258
rect 24882 8206 24894 8258
rect 24946 8206 24958 8258
rect 29250 8206 29262 8258
rect 29314 8206 29326 8258
rect 29810 8206 29822 8258
rect 29874 8206 29886 8258
rect 31826 8206 31838 8258
rect 31890 8206 31902 8258
rect 19294 8194 19346 8206
rect 34750 8194 34802 8206
rect 35758 8258 35810 8270
rect 41570 8206 41582 8258
rect 41634 8206 41646 8258
rect 45154 8206 45166 8258
rect 45218 8206 45230 8258
rect 45938 8206 45950 8258
rect 46002 8206 46014 8258
rect 35758 8194 35810 8206
rect 12574 8146 12626 8158
rect 9762 8094 9774 8146
rect 9826 8094 9838 8146
rect 12574 8082 12626 8094
rect 12798 8146 12850 8158
rect 12798 8082 12850 8094
rect 13582 8146 13634 8158
rect 13582 8082 13634 8094
rect 15262 8146 15314 8158
rect 15262 8082 15314 8094
rect 16382 8146 16434 8158
rect 16382 8082 16434 8094
rect 18174 8146 18226 8158
rect 18174 8082 18226 8094
rect 18510 8146 18562 8158
rect 20190 8146 20242 8158
rect 30382 8146 30434 8158
rect 19618 8094 19630 8146
rect 19682 8094 19694 8146
rect 22082 8094 22094 8146
rect 22146 8094 22158 8146
rect 18510 8082 18562 8094
rect 20190 8082 20242 8094
rect 30382 8082 30434 8094
rect 32398 8146 32450 8158
rect 32398 8082 32450 8094
rect 40574 8146 40626 8158
rect 40574 8082 40626 8094
rect 12686 8034 12738 8046
rect 12686 7970 12738 7982
rect 14030 8034 14082 8046
rect 20526 8034 20578 8046
rect 36206 8034 36258 8046
rect 15586 7982 15598 8034
rect 15650 7982 15662 8034
rect 29922 7982 29934 8034
rect 29986 7982 29998 8034
rect 14030 7970 14082 7982
rect 20526 7970 20578 7982
rect 36206 7970 36258 7982
rect 37886 8034 37938 8046
rect 37886 7970 37938 7982
rect 41358 8034 41410 8046
rect 41358 7970 41410 7982
rect 42478 8034 42530 8046
rect 48290 7982 48302 8034
rect 48354 7982 48366 8034
rect 42478 7970 42530 7982
rect 1344 7866 48720 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48720 7866
rect 1344 7780 48720 7814
rect 2158 7698 2210 7710
rect 2158 7634 2210 7646
rect 4286 7698 4338 7710
rect 4286 7634 4338 7646
rect 5630 7698 5682 7710
rect 5630 7634 5682 7646
rect 6078 7698 6130 7710
rect 6078 7634 6130 7646
rect 7758 7698 7810 7710
rect 7758 7634 7810 7646
rect 8206 7698 8258 7710
rect 8206 7634 8258 7646
rect 10110 7698 10162 7710
rect 16718 7698 16770 7710
rect 16370 7646 16382 7698
rect 16434 7646 16446 7698
rect 10110 7634 10162 7646
rect 16718 7634 16770 7646
rect 20414 7698 20466 7710
rect 20414 7634 20466 7646
rect 21310 7698 21362 7710
rect 21310 7634 21362 7646
rect 23662 7698 23714 7710
rect 23662 7634 23714 7646
rect 24110 7698 24162 7710
rect 24110 7634 24162 7646
rect 24558 7698 24610 7710
rect 32510 7698 32562 7710
rect 29810 7646 29822 7698
rect 29874 7646 29886 7698
rect 30818 7646 30830 7698
rect 30882 7646 30894 7698
rect 24558 7634 24610 7646
rect 32510 7634 32562 7646
rect 33294 7698 33346 7710
rect 33294 7634 33346 7646
rect 34638 7698 34690 7710
rect 34638 7634 34690 7646
rect 34974 7698 35026 7710
rect 34974 7634 35026 7646
rect 35534 7698 35586 7710
rect 35534 7634 35586 7646
rect 35870 7698 35922 7710
rect 35870 7634 35922 7646
rect 36654 7698 36706 7710
rect 41246 7698 41298 7710
rect 46510 7698 46562 7710
rect 38098 7646 38110 7698
rect 38162 7646 38174 7698
rect 43810 7646 43822 7698
rect 43874 7646 43886 7698
rect 36654 7634 36706 7646
rect 41246 7634 41298 7646
rect 46510 7634 46562 7646
rect 2494 7586 2546 7598
rect 2494 7522 2546 7534
rect 11230 7586 11282 7598
rect 11230 7522 11282 7534
rect 11342 7586 11394 7598
rect 17950 7586 18002 7598
rect 12786 7534 12798 7586
rect 12850 7534 12862 7586
rect 13570 7534 13582 7586
rect 13634 7534 13646 7586
rect 15586 7534 15598 7586
rect 15650 7534 15662 7586
rect 11342 7522 11394 7534
rect 17950 7522 18002 7534
rect 20638 7586 20690 7598
rect 20638 7522 20690 7534
rect 20974 7586 21026 7598
rect 28142 7586 28194 7598
rect 34078 7586 34130 7598
rect 44270 7586 44322 7598
rect 21970 7534 21982 7586
rect 22034 7534 22046 7586
rect 29250 7534 29262 7586
rect 29314 7534 29326 7586
rect 29698 7534 29710 7586
rect 29762 7534 29774 7586
rect 32162 7534 32174 7586
rect 32226 7534 32238 7586
rect 42354 7534 42366 7586
rect 42418 7534 42430 7586
rect 47170 7534 47182 7586
rect 47234 7534 47246 7586
rect 47618 7534 47630 7586
rect 47682 7534 47694 7586
rect 20974 7522 21026 7534
rect 28142 7522 28194 7534
rect 34078 7522 34130 7534
rect 44270 7522 44322 7534
rect 10446 7474 10498 7486
rect 10446 7410 10498 7422
rect 11006 7474 11058 7486
rect 11006 7410 11058 7422
rect 11790 7474 11842 7486
rect 11790 7410 11842 7422
rect 12126 7474 12178 7486
rect 13918 7474 13970 7486
rect 12898 7422 12910 7474
rect 12962 7422 12974 7474
rect 12126 7410 12178 7422
rect 13918 7410 13970 7422
rect 18174 7474 18226 7486
rect 18174 7410 18226 7422
rect 18510 7474 18562 7486
rect 18510 7410 18562 7422
rect 18846 7474 18898 7486
rect 18846 7410 18898 7422
rect 19182 7474 19234 7486
rect 26910 7474 26962 7486
rect 25666 7422 25678 7474
rect 25730 7422 25742 7474
rect 26450 7422 26462 7474
rect 26514 7422 26526 7474
rect 19182 7410 19234 7422
rect 26910 7410 26962 7422
rect 27470 7474 27522 7486
rect 27470 7410 27522 7422
rect 27694 7474 27746 7486
rect 27694 7410 27746 7422
rect 28366 7474 28418 7486
rect 38782 7474 38834 7486
rect 29026 7422 29038 7474
rect 29090 7422 29102 7474
rect 30706 7422 30718 7474
rect 30770 7422 30782 7474
rect 30930 7422 30942 7474
rect 30994 7422 31006 7474
rect 31490 7422 31502 7474
rect 31554 7422 31566 7474
rect 37538 7422 37550 7474
rect 37602 7422 37614 7474
rect 37874 7422 37886 7474
rect 37938 7422 37950 7474
rect 39330 7422 39342 7474
rect 39394 7422 39406 7474
rect 40226 7422 40238 7474
rect 40290 7422 40302 7474
rect 42018 7422 42030 7474
rect 42082 7422 42094 7474
rect 43138 7422 43150 7474
rect 43202 7422 43214 7474
rect 43586 7422 43598 7474
rect 43650 7422 43662 7474
rect 45042 7422 45054 7474
rect 45106 7422 45118 7474
rect 45938 7422 45950 7474
rect 46002 7422 46014 7474
rect 28366 7410 28418 7422
rect 38782 7410 38834 7422
rect 4734 7362 4786 7374
rect 4734 7298 4786 7310
rect 5070 7362 5122 7374
rect 5070 7298 5122 7310
rect 6526 7362 6578 7374
rect 6526 7298 6578 7310
rect 7198 7362 7250 7374
rect 7198 7298 7250 7310
rect 8542 7362 8594 7374
rect 8542 7298 8594 7310
rect 9102 7362 9154 7374
rect 9102 7298 9154 7310
rect 9774 7362 9826 7374
rect 18398 7362 18450 7374
rect 14578 7310 14590 7362
rect 14642 7310 14654 7362
rect 9774 7298 9826 7310
rect 18398 7298 18450 7310
rect 19742 7362 19794 7374
rect 27918 7362 27970 7374
rect 20402 7310 20414 7362
rect 20466 7310 20478 7362
rect 22978 7310 22990 7362
rect 23042 7310 23054 7362
rect 25890 7310 25902 7362
rect 25954 7310 25966 7362
rect 19742 7298 19794 7310
rect 27918 7298 27970 7310
rect 33630 7362 33682 7374
rect 33630 7298 33682 7310
rect 37102 7362 37154 7374
rect 37102 7298 37154 7310
rect 42814 7362 42866 7374
rect 42814 7298 42866 7310
rect 48190 7362 48242 7374
rect 48190 7298 48242 7310
rect 17390 7250 17442 7262
rect 7858 7198 7870 7250
rect 7922 7247 7934 7250
rect 8418 7247 8430 7250
rect 7922 7201 8430 7247
rect 7922 7198 7934 7201
rect 8418 7198 8430 7201
rect 8482 7198 8494 7250
rect 17390 7186 17442 7198
rect 17726 7250 17778 7262
rect 41582 7250 41634 7262
rect 25554 7198 25566 7250
rect 25618 7198 25630 7250
rect 17726 7186 17778 7198
rect 41582 7186 41634 7198
rect 46846 7250 46898 7262
rect 46846 7186 46898 7198
rect 1344 7082 48720 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48720 7082
rect 1344 6996 48720 7030
rect 3950 6914 4002 6926
rect 3950 6850 4002 6862
rect 7870 6914 7922 6926
rect 7870 6850 7922 6862
rect 12574 6914 12626 6926
rect 12574 6850 12626 6862
rect 15150 6914 15202 6926
rect 15150 6850 15202 6862
rect 15486 6914 15538 6926
rect 15486 6850 15538 6862
rect 18286 6914 18338 6926
rect 18286 6850 18338 6862
rect 35534 6914 35586 6926
rect 35534 6850 35586 6862
rect 46958 6914 47010 6926
rect 46958 6850 47010 6862
rect 6078 6802 6130 6814
rect 6078 6738 6130 6750
rect 15598 6802 15650 6814
rect 29822 6802 29874 6814
rect 16146 6750 16158 6802
rect 16210 6750 16222 6802
rect 18946 6750 18958 6802
rect 19010 6750 19022 6802
rect 23986 6750 23998 6802
rect 24050 6750 24062 6802
rect 15598 6738 15650 6750
rect 29822 6738 29874 6750
rect 31278 6802 31330 6814
rect 34738 6750 34750 6802
rect 34802 6750 34814 6802
rect 31278 6738 31330 6750
rect 9886 6690 9938 6702
rect 4722 6638 4734 6690
rect 4786 6638 4798 6690
rect 9886 6626 9938 6638
rect 10670 6690 10722 6702
rect 10670 6626 10722 6638
rect 11006 6690 11058 6702
rect 11006 6626 11058 6638
rect 12798 6690 12850 6702
rect 12798 6626 12850 6638
rect 13918 6690 13970 6702
rect 13918 6626 13970 6638
rect 15262 6690 15314 6702
rect 15262 6626 15314 6638
rect 18062 6690 18114 6702
rect 22206 6690 22258 6702
rect 18610 6638 18622 6690
rect 18674 6638 18686 6690
rect 21522 6638 21534 6690
rect 21586 6638 21598 6690
rect 18062 6626 18114 6638
rect 22206 6626 22258 6638
rect 23214 6690 23266 6702
rect 23214 6626 23266 6638
rect 26014 6690 26066 6702
rect 26014 6626 26066 6638
rect 28142 6690 28194 6702
rect 28142 6626 28194 6638
rect 28366 6690 28418 6702
rect 28366 6626 28418 6638
rect 29150 6690 29202 6702
rect 29150 6626 29202 6638
rect 29262 6690 29314 6702
rect 29262 6626 29314 6638
rect 29598 6690 29650 6702
rect 37214 6690 37266 6702
rect 31938 6638 31950 6690
rect 32002 6638 32014 6690
rect 32610 6638 32622 6690
rect 32674 6638 32686 6690
rect 36082 6638 36094 6690
rect 36146 6638 36158 6690
rect 29598 6626 29650 6638
rect 37214 6626 37266 6638
rect 37550 6690 37602 6702
rect 37550 6626 37602 6638
rect 37998 6690 38050 6702
rect 37998 6626 38050 6638
rect 40350 6690 40402 6702
rect 45054 6690 45106 6702
rect 40786 6638 40798 6690
rect 40850 6638 40862 6690
rect 41346 6638 41358 6690
rect 41410 6638 41422 6690
rect 43698 6638 43710 6690
rect 43762 6638 43774 6690
rect 40350 6626 40402 6638
rect 45054 6626 45106 6638
rect 45502 6690 45554 6702
rect 45502 6626 45554 6638
rect 1934 6578 1986 6590
rect 6750 6578 6802 6590
rect 4498 6526 4510 6578
rect 4562 6526 4574 6578
rect 1934 6514 1986 6526
rect 6750 6514 6802 6526
rect 7534 6578 7586 6590
rect 27806 6578 27858 6590
rect 30494 6578 30546 6590
rect 38558 6578 38610 6590
rect 8082 6526 8094 6578
rect 8146 6526 8158 6578
rect 8530 6526 8542 6578
rect 8594 6526 8606 6578
rect 10210 6526 10222 6578
rect 10274 6526 10286 6578
rect 11218 6526 11230 6578
rect 11282 6526 11294 6578
rect 11554 6526 11566 6578
rect 11618 6526 11630 6578
rect 14130 6526 14142 6578
rect 14194 6526 14206 6578
rect 14466 6526 14478 6578
rect 14530 6526 14542 6578
rect 17154 6526 17166 6578
rect 17218 6526 17230 6578
rect 20290 6526 20302 6578
rect 20354 6526 20366 6578
rect 21410 6526 21422 6578
rect 21474 6526 21486 6578
rect 24994 6526 25006 6578
rect 25058 6526 25070 6578
rect 26562 6526 26574 6578
rect 26626 6526 26638 6578
rect 26786 6526 26798 6578
rect 26850 6526 26862 6578
rect 30146 6526 30158 6578
rect 30210 6526 30222 6578
rect 36306 6526 36318 6578
rect 36370 6526 36382 6578
rect 7534 6514 7586 6526
rect 27806 6514 27858 6526
rect 30494 6514 30546 6526
rect 38558 6514 38610 6526
rect 46174 6578 46226 6590
rect 46174 6514 46226 6526
rect 46622 6578 46674 6590
rect 47170 6526 47182 6578
rect 47234 6526 47246 6578
rect 47506 6526 47518 6578
rect 47570 6526 47582 6578
rect 46622 6514 46674 6526
rect 2830 6466 2882 6478
rect 2830 6402 2882 6414
rect 3278 6466 3330 6478
rect 3278 6402 3330 6414
rect 3614 6466 3666 6478
rect 3614 6402 3666 6414
rect 6414 6466 6466 6478
rect 9550 6466 9602 6478
rect 13582 6466 13634 6478
rect 9202 6414 9214 6466
rect 9266 6414 9278 6466
rect 12226 6414 12238 6466
rect 12290 6414 12302 6466
rect 6414 6402 6466 6414
rect 9550 6402 9602 6414
rect 13582 6402 13634 6414
rect 22542 6466 22594 6478
rect 22542 6402 22594 6414
rect 23774 6466 23826 6478
rect 28030 6466 28082 6478
rect 26114 6414 26126 6466
rect 26178 6414 26190 6466
rect 23774 6402 23826 6414
rect 28030 6402 28082 6414
rect 30830 6466 30882 6478
rect 30830 6402 30882 6414
rect 35198 6466 35250 6478
rect 35198 6402 35250 6414
rect 39006 6466 39058 6478
rect 39006 6402 39058 6414
rect 39790 6466 39842 6478
rect 39790 6402 39842 6414
rect 45838 6466 45890 6478
rect 45838 6402 45890 6414
rect 1344 6298 48720 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48720 6298
rect 1344 6212 48720 6246
rect 5182 6130 5234 6142
rect 24222 6130 24274 6142
rect 4722 6078 4734 6130
rect 4786 6078 4798 6130
rect 8642 6078 8654 6130
rect 8706 6078 8718 6130
rect 17714 6078 17726 6130
rect 17778 6078 17790 6130
rect 5182 6066 5234 6078
rect 24222 6066 24274 6078
rect 24446 6130 24498 6142
rect 24446 6066 24498 6078
rect 24670 6130 24722 6142
rect 24670 6066 24722 6078
rect 25342 6130 25394 6142
rect 25342 6066 25394 6078
rect 25566 6130 25618 6142
rect 33742 6130 33794 6142
rect 26338 6078 26350 6130
rect 26402 6078 26414 6130
rect 27234 6078 27246 6130
rect 27298 6078 27310 6130
rect 25566 6066 25618 6078
rect 33742 6066 33794 6078
rect 38222 6130 38274 6142
rect 38222 6066 38274 6078
rect 38670 6130 38722 6142
rect 38670 6066 38722 6078
rect 44942 6130 44994 6142
rect 44942 6066 44994 6078
rect 45390 6130 45442 6142
rect 45390 6066 45442 6078
rect 9774 6018 9826 6030
rect 9774 5954 9826 5966
rect 9998 6018 10050 6030
rect 9998 5954 10050 5966
rect 10670 6018 10722 6030
rect 15038 6018 15090 6030
rect 23550 6018 23602 6030
rect 11778 5966 11790 6018
rect 11842 5966 11854 6018
rect 16370 5966 16382 6018
rect 16434 5966 16446 6018
rect 18386 5966 18398 6018
rect 18450 5966 18462 6018
rect 18722 5966 18734 6018
rect 18786 5966 18798 6018
rect 20514 5966 20526 6018
rect 20578 5966 20590 6018
rect 10670 5954 10722 5966
rect 15038 5954 15090 5966
rect 23550 5954 23602 5966
rect 25230 6018 25282 6030
rect 37438 6018 37490 6030
rect 41470 6018 41522 6030
rect 28242 5966 28254 6018
rect 28306 5966 28318 6018
rect 31714 5966 31726 6018
rect 31778 5966 31790 6018
rect 39666 5966 39678 6018
rect 39730 5966 39742 6018
rect 40226 5966 40238 6018
rect 40290 5966 40302 6018
rect 43138 5966 43150 6018
rect 43202 5966 43214 6018
rect 25230 5954 25282 5966
rect 37438 5954 37490 5966
rect 41470 5954 41522 5966
rect 17390 5906 17442 5918
rect 23214 5906 23266 5918
rect 1698 5854 1710 5906
rect 1762 5854 1774 5906
rect 2258 5854 2270 5906
rect 2322 5854 2334 5906
rect 5730 5854 5742 5906
rect 5794 5854 5806 5906
rect 6290 5854 6302 5906
rect 6354 5854 6366 5906
rect 10434 5854 10446 5906
rect 10498 5854 10510 5906
rect 10994 5854 11006 5906
rect 11058 5854 11070 5906
rect 14802 5854 14814 5906
rect 14866 5854 14878 5906
rect 19730 5854 19742 5906
rect 19794 5854 19806 5906
rect 22978 5854 22990 5906
rect 23042 5854 23054 5906
rect 17390 5842 17442 5854
rect 23214 5842 23266 5854
rect 23438 5906 23490 5918
rect 23438 5842 23490 5854
rect 25790 5906 25842 5918
rect 25790 5842 25842 5854
rect 26910 5906 26962 5918
rect 39454 5906 39506 5918
rect 43710 5906 43762 5918
rect 28354 5854 28366 5906
rect 28418 5854 28430 5906
rect 32498 5854 32510 5906
rect 32562 5854 32574 5906
rect 33506 5854 33518 5906
rect 33570 5854 33582 5906
rect 34066 5854 34078 5906
rect 34130 5854 34142 5906
rect 34626 5854 34638 5906
rect 34690 5854 34702 5906
rect 37650 5854 37662 5906
rect 37714 5854 37726 5906
rect 42914 5854 42926 5906
rect 42978 5854 42990 5906
rect 45714 5854 45726 5906
rect 45778 5854 45790 5906
rect 26910 5842 26962 5854
rect 39454 5842 39506 5854
rect 43710 5842 43762 5854
rect 14366 5794 14418 5806
rect 24558 5794 24610 5806
rect 9650 5742 9662 5794
rect 9714 5742 9726 5794
rect 13906 5742 13918 5794
rect 13970 5742 13982 5794
rect 15362 5742 15374 5794
rect 15426 5742 15438 5794
rect 22642 5742 22654 5794
rect 22706 5742 22718 5794
rect 14366 5730 14418 5742
rect 24558 5730 24610 5742
rect 26014 5794 26066 5806
rect 26014 5730 26066 5742
rect 26686 5794 26738 5806
rect 41022 5794 41074 5806
rect 29586 5742 29598 5794
rect 29650 5742 29662 5794
rect 37090 5742 37102 5794
rect 37154 5742 37166 5794
rect 26686 5730 26738 5742
rect 41022 5730 41074 5742
rect 42142 5794 42194 5806
rect 46834 5742 46846 5794
rect 46898 5742 46910 5794
rect 42142 5730 42194 5742
rect 18958 5682 19010 5694
rect 18958 5618 19010 5630
rect 19294 5682 19346 5694
rect 19294 5618 19346 5630
rect 28814 5682 28866 5694
rect 28814 5618 28866 5630
rect 29150 5682 29202 5694
rect 29150 5618 29202 5630
rect 39118 5682 39170 5694
rect 39118 5618 39170 5630
rect 44046 5682 44098 5694
rect 44046 5618 44098 5630
rect 1344 5514 48720 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48720 5514
rect 1344 5428 48720 5462
rect 4174 5346 4226 5358
rect 12686 5346 12738 5358
rect 12338 5294 12350 5346
rect 12402 5294 12414 5346
rect 4174 5282 4226 5294
rect 12686 5282 12738 5294
rect 29598 5346 29650 5358
rect 29598 5282 29650 5294
rect 31054 5346 31106 5358
rect 31054 5282 31106 5294
rect 37662 5346 37714 5358
rect 37662 5282 37714 5294
rect 37998 5346 38050 5358
rect 37998 5282 38050 5294
rect 1822 5234 1874 5246
rect 1822 5170 1874 5182
rect 3054 5234 3106 5246
rect 3054 5170 3106 5182
rect 3502 5234 3554 5246
rect 3502 5170 3554 5182
rect 5742 5234 5794 5246
rect 20750 5234 20802 5246
rect 9538 5182 9550 5234
rect 9602 5182 9614 5234
rect 11666 5182 11678 5234
rect 11730 5182 11742 5234
rect 15138 5182 15150 5234
rect 15202 5182 15214 5234
rect 16258 5182 16270 5234
rect 16322 5182 16334 5234
rect 18386 5182 18398 5234
rect 18450 5182 18462 5234
rect 18722 5182 18734 5234
rect 18786 5182 18798 5234
rect 5742 5170 5794 5182
rect 20750 5170 20802 5182
rect 24894 5234 24946 5246
rect 35534 5234 35586 5246
rect 31714 5182 31726 5234
rect 31778 5182 31790 5234
rect 24894 5170 24946 5182
rect 35534 5170 35586 5182
rect 35982 5234 36034 5246
rect 35982 5170 36034 5182
rect 36430 5234 36482 5246
rect 36430 5170 36482 5182
rect 36990 5234 37042 5246
rect 36990 5170 37042 5182
rect 43262 5234 43314 5246
rect 43262 5170 43314 5182
rect 44830 5234 44882 5246
rect 48290 5182 48302 5234
rect 48354 5182 48366 5234
rect 44830 5170 44882 5182
rect 2494 5122 2546 5134
rect 2494 5058 2546 5070
rect 3838 5122 3890 5134
rect 6414 5122 6466 5134
rect 4834 5070 4846 5122
rect 4898 5070 4910 5122
rect 3838 5058 3890 5070
rect 6414 5058 6466 5070
rect 7086 5122 7138 5134
rect 12910 5122 12962 5134
rect 21422 5122 21474 5134
rect 27582 5122 27634 5134
rect 7522 5070 7534 5122
rect 7586 5070 7598 5122
rect 8194 5070 8206 5122
rect 8258 5070 8270 5122
rect 8866 5070 8878 5122
rect 8930 5070 8942 5122
rect 15474 5070 15486 5122
rect 15538 5070 15550 5122
rect 22082 5070 22094 5122
rect 22146 5070 22158 5122
rect 27234 5070 27246 5122
rect 27298 5070 27310 5122
rect 7086 5058 7138 5070
rect 12910 5058 12962 5070
rect 21422 5058 21474 5070
rect 27582 5058 27634 5070
rect 28590 5122 28642 5134
rect 28590 5058 28642 5070
rect 29262 5122 29314 5134
rect 30830 5122 30882 5134
rect 35086 5122 35138 5134
rect 42142 5122 42194 5134
rect 30034 5070 30046 5122
rect 30098 5070 30110 5122
rect 34626 5070 34638 5122
rect 34690 5070 34702 5122
rect 38546 5070 38558 5122
rect 38610 5070 38622 5122
rect 39218 5070 39230 5122
rect 39282 5070 39294 5122
rect 43698 5070 43710 5122
rect 43762 5070 43774 5122
rect 45154 5070 45166 5122
rect 45218 5070 45230 5122
rect 45826 5070 45838 5122
rect 45890 5070 45902 5122
rect 29262 5058 29314 5070
rect 30830 5058 30882 5070
rect 35086 5058 35138 5070
rect 42142 5058 42194 5070
rect 2158 5010 2210 5022
rect 28254 5010 28306 5022
rect 4722 4958 4734 5010
rect 4786 4958 4798 5010
rect 8418 4958 8430 5010
rect 8482 4958 8494 5010
rect 14130 4958 14142 5010
rect 14194 4958 14206 5010
rect 19730 4958 19742 5010
rect 19794 4958 19806 5010
rect 30258 4958 30270 5010
rect 30322 4958 30334 5010
rect 33842 4958 33854 5010
rect 33906 4958 33918 5010
rect 38770 4958 38782 5010
rect 38834 4958 38846 5010
rect 2158 4946 2210 4958
rect 28254 4946 28306 4958
rect 6078 4898 6130 4910
rect 6078 4834 6130 4846
rect 6750 4898 6802 4910
rect 6750 4834 6802 4846
rect 7758 4898 7810 4910
rect 7758 4834 7810 4846
rect 22766 4898 22818 4910
rect 22766 4834 22818 4846
rect 27918 4898 27970 4910
rect 37102 4898 37154 4910
rect 31378 4846 31390 4898
rect 31442 4846 31454 4898
rect 27918 4834 27970 4846
rect 37102 4834 37154 4846
rect 40238 4898 40290 4910
rect 40238 4834 40290 4846
rect 42478 4898 42530 4910
rect 42478 4834 42530 4846
rect 43934 4898 43986 4910
rect 43934 4834 43986 4846
rect 1344 4730 48720 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48720 4730
rect 1344 4644 48720 4678
rect 5742 4562 5794 4574
rect 4834 4510 4846 4562
rect 4898 4510 4910 4562
rect 5742 4498 5794 4510
rect 18174 4562 18226 4574
rect 18174 4498 18226 4510
rect 20750 4562 20802 4574
rect 20750 4498 20802 4510
rect 34078 4562 34130 4574
rect 39554 4510 39566 4562
rect 39618 4510 39630 4562
rect 40898 4510 40910 4562
rect 40962 4510 40974 4562
rect 47282 4510 47294 4562
rect 47346 4510 47358 4562
rect 34078 4498 34130 4510
rect 17390 4450 17442 4462
rect 6850 4398 6862 4450
rect 6914 4398 6926 4450
rect 10546 4398 10558 4450
rect 10610 4398 10622 4450
rect 13570 4398 13582 4450
rect 13634 4398 13646 4450
rect 14466 4398 14478 4450
rect 14530 4398 14542 4450
rect 17390 4386 17442 4398
rect 17502 4450 17554 4462
rect 17502 4386 17554 4398
rect 17726 4450 17778 4462
rect 17726 4386 17778 4398
rect 18510 4450 18562 4462
rect 21310 4450 21362 4462
rect 33070 4450 33122 4462
rect 19058 4398 19070 4450
rect 19122 4398 19134 4450
rect 22530 4398 22542 4450
rect 22594 4398 22606 4450
rect 25890 4398 25902 4450
rect 25954 4398 25966 4450
rect 26226 4398 26238 4450
rect 26290 4398 26302 4450
rect 18510 4386 18562 4398
rect 21310 4386 21362 4398
rect 33070 4386 33122 4398
rect 33742 4450 33794 4462
rect 33742 4386 33794 4398
rect 34414 4450 34466 4462
rect 34414 4386 34466 4398
rect 34862 4450 34914 4462
rect 34862 4386 34914 4398
rect 35870 4450 35922 4462
rect 35870 4386 35922 4398
rect 40014 4450 40066 4462
rect 40014 4386 40066 4398
rect 40350 4450 40402 4462
rect 40350 4386 40402 4398
rect 17838 4338 17890 4350
rect 1698 4286 1710 4338
rect 1762 4286 1774 4338
rect 2370 4286 2382 4338
rect 2434 4286 2446 4338
rect 5506 4286 5518 4338
rect 5570 4286 5582 4338
rect 6066 4286 6078 4338
rect 6130 4286 6142 4338
rect 10210 4286 10222 4338
rect 10274 4286 10286 4338
rect 11106 4286 11118 4338
rect 11170 4286 11182 4338
rect 17838 4274 17890 4286
rect 18174 4338 18226 4350
rect 21858 4286 21870 4338
rect 21922 4286 21934 4338
rect 26898 4286 26910 4338
rect 26962 4286 26974 4338
rect 31938 4286 31950 4338
rect 32002 4286 32014 4338
rect 33282 4286 33294 4338
rect 33346 4286 33358 4338
rect 36418 4286 36430 4338
rect 36482 4286 36494 4338
rect 37202 4286 37214 4338
rect 37266 4286 37278 4338
rect 43250 4286 43262 4338
rect 43314 4286 43326 4338
rect 43810 4286 43822 4338
rect 43874 4286 43886 4338
rect 44146 4286 44158 4338
rect 44210 4286 44222 4338
rect 44818 4286 44830 4338
rect 44882 4286 44894 4338
rect 18174 4274 18226 4286
rect 16606 4226 16658 4238
rect 25678 4226 25730 4238
rect 8978 4174 8990 4226
rect 9042 4174 9054 4226
rect 10658 4174 10670 4226
rect 10722 4174 10734 4226
rect 20178 4174 20190 4226
rect 20242 4174 20254 4226
rect 24658 4174 24670 4226
rect 24722 4174 24734 4226
rect 16606 4162 16658 4174
rect 25678 4162 25730 4174
rect 11454 4114 11506 4126
rect 11454 4050 11506 4062
rect 25342 4114 25394 4126
rect 25342 4050 25394 4062
rect 27918 4114 27970 4126
rect 27918 4050 27970 4062
rect 30046 4114 30098 4126
rect 30046 4050 30098 4062
rect 35310 4114 35362 4126
rect 35310 4050 35362 4062
rect 35758 4114 35810 4126
rect 35758 4050 35810 4062
rect 1344 3946 48720 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48720 3946
rect 1344 3860 48720 3894
rect 16830 3778 16882 3790
rect 16830 3714 16882 3726
rect 20750 3778 20802 3790
rect 20750 3714 20802 3726
rect 21086 3778 21138 3790
rect 21086 3714 21138 3726
rect 24558 3778 24610 3790
rect 24558 3714 24610 3726
rect 24894 3778 24946 3790
rect 24894 3714 24946 3726
rect 8206 3666 8258 3678
rect 13470 3666 13522 3678
rect 9314 3614 9326 3666
rect 9378 3614 9390 3666
rect 11106 3614 11118 3666
rect 11170 3614 11182 3666
rect 8206 3602 8258 3614
rect 13470 3602 13522 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 36990 3666 37042 3678
rect 36990 3602 37042 3614
rect 40798 3666 40850 3678
rect 40798 3602 40850 3614
rect 44606 3666 44658 3678
rect 44606 3602 44658 3614
rect 46510 3666 46562 3678
rect 46510 3602 46562 3614
rect 48190 3666 48242 3678
rect 48190 3602 48242 3614
rect 3726 3554 3778 3566
rect 1810 3502 1822 3554
rect 1874 3502 1886 3554
rect 2482 3502 2494 3554
rect 2546 3502 2558 3554
rect 3154 3502 3166 3554
rect 3218 3502 3230 3554
rect 3726 3490 3778 3502
rect 4398 3554 4450 3566
rect 4398 3490 4450 3502
rect 5966 3554 6018 3566
rect 5966 3490 6018 3502
rect 6078 3554 6130 3566
rect 8766 3554 8818 3566
rect 31278 3554 31330 3566
rect 6962 3502 6974 3554
rect 7026 3502 7038 3554
rect 7634 3502 7646 3554
rect 7698 3502 7710 3554
rect 19954 3502 19966 3554
rect 20018 3502 20030 3554
rect 21410 3502 21422 3554
rect 21474 3502 21486 3554
rect 25218 3502 25230 3554
rect 25282 3502 25294 3554
rect 28354 3502 28366 3554
rect 28418 3502 28430 3554
rect 32610 3502 32622 3554
rect 32674 3502 32686 3554
rect 35186 3502 35198 3554
rect 35250 3502 35262 3554
rect 36418 3502 36430 3554
rect 36482 3502 36494 3554
rect 39778 3502 39790 3554
rect 39842 3502 39854 3554
rect 43586 3502 43598 3554
rect 43650 3502 43662 3554
rect 6078 3490 6130 3502
rect 8766 3490 8818 3502
rect 31278 3490 31330 3502
rect 2718 3442 2770 3454
rect 2718 3378 2770 3390
rect 3390 3442 3442 3454
rect 3390 3378 3442 3390
rect 4062 3442 4114 3454
rect 4062 3378 4114 3390
rect 4958 3442 5010 3454
rect 6190 3442 6242 3454
rect 5506 3390 5518 3442
rect 5570 3390 5582 3442
rect 4958 3378 5010 3390
rect 6190 3378 6242 3390
rect 7198 3442 7250 3454
rect 13582 3442 13634 3454
rect 20190 3442 20242 3454
rect 7858 3390 7870 3442
rect 7922 3390 7934 3442
rect 10658 3390 10670 3442
rect 10722 3390 10734 3442
rect 12450 3390 12462 3442
rect 12514 3390 12526 3442
rect 15698 3390 15710 3442
rect 15762 3390 15774 3442
rect 19282 3390 19294 3442
rect 19346 3390 19358 3442
rect 7198 3378 7250 3390
rect 13582 3378 13634 3390
rect 20190 3378 20242 3390
rect 20974 3442 21026 3454
rect 24782 3442 24834 3454
rect 23202 3390 23214 3442
rect 23266 3390 23278 3442
rect 20974 3378 21026 3390
rect 24782 3378 24834 3390
rect 31614 3442 31666 3454
rect 33730 3390 33742 3442
rect 33794 3390 33806 3442
rect 31614 3378 31666 3390
rect 2046 3330 2098 3342
rect 2046 3266 2098 3278
rect 26238 3330 26290 3342
rect 38894 3330 38946 3342
rect 35410 3278 35422 3330
rect 35474 3278 35486 3330
rect 26238 3266 26290 3278
rect 38894 3266 38946 3278
rect 42702 3330 42754 3342
rect 42702 3266 42754 3278
rect 47406 3330 47458 3342
rect 47406 3266 47458 3278
rect 1344 3162 48720 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48720 3162
rect 1344 3076 48720 3110
<< via1 >>
rect 27022 50318 27074 50370
rect 27918 50318 27970 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 27022 49982 27074 50034
rect 29486 49870 29538 49922
rect 32846 49870 32898 49922
rect 26798 49758 26850 49810
rect 29822 49758 29874 49810
rect 32622 49758 32674 49810
rect 21086 49646 21138 49698
rect 21534 49646 21586 49698
rect 28926 49646 28978 49698
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 14478 48974 14530 49026
rect 15038 48974 15090 49026
rect 17614 48974 17666 49026
rect 18286 48974 18338 49026
rect 21422 48974 21474 49026
rect 21870 48974 21922 49026
rect 27918 48974 27970 49026
rect 28702 48974 28754 49026
rect 29262 48974 29314 49026
rect 29710 48974 29762 49026
rect 32622 48974 32674 49026
rect 33294 48974 33346 49026
rect 37102 48974 37154 49026
rect 37550 48974 37602 49026
rect 17390 48750 17442 48802
rect 20750 48750 20802 48802
rect 24334 48750 24386 48802
rect 25566 48750 25618 48802
rect 32174 48750 32226 48802
rect 35758 48750 35810 48802
rect 36206 48750 36258 48802
rect 40014 48750 40066 48802
rect 40462 48750 40514 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 16270 48414 16322 48466
rect 17614 48414 17666 48466
rect 18174 48414 18226 48466
rect 27358 48414 27410 48466
rect 29934 48414 29986 48466
rect 33182 48414 33234 48466
rect 37550 48414 37602 48466
rect 19854 48302 19906 48354
rect 21534 48302 21586 48354
rect 21982 48302 22034 48354
rect 22654 48302 22706 48354
rect 24110 48302 24162 48354
rect 28254 48302 28306 48354
rect 30830 48302 30882 48354
rect 33742 48302 33794 48354
rect 34078 48302 34130 48354
rect 38894 48302 38946 48354
rect 39902 48302 39954 48354
rect 16606 48190 16658 48242
rect 18510 48190 18562 48242
rect 18958 48190 19010 48242
rect 20078 48190 20130 48242
rect 24446 48190 24498 48242
rect 28478 48190 28530 48242
rect 30270 48190 30322 48242
rect 30718 48190 30770 48242
rect 37326 48190 37378 48242
rect 37998 48190 38050 48242
rect 38782 48190 38834 48242
rect 39566 48190 39618 48242
rect 32398 48078 32450 48130
rect 40350 48078 40402 48130
rect 19294 47966 19346 48018
rect 20974 47966 21026 48018
rect 21310 47966 21362 48018
rect 27694 47966 27746 48018
rect 33518 47966 33570 48018
rect 38334 47966 38386 48018
rect 40126 47966 40178 48018
rect 40350 47966 40402 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 17278 47630 17330 47682
rect 38894 47630 38946 47682
rect 9998 47406 10050 47458
rect 10558 47406 10610 47458
rect 17614 47406 17666 47458
rect 18398 47406 18450 47458
rect 21310 47406 21362 47458
rect 23214 47406 23266 47458
rect 23998 47406 24050 47458
rect 32622 47406 32674 47458
rect 33070 47406 33122 47458
rect 38558 47406 38610 47458
rect 39230 47406 39282 47458
rect 39902 47406 39954 47458
rect 18174 47294 18226 47346
rect 21646 47294 21698 47346
rect 31838 47294 31890 47346
rect 32174 47294 32226 47346
rect 37998 47294 38050 47346
rect 38222 47294 38274 47346
rect 12910 47182 12962 47234
rect 13582 47182 13634 47234
rect 22990 47182 23042 47234
rect 26350 47182 26402 47234
rect 35534 47182 35586 47234
rect 35982 47182 36034 47234
rect 42366 47182 42418 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 10894 46846 10946 46898
rect 11678 46846 11730 46898
rect 12910 46846 12962 46898
rect 25342 46846 25394 46898
rect 31278 46846 31330 46898
rect 39454 46846 39506 46898
rect 40238 46846 40290 46898
rect 9550 46734 9602 46786
rect 17390 46734 17442 46786
rect 26350 46734 26402 46786
rect 27806 46734 27858 46786
rect 31950 46734 32002 46786
rect 32398 46734 32450 46786
rect 35198 46734 35250 46786
rect 35758 46734 35810 46786
rect 38670 46734 38722 46786
rect 9886 46622 9938 46674
rect 11230 46622 11282 46674
rect 13134 46622 13186 46674
rect 13918 46622 13970 46674
rect 17614 46622 17666 46674
rect 26126 46622 26178 46674
rect 27470 46622 27522 46674
rect 30606 46622 30658 46674
rect 38894 46622 38946 46674
rect 16270 46510 16322 46562
rect 30158 46510 30210 46562
rect 34974 46510 35026 46562
rect 25678 46398 25730 46450
rect 31614 46398 31666 46450
rect 34638 46398 34690 46450
rect 37774 46398 37826 46450
rect 38110 46398 38162 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 11678 46062 11730 46114
rect 27358 46062 27410 46114
rect 27694 46062 27746 46114
rect 41134 46062 41186 46114
rect 19630 45950 19682 46002
rect 26910 45950 26962 46002
rect 40014 45950 40066 46002
rect 8318 45838 8370 45890
rect 8878 45838 8930 45890
rect 12014 45838 12066 45890
rect 12686 45838 12738 45890
rect 14030 45838 14082 45890
rect 16270 45838 16322 45890
rect 16718 45838 16770 45890
rect 20526 45838 20578 45890
rect 21198 45838 21250 45890
rect 21870 45838 21922 45890
rect 28366 45838 28418 45890
rect 37102 45838 37154 45890
rect 37662 45838 37714 45890
rect 43038 45838 43090 45890
rect 12798 45726 12850 45778
rect 14366 45726 14418 45778
rect 14814 45726 14866 45778
rect 20750 45726 20802 45778
rect 25006 45726 25058 45778
rect 28478 45726 28530 45778
rect 41358 45726 41410 45778
rect 41694 45726 41746 45778
rect 11230 45614 11282 45666
rect 13694 45614 13746 45666
rect 19182 45614 19234 45666
rect 24334 45614 24386 45666
rect 24670 45614 24722 45666
rect 40798 45614 40850 45666
rect 42814 45614 42866 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 10222 45278 10274 45330
rect 13918 45278 13970 45330
rect 17502 45278 17554 45330
rect 20974 45278 21026 45330
rect 25342 45278 25394 45330
rect 29934 45278 29986 45330
rect 31502 45278 31554 45330
rect 37438 45278 37490 45330
rect 37774 45278 37826 45330
rect 11342 45166 11394 45218
rect 18510 45166 18562 45218
rect 26238 45166 26290 45218
rect 40910 45166 40962 45218
rect 11118 45054 11170 45106
rect 13694 45054 13746 45106
rect 18286 45054 18338 45106
rect 26126 45054 26178 45106
rect 27022 45054 27074 45106
rect 27582 45054 27634 45106
rect 30270 45054 30322 45106
rect 31278 45054 31330 45106
rect 34302 45054 34354 45106
rect 35086 45054 35138 45106
rect 37998 45054 38050 45106
rect 39790 45054 39842 45106
rect 42030 45054 42082 45106
rect 42814 45054 42866 45106
rect 30718 44942 30770 44994
rect 33406 44942 33458 44994
rect 33854 44942 33906 44994
rect 39342 44942 39394 44994
rect 41470 44942 41522 44994
rect 45166 44942 45218 44994
rect 10558 44830 10610 44882
rect 17838 44830 17890 44882
rect 20750 44830 20802 44882
rect 21086 44830 21138 44882
rect 25678 44830 25730 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 21646 44494 21698 44546
rect 42478 44494 42530 44546
rect 10446 44382 10498 44434
rect 10894 44382 10946 44434
rect 11678 44382 11730 44434
rect 18398 44382 18450 44434
rect 30158 44382 30210 44434
rect 41806 44382 41858 44434
rect 7534 44270 7586 44322
rect 8094 44270 8146 44322
rect 21982 44270 22034 44322
rect 22430 44270 22482 44322
rect 23326 44270 23378 44322
rect 24110 44270 24162 44322
rect 30494 44270 30546 44322
rect 31166 44270 31218 44322
rect 34414 44270 34466 44322
rect 34862 44270 34914 44322
rect 35870 44270 35922 44322
rect 42814 44270 42866 44322
rect 20190 44158 20242 44210
rect 22766 44158 22818 44210
rect 27918 44158 27970 44210
rect 34974 44158 35026 44210
rect 43038 44158 43090 44210
rect 43374 44158 43426 44210
rect 12126 44046 12178 44098
rect 17950 44046 18002 44098
rect 19854 44046 19906 44098
rect 26462 44046 26514 44098
rect 27358 44046 27410 44098
rect 27582 44046 27634 44098
rect 33630 44046 33682 44098
rect 34078 44046 34130 44098
rect 35646 44046 35698 44098
rect 40238 44046 40290 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 8094 43710 8146 43762
rect 23102 43710 23154 43762
rect 31166 43710 31218 43762
rect 12238 43598 12290 43650
rect 17950 43598 18002 43650
rect 18734 43598 18786 43650
rect 25230 43598 25282 43650
rect 28254 43598 28306 43650
rect 29262 43598 29314 43650
rect 29822 43598 29874 43650
rect 32286 43598 32338 43650
rect 34302 43598 34354 43650
rect 35198 43598 35250 43650
rect 37998 43598 38050 43650
rect 39342 43598 39394 43650
rect 39902 43598 39954 43650
rect 41470 43598 41522 43650
rect 43150 43598 43202 43650
rect 4734 43486 4786 43538
rect 5294 43486 5346 43538
rect 8430 43486 8482 43538
rect 12014 43486 12066 43538
rect 12686 43486 12738 43538
rect 13134 43486 13186 43538
rect 18174 43486 18226 43538
rect 18958 43486 19010 43538
rect 19630 43486 19682 43538
rect 25454 43486 25506 43538
rect 28030 43486 28082 43538
rect 28702 43486 28754 43538
rect 32062 43486 32114 43538
rect 34078 43486 34130 43538
rect 34862 43486 34914 43538
rect 38334 43486 38386 43538
rect 38782 43486 38834 43538
rect 41358 43486 41410 43538
rect 42814 43486 42866 43538
rect 7646 43374 7698 43426
rect 8878 43374 8930 43426
rect 11566 43374 11618 43426
rect 15598 43374 15650 43426
rect 17614 43374 17666 43426
rect 22094 43374 22146 43426
rect 29038 43262 29090 43314
rect 31502 43262 31554 43314
rect 39118 43262 39170 43314
rect 42030 43262 42082 43314
rect 42366 43262 42418 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 8654 42926 8706 42978
rect 13582 42926 13634 42978
rect 21422 42926 21474 42978
rect 42702 42926 42754 42978
rect 10670 42814 10722 42866
rect 18846 42814 18898 42866
rect 23550 42814 23602 42866
rect 36318 42814 36370 42866
rect 8990 42702 9042 42754
rect 9774 42702 9826 42754
rect 11118 42702 11170 42754
rect 11454 42702 11506 42754
rect 12014 42702 12066 42754
rect 13918 42702 13970 42754
rect 14366 42702 14418 42754
rect 15486 42702 15538 42754
rect 16046 42702 16098 42754
rect 18398 42702 18450 42754
rect 21758 42702 21810 42754
rect 22206 42702 22258 42754
rect 23774 42702 23826 42754
rect 24558 42702 24610 42754
rect 37774 42702 37826 42754
rect 38222 42702 38274 42754
rect 43038 42702 43090 42754
rect 43486 42702 43538 42754
rect 5630 42590 5682 42642
rect 5966 42590 6018 42642
rect 9662 42590 9714 42642
rect 14702 42590 14754 42642
rect 22542 42590 22594 42642
rect 35310 42590 35362 42642
rect 43822 42590 43874 42642
rect 26910 42478 26962 42530
rect 35646 42478 35698 42530
rect 40686 42478 40738 42530
rect 41134 42478 41186 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 6526 42142 6578 42194
rect 18958 42142 19010 42194
rect 25342 42142 25394 42194
rect 45726 42142 45778 42194
rect 7646 42030 7698 42082
rect 9998 42030 10050 42082
rect 26238 42030 26290 42082
rect 31054 42030 31106 42082
rect 39790 42030 39842 42082
rect 7534 41918 7586 41970
rect 9662 41918 9714 41970
rect 19182 41918 19234 41970
rect 19966 41918 20018 41970
rect 26126 41918 26178 41970
rect 27806 41918 27858 41970
rect 28254 41918 28306 41970
rect 31278 41918 31330 41970
rect 32958 41918 33010 41970
rect 33630 41918 33682 41970
rect 38782 41918 38834 41970
rect 39342 41918 39394 41970
rect 40014 41918 40066 41970
rect 41022 41918 41074 41970
rect 42366 41918 42418 41970
rect 42590 41918 42642 41970
rect 43262 41918 43314 41970
rect 22318 41806 22370 41858
rect 30718 41806 30770 41858
rect 31838 41806 31890 41858
rect 36094 41806 36146 41858
rect 36430 41806 36482 41858
rect 6862 41694 6914 41746
rect 25678 41694 25730 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 34974 41358 35026 41410
rect 35310 41358 35362 41410
rect 19182 41246 19234 41298
rect 19630 41246 19682 41298
rect 26686 41246 26738 41298
rect 27694 41246 27746 41298
rect 6638 41134 6690 41186
rect 9326 41134 9378 41186
rect 9998 41134 10050 41186
rect 15038 41134 15090 41186
rect 16270 41134 16322 41186
rect 16830 41134 16882 41186
rect 21758 41134 21810 41186
rect 22206 41134 22258 41186
rect 29598 41134 29650 41186
rect 30158 41134 30210 41186
rect 33406 41134 33458 41186
rect 34078 41134 34130 41186
rect 38446 41134 38498 41186
rect 38894 41134 38946 41186
rect 39454 41134 39506 41186
rect 42590 41134 42642 41186
rect 15262 41022 15314 41074
rect 20190 41022 20242 41074
rect 20526 41022 20578 41074
rect 21422 41022 21474 41074
rect 22430 41022 22482 41074
rect 24446 41022 24498 41074
rect 34190 41022 34242 41074
rect 35534 41022 35586 41074
rect 36094 41022 36146 41074
rect 42814 41022 42866 41074
rect 43150 41022 43202 41074
rect 6414 40910 6466 40962
rect 12462 40910 12514 40962
rect 12910 40910 12962 40962
rect 14366 40910 14418 40962
rect 14478 40910 14530 40962
rect 14590 40910 14642 40962
rect 15374 40910 15426 40962
rect 23102 40910 23154 40962
rect 24110 40910 24162 40962
rect 27246 40910 27298 40962
rect 32510 40910 32562 40962
rect 33070 40910 33122 40962
rect 41806 40910 41858 40962
rect 42254 40910 42306 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 9662 40574 9714 40626
rect 15262 40574 15314 40626
rect 15486 40574 15538 40626
rect 22990 40574 23042 40626
rect 25342 40574 25394 40626
rect 30718 40574 30770 40626
rect 33406 40574 33458 40626
rect 39118 40574 39170 40626
rect 41694 40574 41746 40626
rect 8990 40462 9042 40514
rect 10558 40462 10610 40514
rect 15710 40462 15762 40514
rect 17614 40462 17666 40514
rect 26462 40462 26514 40514
rect 31614 40462 31666 40514
rect 33070 40462 33122 40514
rect 40014 40462 40066 40514
rect 2382 40350 2434 40402
rect 3166 40350 3218 40402
rect 5518 40350 5570 40402
rect 5854 40350 5906 40402
rect 6526 40350 6578 40402
rect 10670 40350 10722 40402
rect 12126 40350 12178 40402
rect 12798 40350 12850 40402
rect 15822 40350 15874 40402
rect 16270 40350 16322 40402
rect 17502 40350 17554 40402
rect 18286 40350 18338 40402
rect 19182 40350 19234 40402
rect 20190 40350 20242 40402
rect 23550 40350 23602 40402
rect 26350 40350 26402 40402
rect 27358 40350 27410 40402
rect 27918 40350 27970 40402
rect 31726 40350 31778 40402
rect 32510 40350 32562 40402
rect 40126 40350 40178 40402
rect 41918 40350 41970 40402
rect 42590 40350 42642 40402
rect 45054 40350 45106 40402
rect 19742 40238 19794 40290
rect 20974 40238 21026 40290
rect 21758 40238 21810 40290
rect 24222 40238 24274 40290
rect 24670 40238 24722 40290
rect 30270 40238 30322 40290
rect 9998 40126 10050 40178
rect 18622 40126 18674 40178
rect 19182 40126 19234 40178
rect 19742 40126 19794 40178
rect 25678 40126 25730 40178
rect 31054 40126 31106 40178
rect 39454 40126 39506 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 6750 39790 6802 39842
rect 7086 39790 7138 39842
rect 12238 39790 12290 39842
rect 30494 39678 30546 39730
rect 34974 39678 35026 39730
rect 7534 39566 7586 39618
rect 16942 39566 16994 39618
rect 17502 39566 17554 39618
rect 20526 39566 20578 39618
rect 22094 39566 22146 39618
rect 23326 39566 23378 39618
rect 24110 39566 24162 39618
rect 28142 39566 28194 39618
rect 37102 39566 37154 39618
rect 42254 39566 42306 39618
rect 3278 39454 3330 39506
rect 3614 39454 3666 39506
rect 7646 39454 7698 39506
rect 12462 39454 12514 39506
rect 14030 39454 14082 39506
rect 14702 39454 14754 39506
rect 21758 39454 21810 39506
rect 22318 39454 22370 39506
rect 22878 39454 22930 39506
rect 27918 39454 27970 39506
rect 42590 39454 42642 39506
rect 5742 39342 5794 39394
rect 9214 39342 9266 39394
rect 11678 39342 11730 39394
rect 11902 39342 11954 39394
rect 13022 39342 13074 39394
rect 13694 39342 13746 39394
rect 14366 39342 14418 39394
rect 14590 39342 14642 39394
rect 19854 39342 19906 39394
rect 20750 39342 20802 39394
rect 26462 39342 26514 39394
rect 27134 39342 27186 39394
rect 27470 39342 27522 39394
rect 34526 39342 34578 39394
rect 37326 39342 37378 39394
rect 40350 39342 40402 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 8990 39006 9042 39058
rect 11566 39006 11618 39058
rect 11790 39006 11842 39058
rect 17502 39006 17554 39058
rect 23214 39006 23266 39058
rect 28142 39006 28194 39058
rect 11902 38894 11954 38946
rect 17614 38894 17666 38946
rect 18510 38894 18562 38946
rect 18622 38894 18674 38946
rect 19630 38894 19682 38946
rect 28702 38894 28754 38946
rect 29038 38894 29090 38946
rect 30830 38894 30882 38946
rect 31950 38894 32002 38946
rect 32286 38894 32338 38946
rect 34750 38894 34802 38946
rect 35086 38894 35138 38946
rect 39566 38894 39618 38946
rect 41246 38894 41298 38946
rect 1822 38782 1874 38834
rect 2270 38782 2322 38834
rect 5182 38782 5234 38834
rect 5854 38782 5906 38834
rect 6638 38782 6690 38834
rect 9662 38782 9714 38834
rect 10782 38782 10834 38834
rect 12238 38782 12290 38834
rect 12686 38782 12738 38834
rect 13358 38782 13410 38834
rect 17390 38782 17442 38834
rect 18062 38782 18114 38834
rect 18846 38782 18898 38834
rect 19518 38782 19570 38834
rect 20190 38782 20242 38834
rect 20750 38782 20802 38834
rect 24334 38782 24386 38834
rect 26014 38782 26066 38834
rect 27246 38782 27298 38834
rect 30606 38782 30658 38834
rect 31614 38782 31666 38834
rect 34526 38782 34578 38834
rect 38222 38782 38274 38834
rect 39006 38782 39058 38834
rect 39230 38782 39282 38834
rect 41022 38782 41074 38834
rect 4734 38670 4786 38722
rect 11342 38670 11394 38722
rect 12350 38670 12402 38722
rect 15710 38670 15762 38722
rect 16046 38670 16098 38722
rect 16158 38670 16210 38722
rect 19294 38670 19346 38722
rect 23774 38670 23826 38722
rect 24110 38670 24162 38722
rect 25454 38670 25506 38722
rect 25790 38670 25842 38722
rect 26798 38670 26850 38722
rect 27694 38670 27746 38722
rect 31278 38670 31330 38722
rect 35870 38670 35922 38722
rect 40014 38670 40066 38722
rect 24670 38558 24722 38610
rect 26350 38558 26402 38610
rect 28478 38558 28530 38610
rect 34190 38558 34242 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 3838 38222 3890 38274
rect 10558 38222 10610 38274
rect 37102 38222 37154 38274
rect 37438 38222 37490 38274
rect 38782 38222 38834 38274
rect 6078 38110 6130 38162
rect 9662 38110 9714 38162
rect 12238 38110 12290 38162
rect 14142 38110 14194 38162
rect 14814 38110 14866 38162
rect 16718 38110 16770 38162
rect 17614 38110 17666 38162
rect 21646 38110 21698 38162
rect 22430 38110 22482 38162
rect 22990 38110 23042 38162
rect 24110 38110 24162 38162
rect 27806 38110 27858 38162
rect 33854 38110 33906 38162
rect 4174 37998 4226 38050
rect 4846 37998 4898 38050
rect 11454 37998 11506 38050
rect 12350 37998 12402 38050
rect 13694 37998 13746 38050
rect 14366 37998 14418 38050
rect 17166 37998 17218 38050
rect 18958 37998 19010 38050
rect 19182 37998 19234 38050
rect 19742 37998 19794 38050
rect 20078 37998 20130 38050
rect 23214 37998 23266 38050
rect 25342 37998 25394 38050
rect 25678 37998 25730 38050
rect 26686 37998 26738 38050
rect 27470 37998 27522 38050
rect 27694 37998 27746 38050
rect 28142 37998 28194 38050
rect 30942 37998 30994 38050
rect 31390 37998 31442 38050
rect 35422 37998 35474 38050
rect 39118 37998 39170 38050
rect 39790 37998 39842 38050
rect 40574 37998 40626 38050
rect 41246 37998 41298 38050
rect 2270 37886 2322 37938
rect 2606 37886 2658 37938
rect 4958 37886 5010 37938
rect 5742 37886 5794 37938
rect 6302 37886 6354 37938
rect 6862 37886 6914 37938
rect 7422 37886 7474 37938
rect 7758 37886 7810 37938
rect 9438 37886 9490 37938
rect 10334 37886 10386 37938
rect 11230 37886 11282 37938
rect 12462 37886 12514 37938
rect 16270 37886 16322 37938
rect 16606 37886 16658 37938
rect 16942 37886 16994 37938
rect 17502 37886 17554 37938
rect 17726 37886 17778 37938
rect 20414 37886 20466 37938
rect 20526 37886 20578 37938
rect 24558 37886 24610 37938
rect 24670 37886 24722 37938
rect 26574 37886 26626 37938
rect 35870 37886 35922 37938
rect 37662 37886 37714 37938
rect 37998 37886 38050 37938
rect 39902 37886 39954 37938
rect 9998 37774 10050 37826
rect 10894 37774 10946 37826
rect 14702 37774 14754 37826
rect 14926 37774 14978 37826
rect 15486 37774 15538 37826
rect 18734 37774 18786 37826
rect 19406 37774 19458 37826
rect 19518 37774 19570 37826
rect 19854 37774 19906 37826
rect 20750 37774 20802 37826
rect 21982 37774 22034 37826
rect 23550 37774 23602 37826
rect 24334 37774 24386 37826
rect 25902 37774 25954 37826
rect 26014 37774 26066 37826
rect 26126 37774 26178 37826
rect 26350 37774 26402 37826
rect 27918 37774 27970 37826
rect 29710 37774 29762 37826
rect 34302 37774 34354 37826
rect 43710 37774 43762 37826
rect 44158 37774 44210 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 5182 37438 5234 37490
rect 10222 37438 10274 37490
rect 15486 37438 15538 37490
rect 16382 37438 16434 37490
rect 24334 37438 24386 37490
rect 24558 37438 24610 37490
rect 25566 37438 25618 37490
rect 25790 37438 25842 37490
rect 26462 37438 26514 37490
rect 41134 37438 41186 37490
rect 10110 37326 10162 37378
rect 10894 37326 10946 37378
rect 11006 37326 11058 37378
rect 12014 37326 12066 37378
rect 13918 37326 13970 37378
rect 15038 37326 15090 37378
rect 18286 37326 18338 37378
rect 29486 37326 29538 37378
rect 42254 37326 42306 37378
rect 43150 37326 43202 37378
rect 1822 37214 1874 37266
rect 2382 37214 2434 37266
rect 9102 37214 9154 37266
rect 10446 37214 10498 37266
rect 10670 37214 10722 37266
rect 11342 37214 11394 37266
rect 11790 37214 11842 37266
rect 12462 37214 12514 37266
rect 13246 37214 13298 37266
rect 13470 37214 13522 37266
rect 14142 37214 14194 37266
rect 15598 37214 15650 37266
rect 16046 37214 16098 37266
rect 16382 37214 16434 37266
rect 16718 37214 16770 37266
rect 20078 37214 20130 37266
rect 22206 37214 22258 37266
rect 22766 37214 22818 37266
rect 23102 37214 23154 37266
rect 23886 37214 23938 37266
rect 24110 37214 24162 37266
rect 25342 37214 25394 37266
rect 26014 37214 26066 37266
rect 27022 37214 27074 37266
rect 28926 37214 28978 37266
rect 29262 37214 29314 37266
rect 30046 37214 30098 37266
rect 33070 37214 33122 37266
rect 39678 37214 39730 37266
rect 40462 37214 40514 37266
rect 41470 37214 41522 37266
rect 41918 37214 41970 37266
rect 42926 37214 42978 37266
rect 43374 37214 43426 37266
rect 44046 37214 44098 37266
rect 4734 37102 4786 37154
rect 9886 37102 9938 37154
rect 11454 37102 11506 37154
rect 13694 37102 13746 37154
rect 14702 37102 14754 37154
rect 20638 37102 20690 37154
rect 21310 37102 21362 37154
rect 22318 37102 22370 37154
rect 23774 37102 23826 37154
rect 26126 37102 26178 37154
rect 28254 37102 28306 37154
rect 28702 37102 28754 37154
rect 29822 37102 29874 37154
rect 30830 37102 30882 37154
rect 31726 37102 31778 37154
rect 32062 37102 32114 37154
rect 32510 37102 32562 37154
rect 34526 37102 34578 37154
rect 37326 37102 37378 37154
rect 46510 37102 46562 37154
rect 13358 36990 13410 37042
rect 15710 36990 15762 37042
rect 22094 36990 22146 37042
rect 29150 36990 29202 37042
rect 30382 36990 30434 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 8206 36654 8258 36706
rect 19854 36654 19906 36706
rect 24894 36654 24946 36706
rect 32398 36654 32450 36706
rect 43038 36654 43090 36706
rect 43374 36654 43426 36706
rect 11230 36542 11282 36594
rect 33182 36542 33234 36594
rect 37438 36542 37490 36594
rect 6078 36430 6130 36482
rect 8542 36430 8594 36482
rect 10670 36430 10722 36482
rect 12350 36430 12402 36482
rect 12574 36430 12626 36482
rect 12798 36430 12850 36482
rect 12910 36430 12962 36482
rect 14030 36430 14082 36482
rect 15150 36430 15202 36482
rect 15598 36430 15650 36482
rect 16158 36430 16210 36482
rect 19406 36430 19458 36482
rect 19966 36430 20018 36482
rect 21534 36430 21586 36482
rect 22094 36430 22146 36482
rect 22542 36430 22594 36482
rect 23326 36430 23378 36482
rect 23550 36430 23602 36482
rect 25118 36430 25170 36482
rect 26014 36430 26066 36482
rect 26238 36430 26290 36482
rect 27582 36430 27634 36482
rect 27806 36430 27858 36482
rect 28142 36430 28194 36482
rect 29710 36430 29762 36482
rect 30382 36430 30434 36482
rect 33518 36430 33570 36482
rect 34414 36430 34466 36482
rect 35310 36430 35362 36482
rect 2494 36318 2546 36370
rect 2830 36318 2882 36370
rect 5742 36318 5794 36370
rect 6302 36318 6354 36370
rect 6862 36318 6914 36370
rect 8766 36318 8818 36370
rect 9102 36318 9154 36370
rect 11566 36318 11618 36370
rect 11902 36318 11954 36370
rect 14254 36318 14306 36370
rect 18510 36318 18562 36370
rect 18958 36318 19010 36370
rect 19630 36318 19682 36370
rect 21422 36318 21474 36370
rect 23102 36318 23154 36370
rect 23774 36318 23826 36370
rect 24782 36318 24834 36370
rect 26574 36318 26626 36370
rect 27918 36318 27970 36370
rect 29374 36318 29426 36370
rect 29934 36318 29986 36370
rect 30046 36318 30098 36370
rect 32174 36318 32226 36370
rect 33742 36318 33794 36370
rect 34078 36318 34130 36370
rect 43710 36318 43762 36370
rect 44158 36318 44210 36370
rect 10110 36206 10162 36258
rect 10558 36206 10610 36258
rect 11006 36206 11058 36258
rect 11230 36206 11282 36258
rect 13694 36206 13746 36258
rect 15038 36206 15090 36258
rect 18846 36206 18898 36258
rect 19518 36206 19570 36258
rect 20862 36206 20914 36258
rect 22654 36206 22706 36258
rect 23886 36206 23938 36258
rect 24222 36206 24274 36258
rect 24558 36206 24610 36258
rect 25454 36206 25506 36258
rect 26350 36206 26402 36258
rect 27022 36206 27074 36258
rect 28590 36206 28642 36258
rect 29822 36206 29874 36258
rect 31166 36206 31218 36258
rect 31614 36206 31666 36258
rect 32734 36206 32786 36258
rect 35086 36206 35138 36258
rect 40574 36206 40626 36258
rect 44942 36206 44994 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 8542 35870 8594 35922
rect 10782 35870 10834 35922
rect 14254 35870 14306 35922
rect 14590 35870 14642 35922
rect 15374 35870 15426 35922
rect 15822 35870 15874 35922
rect 16158 35870 16210 35922
rect 16270 35870 16322 35922
rect 16382 35870 16434 35922
rect 21646 35870 21698 35922
rect 23102 35870 23154 35922
rect 28142 35870 28194 35922
rect 29486 35870 29538 35922
rect 30942 35870 30994 35922
rect 32286 35870 32338 35922
rect 43262 35870 43314 35922
rect 9662 35758 9714 35810
rect 10222 35758 10274 35810
rect 16606 35758 16658 35810
rect 22206 35758 22258 35810
rect 22542 35758 22594 35810
rect 22990 35758 23042 35810
rect 24110 35758 24162 35810
rect 26462 35758 26514 35810
rect 27806 35758 27858 35810
rect 28366 35758 28418 35810
rect 29038 35758 29090 35810
rect 29934 35758 29986 35810
rect 31950 35758 32002 35810
rect 32510 35758 32562 35810
rect 33854 35758 33906 35810
rect 42702 35758 42754 35810
rect 5630 35646 5682 35698
rect 6190 35646 6242 35698
rect 13918 35646 13970 35698
rect 18734 35646 18786 35698
rect 21982 35646 22034 35698
rect 22766 35646 22818 35698
rect 23662 35646 23714 35698
rect 28142 35646 28194 35698
rect 29262 35646 29314 35698
rect 29598 35646 29650 35698
rect 30158 35646 30210 35698
rect 30494 35646 30546 35698
rect 32286 35646 32338 35698
rect 33630 35646 33682 35698
rect 34526 35646 34578 35698
rect 35086 35646 35138 35698
rect 39790 35646 39842 35698
rect 41918 35646 41970 35698
rect 42366 35646 42418 35698
rect 10446 35534 10498 35586
rect 12686 35534 12738 35586
rect 18174 35534 18226 35586
rect 20190 35534 20242 35586
rect 23550 35534 23602 35586
rect 25678 35534 25730 35586
rect 26126 35534 26178 35586
rect 26686 35534 26738 35586
rect 27470 35534 27522 35586
rect 30046 35534 30098 35586
rect 31390 35534 31442 35586
rect 37438 35534 37490 35586
rect 39230 35534 39282 35586
rect 41246 35534 41298 35586
rect 23326 35422 23378 35474
rect 27022 35422 27074 35474
rect 30830 35422 30882 35474
rect 31614 35422 31666 35474
rect 33294 35422 33346 35474
rect 41582 35422 41634 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 18846 35086 18898 35138
rect 20190 35086 20242 35138
rect 35198 35086 35250 35138
rect 10334 34974 10386 35026
rect 10558 34974 10610 35026
rect 11118 34974 11170 35026
rect 12238 34974 12290 35026
rect 14254 34974 14306 35026
rect 21646 34974 21698 35026
rect 26238 34974 26290 35026
rect 32622 34974 32674 35026
rect 34526 34974 34578 35026
rect 42142 34974 42194 35026
rect 1822 34862 1874 34914
rect 2382 34862 2434 34914
rect 4734 34862 4786 34914
rect 8318 34862 8370 34914
rect 10782 34862 10834 34914
rect 13806 34862 13858 34914
rect 16606 34862 16658 34914
rect 16942 34862 16994 34914
rect 18062 34862 18114 34914
rect 18286 34862 18338 34914
rect 18622 34862 18674 34914
rect 18958 34862 19010 34914
rect 19742 34862 19794 34914
rect 20078 34862 20130 34914
rect 20526 34862 20578 34914
rect 22878 34862 22930 34914
rect 25006 34862 25058 34914
rect 25118 34862 25170 34914
rect 26686 34862 26738 34914
rect 27022 34862 27074 34914
rect 6414 34750 6466 34802
rect 6750 34750 6802 34802
rect 7982 34750 8034 34802
rect 8542 34750 8594 34802
rect 8878 34750 8930 34802
rect 11678 34750 11730 34802
rect 11790 34750 11842 34802
rect 12014 34750 12066 34802
rect 12574 34750 12626 34802
rect 12910 34750 12962 34802
rect 14590 34750 14642 34802
rect 22318 34750 22370 34802
rect 25454 34750 25506 34802
rect 27246 34806 27298 34858
rect 27470 34862 27522 34914
rect 28030 34862 28082 34914
rect 28142 34862 28194 34914
rect 28254 34862 28306 34914
rect 28590 34862 28642 34914
rect 29710 34862 29762 34914
rect 30494 34862 30546 34914
rect 31054 34862 31106 34914
rect 31502 34862 31554 34914
rect 35534 34862 35586 34914
rect 36206 34862 36258 34914
rect 37662 34862 37714 34914
rect 38222 34862 38274 34914
rect 40574 34862 40626 34914
rect 41246 34862 41298 34914
rect 27358 34750 27410 34802
rect 29822 34750 29874 34802
rect 36094 34750 36146 34802
rect 37102 34750 37154 34802
rect 43038 34750 43090 34802
rect 43374 34750 43426 34802
rect 46510 34750 46562 34802
rect 9662 34638 9714 34690
rect 11454 34638 11506 34690
rect 13470 34638 13522 34690
rect 14926 34638 14978 34690
rect 15374 34638 15426 34690
rect 16830 34638 16882 34690
rect 19070 34638 19122 34690
rect 20526 34638 20578 34690
rect 21982 34638 22034 34690
rect 23214 34638 23266 34690
rect 24558 34638 24610 34690
rect 25342 34638 25394 34690
rect 25790 34638 25842 34690
rect 27806 34638 27858 34690
rect 29262 34638 29314 34690
rect 31054 34638 31106 34690
rect 37886 34638 37938 34690
rect 41582 34638 41634 34690
rect 42478 34638 42530 34690
rect 43710 34638 43762 34690
rect 44158 34638 44210 34690
rect 46174 34638 46226 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 2382 34302 2434 34354
rect 10446 34302 10498 34354
rect 17390 34302 17442 34354
rect 18062 34302 18114 34354
rect 19518 34302 19570 34354
rect 20638 34302 20690 34354
rect 21086 34302 21138 34354
rect 31614 34302 31666 34354
rect 33854 34302 33906 34354
rect 34190 34302 34242 34354
rect 35086 34302 35138 34354
rect 37998 34302 38050 34354
rect 39678 34302 39730 34354
rect 41022 34302 41074 34354
rect 46622 34302 46674 34354
rect 5070 34190 5122 34242
rect 5742 34190 5794 34242
rect 17726 34190 17778 34242
rect 25566 34190 25618 34242
rect 26238 34190 26290 34242
rect 27582 34190 27634 34242
rect 28590 34190 28642 34242
rect 30942 34190 30994 34242
rect 31950 34190 32002 34242
rect 33294 34190 33346 34242
rect 33630 34190 33682 34242
rect 34526 34190 34578 34242
rect 35870 34190 35922 34242
rect 36206 34190 36258 34242
rect 38670 34190 38722 34242
rect 38894 34190 38946 34242
rect 42142 34190 42194 34242
rect 42702 34190 42754 34242
rect 46174 34190 46226 34242
rect 47182 34190 47234 34242
rect 47518 34190 47570 34242
rect 2718 34078 2770 34130
rect 4174 34078 4226 34130
rect 4510 34078 4562 34130
rect 5294 34078 5346 34130
rect 6190 34078 6242 34130
rect 13358 34078 13410 34130
rect 13918 34078 13970 34130
rect 14478 34078 14530 34130
rect 16830 34078 16882 34130
rect 18398 34078 18450 34130
rect 18734 34078 18786 34130
rect 18958 34078 19010 34130
rect 19182 34078 19234 34130
rect 19406 34078 19458 34130
rect 21310 34078 21362 34130
rect 21982 34078 22034 34130
rect 25454 34078 25506 34130
rect 26686 34078 26738 34130
rect 27470 34078 27522 34130
rect 28030 34078 28082 34130
rect 28926 34078 28978 34130
rect 29038 34078 29090 34130
rect 29262 34078 29314 34130
rect 29822 34078 29874 34130
rect 31054 34078 31106 34130
rect 32286 34078 32338 34130
rect 32510 34078 32562 34130
rect 33406 34078 33458 34130
rect 38334 34078 38386 34130
rect 43262 34078 43314 34130
rect 43710 34078 43762 34130
rect 46958 34078 47010 34130
rect 6750 33966 6802 34018
rect 9886 33966 9938 34018
rect 11118 33966 11170 34018
rect 19966 33966 20018 34018
rect 24446 33966 24498 34018
rect 26238 33966 26290 34018
rect 27806 33966 27858 34018
rect 30270 33966 30322 34018
rect 30382 33966 30434 34018
rect 32062 33966 32114 34018
rect 33518 33966 33570 34018
rect 36430 33854 36482 33906
rect 36766 33854 36818 33906
rect 41582 33854 41634 33906
rect 41918 33854 41970 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 3838 33518 3890 33570
rect 16382 33518 16434 33570
rect 17166 33518 17218 33570
rect 18062 33518 18114 33570
rect 18286 33518 18338 33570
rect 18734 33518 18786 33570
rect 22542 33518 22594 33570
rect 24558 33518 24610 33570
rect 25006 33518 25058 33570
rect 34750 33518 34802 33570
rect 43038 33518 43090 33570
rect 8990 33406 9042 33458
rect 15598 33406 15650 33458
rect 17166 33406 17218 33458
rect 17726 33406 17778 33458
rect 19406 33406 19458 33458
rect 24334 33406 24386 33458
rect 29374 33406 29426 33458
rect 33966 33406 34018 33458
rect 38558 33406 38610 33458
rect 41246 33406 41298 33458
rect 4398 33294 4450 33346
rect 6078 33294 6130 33346
rect 6638 33294 6690 33346
rect 10334 33294 10386 33346
rect 15822 33294 15874 33346
rect 16718 33294 16770 33346
rect 19518 33294 19570 33346
rect 19966 33294 20018 33346
rect 22878 33294 22930 33346
rect 24110 33294 24162 33346
rect 25342 33294 25394 33346
rect 28702 33294 28754 33346
rect 29934 33294 29986 33346
rect 30942 33294 30994 33346
rect 32734 33294 32786 33346
rect 33294 33294 33346 33346
rect 35086 33294 35138 33346
rect 36990 33294 37042 33346
rect 38222 33294 38274 33346
rect 39566 33294 39618 33346
rect 42142 33294 42194 33346
rect 42590 33294 42642 33346
rect 43374 33294 43426 33346
rect 43822 33294 43874 33346
rect 45278 33294 45330 33346
rect 45950 33294 46002 33346
rect 4622 33182 4674 33234
rect 10222 33182 10274 33234
rect 10670 33182 10722 33234
rect 12126 33182 12178 33234
rect 13806 33182 13858 33234
rect 15486 33182 15538 33234
rect 16046 33182 16098 33234
rect 16494 33182 16546 33234
rect 23214 33182 23266 33234
rect 23662 33182 23714 33234
rect 27134 33182 27186 33234
rect 28366 33182 28418 33234
rect 28478 33182 28530 33234
rect 29710 33182 29762 33234
rect 30718 33182 30770 33234
rect 32846 33182 32898 33234
rect 35310 33182 35362 33234
rect 35870 33182 35922 33234
rect 41918 33182 41970 33234
rect 43934 33182 43986 33234
rect 3502 33070 3554 33122
rect 10894 33070 10946 33122
rect 11006 33070 11058 33122
rect 11790 33070 11842 33122
rect 12462 33070 12514 33122
rect 12910 33070 12962 33122
rect 13470 33070 13522 33122
rect 14366 33070 14418 33122
rect 18174 33070 18226 33122
rect 18622 33070 18674 33122
rect 19294 33070 19346 33122
rect 20414 33070 20466 33122
rect 20862 33070 20914 33122
rect 26798 33070 26850 33122
rect 27582 33070 27634 33122
rect 28142 33070 28194 33122
rect 31502 33070 31554 33122
rect 32398 33070 32450 33122
rect 32958 33070 33010 33122
rect 37326 33070 37378 33122
rect 37774 33070 37826 33122
rect 42254 33070 42306 33122
rect 48302 33070 48354 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4734 32734 4786 32786
rect 6974 32734 7026 32786
rect 9662 32734 9714 32786
rect 11006 32734 11058 32786
rect 11230 32734 11282 32786
rect 12126 32734 12178 32786
rect 12574 32734 12626 32786
rect 14254 32734 14306 32786
rect 15150 32734 15202 32786
rect 29150 32734 29202 32786
rect 30606 32734 30658 32786
rect 35422 32734 35474 32786
rect 39342 32734 39394 32786
rect 43038 32734 43090 32786
rect 8654 32622 8706 32674
rect 9998 32622 10050 32674
rect 10110 32622 10162 32674
rect 12910 32622 12962 32674
rect 13806 32622 13858 32674
rect 15486 32622 15538 32674
rect 20526 32622 20578 32674
rect 29934 32622 29986 32674
rect 31614 32622 31666 32674
rect 31950 32622 32002 32674
rect 33406 32622 33458 32674
rect 33742 32622 33794 32674
rect 46286 32622 46338 32674
rect 1822 32510 1874 32562
rect 2270 32510 2322 32562
rect 5742 32510 5794 32562
rect 7310 32510 7362 32562
rect 7758 32510 7810 32562
rect 8094 32510 8146 32562
rect 8766 32510 8818 32562
rect 10334 32510 10386 32562
rect 10782 32510 10834 32562
rect 11454 32510 11506 32562
rect 11566 32510 11618 32562
rect 12238 32510 12290 32562
rect 12574 32510 12626 32562
rect 13134 32510 13186 32562
rect 13470 32510 13522 32562
rect 17950 32510 18002 32562
rect 20862 32510 20914 32562
rect 26238 32510 26290 32562
rect 26798 32510 26850 32562
rect 30158 32510 30210 32562
rect 30942 32510 30994 32562
rect 33518 32510 33570 32562
rect 33966 32510 34018 32562
rect 37774 32510 37826 32562
rect 38558 32510 38610 32562
rect 39790 32510 39842 32562
rect 40910 32510 40962 32562
rect 41246 32510 41298 32562
rect 42142 32510 42194 32562
rect 46622 32510 46674 32562
rect 5182 32398 5234 32450
rect 6190 32398 6242 32450
rect 13358 32398 13410 32450
rect 17390 32398 17442 32450
rect 18398 32398 18450 32450
rect 18846 32398 18898 32450
rect 19742 32398 19794 32450
rect 20302 32398 20354 32450
rect 21310 32398 21362 32450
rect 29598 32398 29650 32450
rect 32510 32398 32562 32450
rect 33630 32398 33682 32450
rect 39566 32398 39618 32450
rect 40126 32398 40178 32450
rect 41134 32398 41186 32450
rect 42478 32398 42530 32450
rect 5966 32286 6018 32338
rect 6190 32286 6242 32338
rect 18174 32286 18226 32338
rect 18398 32286 18450 32338
rect 19518 32286 19570 32338
rect 19742 32286 19794 32338
rect 20078 32286 20130 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 3950 31950 4002 32002
rect 21534 31950 21586 32002
rect 33518 31950 33570 32002
rect 11678 31838 11730 31890
rect 18510 31838 18562 31890
rect 18846 31838 18898 31890
rect 23662 31838 23714 31890
rect 32062 31838 32114 31890
rect 40126 31838 40178 31890
rect 43038 31838 43090 31890
rect 2494 31726 2546 31778
rect 4734 31726 4786 31778
rect 15262 31726 15314 31778
rect 15822 31726 15874 31778
rect 19630 31726 19682 31778
rect 19966 31726 20018 31778
rect 21870 31726 21922 31778
rect 22542 31726 22594 31778
rect 26014 31726 26066 31778
rect 27022 31726 27074 31778
rect 27470 31726 27522 31778
rect 30270 31726 30322 31778
rect 31166 31726 31218 31778
rect 32622 31726 32674 31778
rect 32958 31726 33010 31778
rect 33854 31726 33906 31778
rect 34078 31726 34130 31778
rect 37214 31726 37266 31778
rect 40574 31726 40626 31778
rect 41022 31726 41074 31778
rect 42254 31726 42306 31778
rect 45278 31726 45330 31778
rect 45950 31726 46002 31778
rect 2158 31614 2210 31666
rect 4510 31614 4562 31666
rect 11566 31614 11618 31666
rect 11902 31614 11954 31666
rect 12126 31614 12178 31666
rect 18734 31614 18786 31666
rect 20414 31614 20466 31666
rect 20638 31614 20690 31666
rect 22654 31614 22706 31666
rect 23886 31614 23938 31666
rect 24222 31614 24274 31666
rect 26126 31614 26178 31666
rect 26686 31614 26738 31666
rect 29934 31614 29986 31666
rect 33182 31614 33234 31666
rect 40462 31614 40514 31666
rect 40910 31614 40962 31666
rect 43262 31614 43314 31666
rect 43598 31614 43650 31666
rect 3614 31502 3666 31554
rect 12686 31502 12738 31554
rect 18174 31502 18226 31554
rect 19406 31502 19458 31554
rect 19518 31502 19570 31554
rect 20526 31502 20578 31554
rect 23326 31502 23378 31554
rect 25118 31502 25170 31554
rect 25454 31502 25506 31554
rect 27918 31502 27970 31554
rect 30606 31502 30658 31554
rect 31502 31502 31554 31554
rect 32846 31502 32898 31554
rect 34526 31502 34578 31554
rect 35982 31502 36034 31554
rect 37438 31502 37490 31554
rect 39902 31502 39954 31554
rect 42702 31502 42754 31554
rect 43934 31502 43986 31554
rect 48302 31502 48354 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 5406 31166 5458 31218
rect 8878 31166 8930 31218
rect 17502 31166 17554 31218
rect 19070 31166 19122 31218
rect 22766 31166 22818 31218
rect 24670 31166 24722 31218
rect 26126 31166 26178 31218
rect 27134 31166 27186 31218
rect 30046 31166 30098 31218
rect 30830 31166 30882 31218
rect 31726 31166 31778 31218
rect 35646 31166 35698 31218
rect 41022 31166 41074 31218
rect 41134 31166 41186 31218
rect 46622 31166 46674 31218
rect 48302 31166 48354 31218
rect 2158 31054 2210 31106
rect 2494 31054 2546 31106
rect 4398 31054 4450 31106
rect 4846 31054 4898 31106
rect 14590 31054 14642 31106
rect 17390 31054 17442 31106
rect 17726 31054 17778 31106
rect 17950 31054 18002 31106
rect 23886 31054 23938 31106
rect 26462 31054 26514 31106
rect 28254 31054 28306 31106
rect 35086 31054 35138 31106
rect 40910 31054 40962 31106
rect 41470 31054 41522 31106
rect 47182 31054 47234 31106
rect 47518 31054 47570 31106
rect 5070 30942 5122 30994
rect 5966 30942 6018 30994
rect 6526 30942 6578 30994
rect 9662 30942 9714 30994
rect 10222 30942 10274 30994
rect 14814 30942 14866 30994
rect 18622 30942 18674 30994
rect 18958 30942 19010 30994
rect 19406 30942 19458 30994
rect 19742 30942 19794 30994
rect 20302 30942 20354 30994
rect 24110 30942 24162 30994
rect 24446 30942 24498 30994
rect 25230 30942 25282 30994
rect 25454 30942 25506 30994
rect 28030 30942 28082 30994
rect 30270 30942 30322 30994
rect 38670 30942 38722 30994
rect 39454 30942 39506 30994
rect 41358 30942 41410 30994
rect 44718 30942 44770 30994
rect 45278 30942 45330 30994
rect 46958 30942 47010 30994
rect 12574 30830 12626 30882
rect 15374 30830 15426 30882
rect 23550 30830 23602 30882
rect 31278 30830 31330 30882
rect 32174 30830 32226 30882
rect 33182 30830 33234 30882
rect 36318 30830 36370 30882
rect 40350 30830 40402 30882
rect 42366 30830 42418 30882
rect 13694 30718 13746 30770
rect 14030 30718 14082 30770
rect 19182 30718 19234 30770
rect 24334 30718 24386 30770
rect 25678 30718 25730 30770
rect 27470 30718 27522 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 12014 30382 12066 30434
rect 20078 30382 20130 30434
rect 22094 30382 22146 30434
rect 22654 30382 22706 30434
rect 37774 30382 37826 30434
rect 8430 30270 8482 30322
rect 19630 30270 19682 30322
rect 26574 30270 26626 30322
rect 29934 30270 29986 30322
rect 35086 30270 35138 30322
rect 40798 30270 40850 30322
rect 43374 30270 43426 30322
rect 47182 30270 47234 30322
rect 1822 30158 1874 30210
rect 2270 30158 2322 30210
rect 5742 30158 5794 30210
rect 10670 30158 10722 30210
rect 11678 30158 11730 30210
rect 19854 30158 19906 30210
rect 20078 30158 20130 30210
rect 23102 30158 23154 30210
rect 26686 30158 26738 30210
rect 27022 30158 27074 30210
rect 30382 30158 30434 30210
rect 32286 30158 32338 30210
rect 35534 30158 35586 30210
rect 38110 30158 38162 30210
rect 40686 30158 40738 30210
rect 40910 30158 40962 30210
rect 43038 30158 43090 30210
rect 44158 30158 44210 30210
rect 46062 30158 46114 30210
rect 6862 30046 6914 30098
rect 7198 30046 7250 30098
rect 8094 30046 8146 30098
rect 8766 30046 8818 30098
rect 8990 30046 9042 30098
rect 10334 30046 10386 30098
rect 12238 30046 12290 30098
rect 12574 30046 12626 30098
rect 16046 30046 16098 30098
rect 17726 30046 17778 30098
rect 19518 30046 19570 30098
rect 22878 30046 22930 30098
rect 32958 30046 33010 30098
rect 38446 30046 38498 30098
rect 38670 30046 38722 30098
rect 41246 30046 41298 30098
rect 41582 30046 41634 30098
rect 41918 30046 41970 30098
rect 43934 30046 43986 30098
rect 4734 29934 4786 29986
rect 16382 29934 16434 29986
rect 18062 29934 18114 29986
rect 18510 29934 18562 29986
rect 20862 29934 20914 29986
rect 22430 29934 22482 29986
rect 23662 29934 23714 29986
rect 24894 29934 24946 29986
rect 26238 29934 26290 29986
rect 30942 29934 30994 29986
rect 39454 29934 39506 29986
rect 45614 29934 45666 29986
rect 45838 29934 45890 29986
rect 46734 29934 46786 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 23214 29598 23266 29650
rect 24334 29598 24386 29650
rect 28142 29598 28194 29650
rect 30270 29598 30322 29650
rect 36766 29598 36818 29650
rect 44942 29598 44994 29650
rect 13918 29486 13970 29538
rect 14478 29486 14530 29538
rect 18622 29486 18674 29538
rect 19182 29486 19234 29538
rect 22542 29486 22594 29538
rect 29374 29486 29426 29538
rect 31838 29486 31890 29538
rect 33182 29486 33234 29538
rect 34526 29486 34578 29538
rect 39566 29486 39618 29538
rect 41246 29486 41298 29538
rect 15710 29374 15762 29426
rect 18174 29374 18226 29426
rect 21758 29374 21810 29426
rect 22878 29374 22930 29426
rect 23438 29374 23490 29426
rect 23886 29374 23938 29426
rect 24334 29374 24386 29426
rect 24670 29374 24722 29426
rect 25230 29374 25282 29426
rect 26014 29374 26066 29426
rect 28366 29374 28418 29426
rect 28814 29374 28866 29426
rect 30606 29374 30658 29426
rect 31390 29374 31442 29426
rect 34302 29374 34354 29426
rect 34974 29374 35026 29426
rect 35982 29374 36034 29426
rect 37102 29374 37154 29426
rect 38670 29374 38722 29426
rect 39790 29374 39842 29426
rect 41806 29374 41858 29426
rect 42590 29374 42642 29426
rect 45278 29374 45330 29426
rect 45838 29374 45890 29426
rect 48302 29374 48354 29426
rect 16158 29262 16210 29314
rect 17838 29262 17890 29314
rect 22094 29262 22146 29314
rect 32510 29262 32562 29314
rect 33070 29262 33122 29314
rect 33406 29262 33458 29314
rect 33966 29262 34018 29314
rect 35534 29262 35586 29314
rect 36430 29262 36482 29314
rect 38334 29262 38386 29314
rect 39230 29262 39282 29314
rect 13358 29150 13410 29202
rect 13694 29150 13746 29202
rect 24222 29150 24274 29202
rect 25230 29150 25282 29202
rect 25566 29150 25618 29202
rect 40126 29150 40178 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 16606 28814 16658 28866
rect 45950 28814 46002 28866
rect 9886 28702 9938 28754
rect 14254 28702 14306 28754
rect 17390 28702 17442 28754
rect 20414 28702 20466 28754
rect 27470 28702 27522 28754
rect 30718 28702 30770 28754
rect 34190 28702 34242 28754
rect 36094 28702 36146 28754
rect 37438 28702 37490 28754
rect 1822 28590 1874 28642
rect 2494 28590 2546 28642
rect 4846 28590 4898 28642
rect 8206 28590 8258 28642
rect 8318 28590 8370 28642
rect 8766 28590 8818 28642
rect 9774 28590 9826 28642
rect 11006 28590 11058 28642
rect 11902 28590 11954 28642
rect 13582 28590 13634 28642
rect 13806 28590 13858 28642
rect 14030 28590 14082 28642
rect 14926 28590 14978 28642
rect 16942 28590 16994 28642
rect 18398 28590 18450 28642
rect 19518 28590 19570 28642
rect 19742 28590 19794 28642
rect 20078 28590 20130 28642
rect 22430 28590 22482 28642
rect 23550 28590 23602 28642
rect 23662 28590 23714 28642
rect 24334 28590 24386 28642
rect 25006 28590 25058 28642
rect 29486 28590 29538 28642
rect 30158 28590 30210 28642
rect 32622 28590 32674 28642
rect 34862 28590 34914 28642
rect 38558 28590 38610 28642
rect 38894 28590 38946 28642
rect 39118 28590 39170 28642
rect 39902 28590 39954 28642
rect 40238 28590 40290 28642
rect 40910 28590 40962 28642
rect 41694 28590 41746 28642
rect 45502 28590 45554 28642
rect 46286 28590 46338 28642
rect 47070 28590 47122 28642
rect 47518 28590 47570 28642
rect 47966 28590 48018 28642
rect 10670 28478 10722 28530
rect 14478 28478 14530 28530
rect 18174 28478 18226 28530
rect 20526 28478 20578 28530
rect 20750 28478 20802 28530
rect 22654 28478 22706 28530
rect 23886 28478 23938 28530
rect 24110 28478 24162 28530
rect 29822 28478 29874 28530
rect 31614 28478 31666 28530
rect 34526 28478 34578 28530
rect 39230 28478 39282 28530
rect 41918 28478 41970 28530
rect 42702 28478 42754 28530
rect 43038 28478 43090 28530
rect 46846 28478 46898 28530
rect 8094 28366 8146 28418
rect 10446 28366 10498 28418
rect 10782 28366 10834 28418
rect 11566 28366 11618 28418
rect 14590 28366 14642 28418
rect 16718 28366 16770 28418
rect 19630 28366 19682 28418
rect 31726 28366 31778 28418
rect 35422 28366 35474 28418
rect 35982 28366 36034 28418
rect 37998 28366 38050 28418
rect 41022 28366 41074 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 2494 28030 2546 28082
rect 8990 28030 9042 28082
rect 9662 28030 9714 28082
rect 13806 28030 13858 28082
rect 16494 28030 16546 28082
rect 18622 28030 18674 28082
rect 21982 28030 22034 28082
rect 22430 28030 22482 28082
rect 24110 28030 24162 28082
rect 25342 28030 25394 28082
rect 25454 28030 25506 28082
rect 29934 28030 29986 28082
rect 30270 28030 30322 28082
rect 31950 28030 32002 28082
rect 42478 28030 42530 28082
rect 45502 28030 45554 28082
rect 47182 28030 47234 28082
rect 5182 27918 5234 27970
rect 9774 27918 9826 27970
rect 10110 27918 10162 27970
rect 14142 27918 14194 27970
rect 14478 27918 14530 27970
rect 14814 27918 14866 27970
rect 16830 27918 16882 27970
rect 26014 27918 26066 27970
rect 30606 27918 30658 27970
rect 33518 27918 33570 27970
rect 44494 27918 44546 27970
rect 46062 27918 46114 27970
rect 46398 27918 46450 27970
rect 2830 27806 2882 27858
rect 4062 27806 4114 27858
rect 4398 27806 4450 27858
rect 4846 27806 4898 27858
rect 6078 27806 6130 27858
rect 6638 27806 6690 27858
rect 9438 27806 9490 27858
rect 10334 27806 10386 27858
rect 10894 27806 10946 27858
rect 11454 27806 11506 27858
rect 15038 27806 15090 27858
rect 17390 27806 17442 27858
rect 17726 27806 17778 27858
rect 18174 27806 18226 27858
rect 19070 27806 19122 27858
rect 19630 27806 19682 27858
rect 26350 27806 26402 27858
rect 26574 27806 26626 27858
rect 27022 27806 27074 27858
rect 27470 27806 27522 27858
rect 31390 27806 31442 27858
rect 33630 27806 33682 27858
rect 34638 27806 34690 27858
rect 35198 27806 35250 27858
rect 35646 27806 35698 27858
rect 38894 27806 38946 27858
rect 41134 27806 41186 27858
rect 42366 27806 42418 27858
rect 42702 27806 42754 27858
rect 44718 27806 44770 27858
rect 17502 27694 17554 27746
rect 17838 27694 17890 27746
rect 26126 27694 26178 27746
rect 30942 27694 30994 27746
rect 33182 27694 33234 27746
rect 34190 27694 34242 27746
rect 36094 27694 36146 27746
rect 38222 27694 38274 27746
rect 39566 27694 39618 27746
rect 40350 27694 40402 27746
rect 48302 27694 48354 27746
rect 25566 27582 25618 27634
rect 45838 27582 45890 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 17502 27246 17554 27298
rect 21646 27246 21698 27298
rect 24446 27246 24498 27298
rect 26574 27246 26626 27298
rect 36990 27246 37042 27298
rect 37326 27246 37378 27298
rect 43038 27246 43090 27298
rect 9998 27134 10050 27186
rect 11118 27134 11170 27186
rect 11678 27134 11730 27186
rect 16606 27134 16658 27186
rect 20638 27134 20690 27186
rect 26686 27134 26738 27186
rect 27358 27134 27410 27186
rect 30494 27134 30546 27186
rect 32622 27134 32674 27186
rect 38446 27134 38498 27186
rect 38894 27134 38946 27186
rect 42702 27134 42754 27186
rect 4174 27022 4226 27074
rect 4846 27022 4898 27074
rect 5630 27022 5682 27074
rect 8094 27022 8146 27074
rect 8766 27022 8818 27074
rect 9326 27022 9378 27074
rect 9438 27022 9490 27074
rect 10782 27022 10834 27074
rect 11566 27022 11618 27074
rect 12014 27022 12066 27074
rect 13694 27022 13746 27074
rect 14142 27034 14194 27086
rect 17726 27022 17778 27074
rect 19630 27022 19682 27074
rect 19742 27022 19794 27074
rect 20302 27022 20354 27074
rect 21310 27022 21362 27074
rect 26910 27022 26962 27074
rect 30830 27022 30882 27074
rect 31278 27022 31330 27074
rect 32958 27022 33010 27074
rect 33966 27022 34018 27074
rect 34862 27022 34914 27074
rect 35086 27022 35138 27074
rect 37886 27022 37938 27074
rect 39230 27022 39282 27074
rect 39454 27022 39506 27074
rect 39902 27022 39954 27074
rect 40686 27022 40738 27074
rect 41246 27022 41298 27074
rect 41582 27022 41634 27074
rect 41918 27022 41970 27074
rect 42254 27022 42306 27074
rect 43374 27022 43426 27074
rect 44158 27022 44210 27074
rect 47182 27022 47234 27074
rect 2606 26910 2658 26962
rect 3838 26910 3890 26962
rect 4734 26910 4786 26962
rect 8990 26910 9042 26962
rect 9550 26910 9602 26962
rect 12686 26910 12738 26962
rect 16942 26910 16994 26962
rect 17166 26910 17218 26962
rect 23662 26910 23714 26962
rect 23774 26910 23826 26962
rect 24558 26910 24610 26962
rect 25118 26910 25170 26962
rect 29150 26910 29202 26962
rect 29486 26910 29538 26962
rect 31614 26910 31666 26962
rect 31838 26910 31890 26962
rect 35198 26910 35250 26962
rect 37214 26910 37266 26962
rect 37662 26910 37714 26962
rect 40126 26910 40178 26962
rect 44046 26910 44098 26962
rect 46398 26910 46450 26962
rect 46846 26910 46898 26962
rect 47406 26910 47458 26962
rect 47966 26910 48018 26962
rect 2270 26798 2322 26850
rect 17726 26798 17778 26850
rect 19854 26798 19906 26850
rect 21534 26798 21586 26850
rect 23438 26798 23490 26850
rect 30046 26798 30098 26850
rect 35646 26798 35698 26850
rect 39678 26798 39730 26850
rect 41134 26798 41186 26850
rect 42030 26798 42082 26850
rect 46062 26798 46114 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 8878 26462 8930 26514
rect 12462 26462 12514 26514
rect 14142 26462 14194 26514
rect 18510 26462 18562 26514
rect 19854 26462 19906 26514
rect 20750 26462 20802 26514
rect 24670 26462 24722 26514
rect 30830 26462 30882 26514
rect 32398 26462 32450 26514
rect 35310 26462 35362 26514
rect 39902 26462 39954 26514
rect 40350 26462 40402 26514
rect 40798 26462 40850 26514
rect 48302 26462 48354 26514
rect 9998 26350 10050 26402
rect 10110 26350 10162 26402
rect 10670 26350 10722 26402
rect 18846 26350 18898 26402
rect 20190 26350 20242 26402
rect 31502 26350 31554 26402
rect 33630 26350 33682 26402
rect 33966 26350 34018 26402
rect 37326 26350 37378 26402
rect 42030 26350 42082 26402
rect 42702 26350 42754 26402
rect 1822 26238 1874 26290
rect 2270 26238 2322 26290
rect 5182 26238 5234 26290
rect 10334 26238 10386 26290
rect 13806 26238 13858 26290
rect 14254 26238 14306 26290
rect 14478 26238 14530 26290
rect 14926 26238 14978 26290
rect 15150 26238 15202 26290
rect 17614 26238 17666 26290
rect 17838 26238 17890 26290
rect 19518 26238 19570 26290
rect 19854 26238 19906 26290
rect 21646 26238 21698 26290
rect 22206 26238 22258 26290
rect 25230 26238 25282 26290
rect 31166 26238 31218 26290
rect 31838 26238 31890 26290
rect 33406 26238 33458 26290
rect 40910 26238 40962 26290
rect 41918 26238 41970 26290
rect 43038 26238 43090 26290
rect 45166 26238 45218 26290
rect 45950 26238 46002 26290
rect 4734 26126 4786 26178
rect 8990 26126 9042 26178
rect 9662 26126 9714 26178
rect 11118 26126 11170 26178
rect 16606 26126 16658 26178
rect 17390 26126 17442 26178
rect 19294 26126 19346 26178
rect 28702 26126 28754 26178
rect 34414 26126 34466 26178
rect 35758 26126 35810 26178
rect 44942 26126 44994 26178
rect 8654 26014 8706 26066
rect 10446 26014 10498 26066
rect 10894 26014 10946 26066
rect 14814 26014 14866 26066
rect 18286 26014 18338 26066
rect 33070 26014 33122 26066
rect 37438 26014 37490 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 8654 25678 8706 25730
rect 18286 25678 18338 25730
rect 25902 25678 25954 25730
rect 31502 25678 31554 25730
rect 42702 25678 42754 25730
rect 45838 25678 45890 25730
rect 9662 25566 9714 25618
rect 12014 25566 12066 25618
rect 13582 25566 13634 25618
rect 23102 25566 23154 25618
rect 24222 25566 24274 25618
rect 26910 25566 26962 25618
rect 28030 25566 28082 25618
rect 29822 25566 29874 25618
rect 30830 25566 30882 25618
rect 36990 25566 37042 25618
rect 45390 25566 45442 25618
rect 8318 25454 8370 25506
rect 9214 25454 9266 25506
rect 10334 25454 10386 25506
rect 10894 25454 10946 25506
rect 12350 25454 12402 25506
rect 12910 25454 12962 25506
rect 13470 25454 13522 25506
rect 18398 25454 18450 25506
rect 18622 25454 18674 25506
rect 19742 25454 19794 25506
rect 22430 25454 22482 25506
rect 23214 25454 23266 25506
rect 23550 25454 23602 25506
rect 25342 25454 25394 25506
rect 25566 25454 25618 25506
rect 26126 25454 26178 25506
rect 26574 25454 26626 25506
rect 27022 25454 27074 25506
rect 27806 25454 27858 25506
rect 28142 25454 28194 25506
rect 28478 25454 28530 25506
rect 29374 25454 29426 25506
rect 30270 25454 30322 25506
rect 31838 25454 31890 25506
rect 39902 25454 39954 25506
rect 41918 25454 41970 25506
rect 43038 25454 43090 25506
rect 43598 25454 43650 25506
rect 46174 25454 46226 25506
rect 9886 25342 9938 25394
rect 9998 25342 10050 25394
rect 11342 25342 11394 25394
rect 11566 25342 11618 25394
rect 12686 25342 12738 25394
rect 13806 25342 13858 25394
rect 18286 25342 18338 25394
rect 19294 25342 19346 25394
rect 19966 25342 20018 25394
rect 21310 25342 21362 25394
rect 22318 25342 22370 25394
rect 22990 25342 23042 25394
rect 24446 25342 24498 25394
rect 24558 25342 24610 25394
rect 27134 25342 27186 25394
rect 31278 25342 31330 25394
rect 32734 25342 32786 25394
rect 39118 25342 39170 25394
rect 43822 25342 43874 25394
rect 46510 25342 46562 25394
rect 46958 25342 47010 25394
rect 8542 25230 8594 25282
rect 11230 25230 11282 25282
rect 12462 25230 12514 25282
rect 19070 25230 19122 25282
rect 19182 25230 19234 25282
rect 20414 25230 20466 25282
rect 21422 25230 21474 25282
rect 21534 25230 21586 25282
rect 21758 25230 21810 25282
rect 22094 25230 22146 25282
rect 24782 25230 24834 25282
rect 25454 25230 25506 25282
rect 26798 25230 26850 25282
rect 27694 25230 27746 25282
rect 31390 25230 31442 25282
rect 32174 25230 32226 25282
rect 32398 25230 32450 25282
rect 32622 25230 32674 25282
rect 40350 25230 40402 25282
rect 42254 25230 42306 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 9438 24894 9490 24946
rect 10894 24894 10946 24946
rect 14254 24894 14306 24946
rect 20750 24894 20802 24946
rect 1934 24670 1986 24722
rect 2606 24670 2658 24722
rect 7982 24670 8034 24722
rect 8542 24670 8594 24722
rect 8990 24670 9042 24722
rect 4958 24558 5010 24610
rect 5518 24558 5570 24610
rect 23998 24894 24050 24946
rect 27134 24894 27186 24946
rect 28814 24894 28866 24946
rect 29710 24894 29762 24946
rect 31054 24894 31106 24946
rect 40350 24894 40402 24946
rect 45166 24894 45218 24946
rect 9886 24782 9938 24834
rect 24222 24782 24274 24834
rect 26350 24782 26402 24834
rect 26798 24782 26850 24834
rect 30046 24782 30098 24834
rect 35758 24782 35810 24834
rect 36766 24782 36818 24834
rect 38558 24782 38610 24834
rect 40910 24782 40962 24834
rect 9774 24670 9826 24722
rect 11342 24670 11394 24722
rect 11902 24670 11954 24722
rect 14702 24670 14754 24722
rect 17502 24670 17554 24722
rect 18062 24670 18114 24722
rect 20414 24670 20466 24722
rect 20862 24670 20914 24722
rect 24670 24670 24722 24722
rect 27134 24670 27186 24722
rect 27470 24670 27522 24722
rect 29150 24670 29202 24722
rect 30382 24670 30434 24722
rect 30494 24670 30546 24722
rect 32286 24670 32338 24722
rect 35982 24670 36034 24722
rect 36542 24670 36594 24722
rect 38782 24670 38834 24722
rect 41134 24670 41186 24722
rect 42030 24670 42082 24722
rect 42702 24670 42754 24722
rect 10446 24558 10498 24610
rect 15150 24558 15202 24610
rect 24110 24558 24162 24610
rect 26462 24558 26514 24610
rect 27806 24558 27858 24610
rect 28254 24558 28306 24610
rect 30158 24558 30210 24610
rect 31614 24558 31666 24610
rect 32510 24558 32562 24610
rect 45614 24558 45666 24610
rect 9550 24446 9602 24498
rect 9886 24446 9938 24498
rect 10334 24446 10386 24498
rect 11006 24446 11058 24498
rect 31950 24446 32002 24498
rect 36318 24446 36370 24498
rect 41470 24446 41522 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12126 24110 12178 24162
rect 15486 24110 15538 24162
rect 22094 24110 22146 24162
rect 38334 24110 38386 24162
rect 38670 24110 38722 24162
rect 41358 24110 41410 24162
rect 5742 23998 5794 24050
rect 7758 23998 7810 24050
rect 8094 23998 8146 24050
rect 13582 23998 13634 24050
rect 26462 23998 26514 24050
rect 26798 23998 26850 24050
rect 28366 23998 28418 24050
rect 30942 23998 30994 24050
rect 31278 23998 31330 24050
rect 32622 23998 32674 24050
rect 33854 23998 33906 24050
rect 35982 23998 36034 24050
rect 36430 23998 36482 24050
rect 4174 23886 4226 23938
rect 4958 23886 5010 23938
rect 7870 23886 7922 23938
rect 8206 23886 8258 23938
rect 8430 23886 8482 23938
rect 9438 23886 9490 23938
rect 9998 23886 10050 23938
rect 10334 23886 10386 23938
rect 10558 23886 10610 23938
rect 10782 23886 10834 23938
rect 11678 23886 11730 23938
rect 12126 23886 12178 23938
rect 12238 23886 12290 23938
rect 14142 23886 14194 23938
rect 14478 23886 14530 23938
rect 14702 23886 14754 23938
rect 15150 23886 15202 23938
rect 16046 23886 16098 23938
rect 16382 23886 16434 23938
rect 23326 23886 23378 23938
rect 24110 23886 24162 23938
rect 29150 23886 29202 23938
rect 29598 23886 29650 23938
rect 33182 23886 33234 23938
rect 37102 23886 37154 23938
rect 37438 23886 37490 23938
rect 39230 23886 39282 23938
rect 40462 23886 40514 23938
rect 40686 23886 40738 23938
rect 41470 23886 41522 23938
rect 2606 23774 2658 23826
rect 2942 23774 2994 23826
rect 3838 23774 3890 23826
rect 4846 23774 4898 23826
rect 8990 23774 9042 23826
rect 9102 23774 9154 23826
rect 9550 23774 9602 23826
rect 14030 23774 14082 23826
rect 15374 23774 15426 23826
rect 15486 23774 15538 23826
rect 16718 23774 16770 23826
rect 17054 23774 17106 23826
rect 22206 23774 22258 23826
rect 30046 23774 30098 23826
rect 30382 23774 30434 23826
rect 32398 23774 32450 23826
rect 37998 23774 38050 23826
rect 38558 23774 38610 23826
rect 39678 23774 39730 23826
rect 41694 23774 41746 23826
rect 46734 23774 46786 23826
rect 8766 23662 8818 23714
rect 9774 23662 9826 23714
rect 10110 23662 10162 23714
rect 13806 23662 13858 23714
rect 14590 23662 14642 23714
rect 16270 23662 16322 23714
rect 17166 23662 17218 23714
rect 17614 23662 17666 23714
rect 27358 23662 27410 23714
rect 27806 23662 27858 23714
rect 32174 23662 32226 23714
rect 32622 23662 32674 23714
rect 46398 23662 46450 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 7982 23326 8034 23378
rect 9102 23326 9154 23378
rect 10222 23326 10274 23378
rect 10782 23326 10834 23378
rect 11678 23326 11730 23378
rect 12910 23326 12962 23378
rect 16830 23326 16882 23378
rect 23102 23326 23154 23378
rect 31054 23326 31106 23378
rect 34078 23326 34130 23378
rect 38782 23326 38834 23378
rect 48302 23326 48354 23378
rect 5854 23214 5906 23266
rect 6414 23214 6466 23266
rect 10446 23214 10498 23266
rect 11230 23214 11282 23266
rect 27022 23214 27074 23266
rect 27358 23214 27410 23266
rect 30158 23214 30210 23266
rect 31726 23214 31778 23266
rect 34526 23214 34578 23266
rect 36094 23214 36146 23266
rect 36542 23214 36594 23266
rect 36766 23214 36818 23266
rect 40350 23214 40402 23266
rect 42142 23214 42194 23266
rect 44158 23214 44210 23266
rect 44718 23214 44770 23266
rect 1822 23102 1874 23154
rect 2270 23102 2322 23154
rect 4734 23102 4786 23154
rect 5630 23102 5682 23154
rect 8206 23102 8258 23154
rect 8654 23102 8706 23154
rect 10110 23102 10162 23154
rect 10558 23102 10610 23154
rect 10894 23102 10946 23154
rect 12126 23102 12178 23154
rect 13022 23102 13074 23154
rect 13134 23102 13186 23154
rect 13582 23102 13634 23154
rect 13918 23102 13970 23154
rect 14478 23102 14530 23154
rect 17390 23102 17442 23154
rect 17950 23102 18002 23154
rect 20190 23102 20242 23154
rect 20750 23102 20802 23154
rect 26574 23102 26626 23154
rect 30270 23102 30322 23154
rect 31838 23102 31890 23154
rect 34750 23102 34802 23154
rect 35758 23102 35810 23154
rect 40126 23102 40178 23154
rect 41022 23102 41074 23154
rect 41358 23102 41410 23154
rect 41918 23102 41970 23154
rect 45166 23102 45218 23154
rect 45950 23102 46002 23154
rect 8094 22990 8146 23042
rect 9774 22990 9826 23042
rect 12574 22990 12626 23042
rect 26238 22990 26290 23042
rect 31950 22990 32002 23042
rect 32510 22990 32562 23042
rect 34190 22990 34242 23042
rect 37326 22990 37378 23042
rect 37998 22990 38050 23042
rect 39678 22990 39730 23042
rect 5294 22878 5346 22930
rect 12126 22878 12178 22930
rect 12686 22878 12738 22930
rect 30718 22878 30770 22930
rect 30942 22878 30994 22930
rect 34974 22878 35026 22930
rect 36878 22878 36930 22930
rect 43598 22878 43650 22930
rect 43934 22878 43986 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 9998 22542 10050 22594
rect 46846 22542 46898 22594
rect 47182 22542 47234 22594
rect 6302 22430 6354 22482
rect 10670 22430 10722 22482
rect 11678 22430 11730 22482
rect 12910 22430 12962 22482
rect 13582 22430 13634 22482
rect 17390 22430 17442 22482
rect 17726 22430 17778 22482
rect 23438 22430 23490 22482
rect 24222 22430 24274 22482
rect 25230 22430 25282 22482
rect 27918 22430 27970 22482
rect 35198 22430 35250 22482
rect 36206 22430 36258 22482
rect 37550 22430 37602 22482
rect 42814 22430 42866 22482
rect 43262 22430 43314 22482
rect 44942 22430 44994 22482
rect 45390 22430 45442 22482
rect 2606 22318 2658 22370
rect 4958 22318 5010 22370
rect 6526 22318 6578 22370
rect 7310 22318 7362 22370
rect 11566 22318 11618 22370
rect 12462 22318 12514 22370
rect 16942 22318 16994 22370
rect 20078 22318 20130 22370
rect 20862 22318 20914 22370
rect 21982 22318 22034 22370
rect 22990 22318 23042 22370
rect 24782 22318 24834 22370
rect 27470 22318 27522 22370
rect 28254 22318 28306 22370
rect 29486 22318 29538 22370
rect 29710 22318 29762 22370
rect 30158 22318 30210 22370
rect 30606 22318 30658 22370
rect 31502 22318 31554 22370
rect 31838 22318 31890 22370
rect 33966 22318 34018 22370
rect 34862 22318 34914 22370
rect 35870 22318 35922 22370
rect 37774 22318 37826 22370
rect 37998 22318 38050 22370
rect 39678 22318 39730 22370
rect 40350 22318 40402 22370
rect 43710 22318 43762 22370
rect 2270 22206 2322 22258
rect 9662 22206 9714 22258
rect 10110 22206 10162 22258
rect 11006 22206 11058 22258
rect 12126 22206 12178 22258
rect 29150 22206 29202 22258
rect 29598 22206 29650 22258
rect 30718 22206 30770 22258
rect 32174 22206 32226 22258
rect 33070 22206 33122 22258
rect 33742 22206 33794 22258
rect 34414 22206 34466 22258
rect 44046 22206 44098 22258
rect 47406 22206 47458 22258
rect 47966 22206 48018 22258
rect 5742 22094 5794 22146
rect 14030 22094 14082 22146
rect 22542 22094 22594 22146
rect 25790 22094 25842 22146
rect 27134 22094 27186 22146
rect 32734 22094 32786 22146
rect 37102 22094 37154 22146
rect 37214 22094 37266 22146
rect 37326 22094 37378 22146
rect 39006 22094 39058 22146
rect 39454 22094 39506 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 9102 21758 9154 21810
rect 10670 21758 10722 21810
rect 16494 21758 16546 21810
rect 23438 21758 23490 21810
rect 27806 21758 27858 21810
rect 31726 21758 31778 21810
rect 37102 21758 37154 21810
rect 47630 21758 47682 21810
rect 6414 21646 6466 21698
rect 9662 21646 9714 21698
rect 10334 21646 10386 21698
rect 18174 21646 18226 21698
rect 19070 21646 19122 21698
rect 21086 21646 21138 21698
rect 22206 21646 22258 21698
rect 23774 21646 23826 21698
rect 25454 21646 25506 21698
rect 26014 21646 26066 21698
rect 26798 21646 26850 21698
rect 27582 21646 27634 21698
rect 28254 21646 28306 21698
rect 29710 21646 29762 21698
rect 32286 21646 32338 21698
rect 33182 21646 33234 21698
rect 37774 21646 37826 21698
rect 37998 21646 38050 21698
rect 38334 21646 38386 21698
rect 39454 21646 39506 21698
rect 40126 21646 40178 21698
rect 47966 21646 48018 21698
rect 1934 21534 1986 21586
rect 2494 21534 2546 21586
rect 4846 21534 4898 21586
rect 5630 21534 5682 21586
rect 6302 21534 6354 21586
rect 9774 21534 9826 21586
rect 10782 21534 10834 21586
rect 11342 21534 11394 21586
rect 12238 21534 12290 21586
rect 13134 21534 13186 21586
rect 13582 21534 13634 21586
rect 16830 21534 16882 21586
rect 17726 21534 17778 21586
rect 19630 21534 19682 21586
rect 20190 21534 20242 21586
rect 22542 21534 22594 21586
rect 24334 21534 24386 21586
rect 25790 21534 25842 21586
rect 26686 21534 26738 21586
rect 28030 21534 28082 21586
rect 28702 21534 28754 21586
rect 29262 21534 29314 21586
rect 29598 21534 29650 21586
rect 31838 21534 31890 21586
rect 32174 21534 32226 21586
rect 33294 21534 33346 21586
rect 34078 21534 34130 21586
rect 34526 21534 34578 21586
rect 35758 21534 35810 21586
rect 36094 21534 36146 21586
rect 36318 21534 36370 21586
rect 37438 21534 37490 21586
rect 38446 21534 38498 21586
rect 38670 21534 38722 21586
rect 41134 21534 41186 21586
rect 42366 21534 42418 21586
rect 42814 21534 42866 21586
rect 44494 21534 44546 21586
rect 45166 21534 45218 21586
rect 48190 21534 48242 21586
rect 6974 21422 7026 21474
rect 12686 21422 12738 21474
rect 16046 21422 16098 21474
rect 18510 21422 18562 21474
rect 20526 21422 20578 21474
rect 22878 21422 22930 21474
rect 26574 21422 26626 21474
rect 28366 21422 28418 21474
rect 33630 21422 33682 21474
rect 39342 21422 39394 21474
rect 40126 21422 40178 21474
rect 43038 21422 43090 21474
rect 5294 21310 5346 21362
rect 29710 21310 29762 21362
rect 31726 21310 31778 21362
rect 32286 21310 32338 21362
rect 37214 21310 37266 21362
rect 38782 21310 38834 21362
rect 39230 21310 39282 21362
rect 39902 21310 39954 21362
rect 43598 21310 43650 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 6414 20974 6466 21026
rect 13582 20974 13634 21026
rect 14254 20974 14306 21026
rect 14366 20974 14418 21026
rect 15150 20974 15202 21026
rect 25342 20974 25394 21026
rect 25902 20974 25954 21026
rect 26126 20974 26178 21026
rect 34190 20974 34242 21026
rect 43486 20974 43538 21026
rect 5070 20862 5122 20914
rect 8990 20862 9042 20914
rect 9326 20862 9378 20914
rect 15262 20862 15314 20914
rect 19518 20862 19570 20914
rect 20638 20862 20690 20914
rect 22094 20862 22146 20914
rect 23998 20862 24050 20914
rect 26686 20862 26738 20914
rect 28254 20862 28306 20914
rect 31054 20862 31106 20914
rect 31950 20862 32002 20914
rect 36990 20862 37042 20914
rect 41582 20862 41634 20914
rect 44046 20862 44098 20914
rect 44942 20862 44994 20914
rect 48302 20862 48354 20914
rect 2942 20750 2994 20802
rect 9998 20750 10050 20802
rect 10558 20750 10610 20802
rect 11566 20750 11618 20802
rect 12126 20750 12178 20802
rect 13806 20750 13858 20802
rect 14814 20750 14866 20802
rect 18062 20750 18114 20802
rect 22318 20750 22370 20802
rect 22990 20750 23042 20802
rect 24782 20750 24834 20802
rect 25566 20750 25618 20802
rect 26462 20750 26514 20802
rect 26574 20750 26626 20802
rect 27246 20750 27298 20802
rect 27806 20750 27858 20802
rect 29822 20750 29874 20802
rect 30046 20750 30098 20802
rect 30270 20750 30322 20802
rect 30494 20750 30546 20802
rect 30830 20750 30882 20802
rect 31166 20750 31218 20802
rect 33406 20750 33458 20802
rect 33742 20750 33794 20802
rect 34862 20750 34914 20802
rect 37326 20750 37378 20802
rect 37886 20750 37938 20802
rect 39230 20750 39282 20802
rect 40126 20750 40178 20802
rect 42926 20750 42978 20802
rect 43822 20750 43874 20802
rect 45166 20750 45218 20802
rect 45950 20750 46002 20802
rect 2606 20638 2658 20690
rect 6638 20638 6690 20690
rect 6974 20638 7026 20690
rect 9662 20638 9714 20690
rect 10782 20638 10834 20690
rect 11118 20638 11170 20690
rect 14142 20638 14194 20690
rect 23438 20638 23490 20690
rect 25006 20638 25058 20690
rect 31502 20638 31554 20690
rect 32286 20638 32338 20690
rect 32398 20638 32450 20690
rect 32622 20638 32674 20690
rect 32846 20638 32898 20690
rect 33518 20638 33570 20690
rect 34526 20638 34578 20690
rect 34974 20638 35026 20690
rect 38446 20638 38498 20690
rect 6078 20526 6130 20578
rect 8094 20526 8146 20578
rect 8430 20526 8482 20578
rect 11454 20526 11506 20578
rect 17054 20526 17106 20578
rect 21534 20526 21586 20578
rect 22430 20526 22482 20578
rect 22654 20526 22706 20578
rect 24446 20526 24498 20578
rect 25230 20526 25282 20578
rect 26798 20526 26850 20578
rect 30606 20526 30658 20578
rect 32958 20526 33010 20578
rect 33182 20526 33234 20578
rect 34302 20526 34354 20578
rect 35198 20526 35250 20578
rect 37998 20526 38050 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 25902 20190 25954 20242
rect 27246 20190 27298 20242
rect 28702 20190 28754 20242
rect 39118 20190 39170 20242
rect 43822 20190 43874 20242
rect 5630 20078 5682 20130
rect 8990 20078 9042 20130
rect 13918 20078 13970 20130
rect 14366 20078 14418 20130
rect 15150 20078 15202 20130
rect 23886 20078 23938 20130
rect 25342 20078 25394 20130
rect 26798 20078 26850 20130
rect 27806 20078 27858 20130
rect 29710 20078 29762 20130
rect 29822 20078 29874 20130
rect 29934 20078 29986 20130
rect 30382 20078 30434 20130
rect 32174 20078 32226 20130
rect 32398 20078 32450 20130
rect 35534 20078 35586 20130
rect 36430 20078 36482 20130
rect 39678 20078 39730 20130
rect 40014 20078 40066 20130
rect 44158 20078 44210 20130
rect 5406 19966 5458 20018
rect 5854 19966 5906 20018
rect 6526 19966 6578 20018
rect 9998 19966 10050 20018
rect 10446 19966 10498 20018
rect 13358 19966 13410 20018
rect 14702 19966 14754 20018
rect 16830 19966 16882 20018
rect 18174 19966 18226 20018
rect 21310 19966 21362 20018
rect 22542 19966 22594 20018
rect 23438 19966 23490 20018
rect 25902 19966 25954 20018
rect 26910 19966 26962 20018
rect 27358 19966 27410 20018
rect 28254 19966 28306 20018
rect 29038 19966 29090 20018
rect 29262 19966 29314 20018
rect 30270 19966 30322 20018
rect 32510 19966 32562 20018
rect 33406 19966 33458 20018
rect 33742 19965 33794 20017
rect 34414 19966 34466 20018
rect 36206 19966 36258 20018
rect 38110 19966 38162 20018
rect 42926 19966 42978 20018
rect 44270 19966 44322 20018
rect 45390 19966 45442 20018
rect 46062 19966 46114 20018
rect 46286 19966 46338 20018
rect 11006 19854 11058 19906
rect 16270 19854 16322 19906
rect 17614 19854 17666 19906
rect 18846 19854 18898 19906
rect 20974 19854 21026 19906
rect 33630 19854 33682 19906
rect 36430 19854 36482 19906
rect 38558 19854 38610 19906
rect 41918 19854 41970 19906
rect 24558 19742 24610 19794
rect 39454 19742 39506 19794
rect 44606 19742 44658 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 28030 19406 28082 19458
rect 37214 19406 37266 19458
rect 43150 19406 43202 19458
rect 45502 19406 45554 19458
rect 48078 19406 48130 19458
rect 5742 19294 5794 19346
rect 7310 19294 7362 19346
rect 8430 19294 8482 19346
rect 8990 19294 9042 19346
rect 10558 19294 10610 19346
rect 17278 19294 17330 19346
rect 19966 19294 20018 19346
rect 20750 19294 20802 19346
rect 23998 19294 24050 19346
rect 26014 19294 26066 19346
rect 26798 19294 26850 19346
rect 28590 19294 28642 19346
rect 29598 19294 29650 19346
rect 33406 19294 33458 19346
rect 35982 19294 36034 19346
rect 37662 19294 37714 19346
rect 39342 19294 39394 19346
rect 41806 19294 41858 19346
rect 42590 19294 42642 19346
rect 43486 19294 43538 19346
rect 45278 19294 45330 19346
rect 1822 19182 1874 19234
rect 2270 19182 2322 19234
rect 6862 19182 6914 19234
rect 9998 19182 10050 19234
rect 12798 19182 12850 19234
rect 13694 19182 13746 19234
rect 14366 19182 14418 19234
rect 18062 19182 18114 19234
rect 21422 19182 21474 19234
rect 21982 19182 22034 19234
rect 22430 19182 22482 19234
rect 24110 19182 24162 19234
rect 26686 19182 26738 19234
rect 28366 19182 28418 19234
rect 29150 19182 29202 19234
rect 30830 19182 30882 19234
rect 34526 19182 34578 19234
rect 36430 19182 36482 19234
rect 37102 19182 37154 19234
rect 37550 19182 37602 19234
rect 40350 19182 40402 19234
rect 41022 19182 41074 19234
rect 42814 19182 42866 19234
rect 43710 19182 43762 19234
rect 45054 19182 45106 19234
rect 46286 19182 46338 19234
rect 47742 19182 47794 19234
rect 6302 19070 6354 19122
rect 9438 19070 9490 19122
rect 9550 19070 9602 19122
rect 15150 19070 15202 19122
rect 22990 19070 23042 19122
rect 24222 19070 24274 19122
rect 27358 19070 27410 19122
rect 27694 19070 27746 19122
rect 29374 19070 29426 19122
rect 31950 19070 32002 19122
rect 33966 19070 34018 19122
rect 37774 19070 37826 19122
rect 45838 19070 45890 19122
rect 47182 19070 47234 19122
rect 47406 19070 47458 19122
rect 4734 18958 4786 19010
rect 9214 18958 9266 19010
rect 9326 18958 9378 19010
rect 13470 18958 13522 19010
rect 34974 18958 35026 19010
rect 35310 18958 35362 19010
rect 44046 18958 44098 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 2270 18622 2322 18674
rect 14926 18622 14978 18674
rect 25566 18622 25618 18674
rect 27694 18622 27746 18674
rect 29262 18622 29314 18674
rect 29486 18622 29538 18674
rect 32510 18622 32562 18674
rect 34078 18622 34130 18674
rect 37438 18622 37490 18674
rect 43598 18622 43650 18674
rect 5182 18510 5234 18562
rect 6750 18510 6802 18562
rect 19294 18510 19346 18562
rect 25230 18510 25282 18562
rect 28590 18510 28642 18562
rect 29038 18510 29090 18562
rect 29598 18510 29650 18562
rect 34302 18510 34354 18562
rect 36654 18510 36706 18562
rect 36990 18510 37042 18562
rect 41022 18510 41074 18562
rect 42814 18510 42866 18562
rect 44942 18510 44994 18562
rect 2606 18398 2658 18450
rect 4062 18398 4114 18450
rect 4398 18398 4450 18450
rect 4846 18398 4898 18450
rect 6414 18398 6466 18450
rect 9998 18398 10050 18450
rect 10334 18398 10386 18450
rect 10670 18398 10722 18450
rect 10894 18398 10946 18450
rect 11454 18398 11506 18450
rect 11790 18398 11842 18450
rect 12350 18398 12402 18450
rect 12462 18398 12514 18450
rect 14254 18398 14306 18450
rect 14702 18398 14754 18450
rect 15262 18398 15314 18450
rect 15710 18398 15762 18450
rect 17950 18398 18002 18450
rect 18286 18398 18338 18450
rect 19630 18398 19682 18450
rect 20414 18398 20466 18450
rect 24558 18398 24610 18450
rect 26462 18398 26514 18450
rect 26686 18398 26738 18450
rect 26910 18398 26962 18450
rect 28814 18398 28866 18450
rect 30494 18398 30546 18450
rect 30942 18398 30994 18450
rect 31950 18398 32002 18450
rect 33182 18398 33234 18450
rect 33406 18398 33458 18450
rect 34190 18398 34242 18450
rect 35534 18398 35586 18450
rect 36430 18398 36482 18450
rect 37214 18398 37266 18450
rect 37550 18398 37602 18450
rect 37998 18398 38050 18450
rect 38222 18398 38274 18450
rect 38334 18398 38386 18450
rect 38670 18398 38722 18450
rect 39006 18398 39058 18450
rect 39230 18398 39282 18450
rect 39454 18398 39506 18450
rect 39678 18398 39730 18450
rect 40910 18398 40962 18450
rect 41918 18398 41970 18450
rect 43038 18398 43090 18450
rect 44718 18398 44770 18450
rect 45166 18398 45218 18450
rect 45838 18398 45890 18450
rect 9774 18286 9826 18338
rect 10782 18286 10834 18338
rect 12238 18286 12290 18338
rect 13134 18286 13186 18338
rect 13806 18286 13858 18338
rect 18398 18286 18450 18338
rect 20862 18286 20914 18338
rect 22094 18286 22146 18338
rect 23774 18286 23826 18338
rect 24110 18286 24162 18338
rect 31278 18286 31330 18338
rect 35086 18286 35138 18338
rect 35982 18286 36034 18338
rect 40014 18286 40066 18338
rect 42366 18286 42418 18338
rect 44046 18286 44098 18338
rect 48302 18286 48354 18338
rect 10446 18174 10498 18226
rect 12014 18174 12066 18226
rect 14030 18174 14082 18226
rect 17726 18174 17778 18226
rect 28702 18174 28754 18226
rect 37438 18174 37490 18226
rect 41022 18174 41074 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 4174 17838 4226 17890
rect 6190 17838 6242 17890
rect 9102 17838 9154 17890
rect 11790 17838 11842 17890
rect 16046 17838 16098 17890
rect 17950 17838 18002 17890
rect 18958 17838 19010 17890
rect 45726 17838 45778 17890
rect 46062 17838 46114 17890
rect 8542 17726 8594 17778
rect 11118 17726 11170 17778
rect 12126 17726 12178 17778
rect 12910 17726 12962 17778
rect 13582 17726 13634 17778
rect 14702 17726 14754 17778
rect 19182 17726 19234 17778
rect 19406 17726 19458 17778
rect 23662 17726 23714 17778
rect 29934 17726 29986 17778
rect 32174 17726 32226 17778
rect 32734 17726 32786 17778
rect 34750 17726 34802 17778
rect 35534 17726 35586 17778
rect 37214 17726 37266 17778
rect 39902 17726 39954 17778
rect 40798 17726 40850 17778
rect 44270 17726 44322 17778
rect 45054 17726 45106 17778
rect 4622 17614 4674 17666
rect 6526 17614 6578 17666
rect 8766 17614 8818 17666
rect 9326 17614 9378 17666
rect 9662 17614 9714 17666
rect 9886 17614 9938 17666
rect 10110 17614 10162 17666
rect 11230 17614 11282 17666
rect 11566 17614 11618 17666
rect 12014 17614 12066 17666
rect 15822 17614 15874 17666
rect 16158 17614 16210 17666
rect 17054 17614 17106 17666
rect 17390 17614 17442 17666
rect 17614 17614 17666 17666
rect 18734 17614 18786 17666
rect 20414 17614 20466 17666
rect 21198 17614 21250 17666
rect 21534 17614 21586 17666
rect 23214 17614 23266 17666
rect 27022 17614 27074 17666
rect 27470 17614 27522 17666
rect 28254 17614 28306 17666
rect 29486 17614 29538 17666
rect 30606 17614 30658 17666
rect 30830 17614 30882 17666
rect 31054 17614 31106 17666
rect 33182 17614 33234 17666
rect 33518 17614 33570 17666
rect 35422 17614 35474 17666
rect 39006 17614 39058 17666
rect 40574 17614 40626 17666
rect 41134 17614 41186 17666
rect 41806 17614 41858 17666
rect 46734 17614 46786 17666
rect 2494 17502 2546 17554
rect 3838 17502 3890 17554
rect 4958 17502 5010 17554
rect 6750 17502 6802 17554
rect 7086 17502 7138 17554
rect 10334 17502 10386 17554
rect 12238 17502 12290 17554
rect 13694 17502 13746 17554
rect 13806 17502 13858 17554
rect 13918 17502 13970 17554
rect 20078 17502 20130 17554
rect 21758 17502 21810 17554
rect 21870 17502 21922 17554
rect 22094 17502 22146 17554
rect 24446 17502 24498 17554
rect 26910 17502 26962 17554
rect 27694 17502 27746 17554
rect 28478 17502 28530 17554
rect 28590 17502 28642 17554
rect 29150 17502 29202 17554
rect 33070 17502 33122 17554
rect 35646 17502 35698 17554
rect 46622 17502 46674 17554
rect 2158 17390 2210 17442
rect 9886 17390 9938 17442
rect 13470 17390 13522 17442
rect 16158 17390 16210 17442
rect 16718 17390 16770 17442
rect 18286 17390 18338 17442
rect 20190 17390 20242 17442
rect 22206 17390 22258 17442
rect 22430 17390 22482 17442
rect 22878 17390 22930 17442
rect 27470 17390 27522 17442
rect 30942 17390 30994 17442
rect 31278 17390 31330 17442
rect 31726 17390 31778 17442
rect 34190 17390 34242 17442
rect 35198 17390 35250 17442
rect 36094 17390 36146 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 4734 17054 4786 17106
rect 9662 17054 9714 17106
rect 10894 17054 10946 17106
rect 11342 17054 11394 17106
rect 12462 17054 12514 17106
rect 13022 17054 13074 17106
rect 13470 17054 13522 17106
rect 14030 17054 14082 17106
rect 14254 17054 14306 17106
rect 15374 17054 15426 17106
rect 18286 17054 18338 17106
rect 19070 17054 19122 17106
rect 19854 17054 19906 17106
rect 27358 17054 27410 17106
rect 28254 17054 28306 17106
rect 29934 17054 29986 17106
rect 35198 17054 35250 17106
rect 36094 17054 36146 17106
rect 36990 17054 37042 17106
rect 37438 17054 37490 17106
rect 37662 17054 37714 17106
rect 37774 17054 37826 17106
rect 38222 17054 38274 17106
rect 40014 17054 40066 17106
rect 40910 17054 40962 17106
rect 41358 17054 41410 17106
rect 41918 17054 41970 17106
rect 42366 17054 42418 17106
rect 42814 17054 42866 17106
rect 47294 17054 47346 17106
rect 8990 16942 9042 16994
rect 11902 16942 11954 16994
rect 14590 16942 14642 16994
rect 15486 16942 15538 16994
rect 16046 16942 16098 16994
rect 16494 16942 16546 16994
rect 16830 16942 16882 16994
rect 17614 16942 17666 16994
rect 20190 16942 20242 16994
rect 20974 16942 21026 16994
rect 21310 16942 21362 16994
rect 21758 16942 21810 16994
rect 25230 16942 25282 16994
rect 27470 16942 27522 16994
rect 27918 16942 27970 16994
rect 28478 16942 28530 16994
rect 30046 16942 30098 16994
rect 30382 16942 30434 16994
rect 31502 16942 31554 16994
rect 33742 16942 33794 16994
rect 34190 16942 34242 16994
rect 34302 16942 34354 16994
rect 38558 16942 38610 16994
rect 39454 16942 39506 16994
rect 41470 16942 41522 16994
rect 43822 16942 43874 16994
rect 45726 16942 45778 16994
rect 46062 16942 46114 16994
rect 1710 16830 1762 16882
rect 2270 16830 2322 16882
rect 5854 16830 5906 16882
rect 6638 16830 6690 16882
rect 17838 16830 17890 16882
rect 18062 16830 18114 16882
rect 18286 16830 18338 16882
rect 19294 16830 19346 16882
rect 20414 16830 20466 16882
rect 20750 16830 20802 16882
rect 22430 16830 22482 16882
rect 23326 16830 23378 16882
rect 23774 16830 23826 16882
rect 24334 16830 24386 16882
rect 27694 16830 27746 16882
rect 28030 16830 28082 16882
rect 28590 16830 28642 16882
rect 30942 16830 30994 16882
rect 31166 16830 31218 16882
rect 31726 16830 31778 16882
rect 33182 16830 33234 16882
rect 35534 16830 35586 16882
rect 36318 16830 36370 16882
rect 36766 16830 36818 16882
rect 37886 16830 37938 16882
rect 38894 16830 38946 16882
rect 41022 16830 41074 16882
rect 43598 16830 43650 16882
rect 46734 16830 46786 16882
rect 5182 16718 5234 16770
rect 10222 16718 10274 16770
rect 18846 16718 18898 16770
rect 19182 16718 19234 16770
rect 20078 16718 20130 16770
rect 21646 16718 21698 16770
rect 21982 16718 22034 16770
rect 22766 16718 22818 16770
rect 25454 16718 25506 16770
rect 33518 16718 33570 16770
rect 34638 16718 34690 16770
rect 34862 16718 34914 16770
rect 35758 16718 35810 16770
rect 36878 16718 36930 16770
rect 39902 16718 39954 16770
rect 44718 16718 44770 16770
rect 47742 16718 47794 16770
rect 10222 16606 10274 16658
rect 11566 16606 11618 16658
rect 12126 16606 12178 16658
rect 15374 16606 15426 16658
rect 15822 16606 15874 16658
rect 16158 16606 16210 16658
rect 18622 16606 18674 16658
rect 22990 16606 23042 16658
rect 27358 16606 27410 16658
rect 29934 16606 29986 16658
rect 31950 16606 32002 16658
rect 32174 16606 32226 16658
rect 32622 16606 32674 16658
rect 34190 16606 34242 16658
rect 39790 16606 39842 16658
rect 43150 16606 43202 16658
rect 45166 16606 45218 16658
rect 45502 16606 45554 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 4174 16270 4226 16322
rect 27134 16270 27186 16322
rect 37326 16270 37378 16322
rect 43262 16270 43314 16322
rect 8318 16158 8370 16210
rect 8878 16158 8930 16210
rect 9998 16158 10050 16210
rect 11118 16158 11170 16210
rect 11566 16158 11618 16210
rect 12798 16158 12850 16210
rect 28366 16158 28418 16210
rect 29374 16158 29426 16210
rect 30494 16158 30546 16210
rect 31278 16158 31330 16210
rect 35982 16158 36034 16210
rect 36990 16158 37042 16210
rect 38110 16158 38162 16210
rect 39118 16158 39170 16210
rect 41246 16158 41298 16210
rect 41694 16158 41746 16210
rect 48302 16158 48354 16210
rect 4846 16046 4898 16098
rect 8542 16046 8594 16098
rect 14702 16046 14754 16098
rect 15822 16046 15874 16098
rect 16270 16046 16322 16098
rect 17614 16046 17666 16098
rect 19406 16046 19458 16098
rect 22430 16046 22482 16098
rect 23998 16046 24050 16098
rect 26462 16046 26514 16098
rect 27022 16046 27074 16098
rect 28254 16046 28306 16098
rect 29486 16046 29538 16098
rect 33406 16046 33458 16098
rect 33742 16046 33794 16098
rect 35870 16046 35922 16098
rect 36542 16046 36594 16098
rect 38446 16046 38498 16098
rect 43710 16046 43762 16098
rect 45166 16046 45218 16098
rect 45838 16046 45890 16098
rect 4958 15934 5010 15986
rect 9550 15934 9602 15986
rect 9662 15934 9714 15986
rect 10670 15934 10722 15986
rect 10782 15934 10834 15986
rect 15374 15934 15426 15986
rect 16830 15934 16882 15986
rect 17950 15934 18002 15986
rect 18510 15934 18562 15986
rect 18958 15934 19010 15986
rect 22318 15934 22370 15986
rect 25678 15934 25730 15986
rect 30158 15934 30210 15986
rect 31838 15934 31890 15986
rect 34302 15934 34354 15986
rect 36094 15934 36146 15986
rect 37550 15934 37602 15986
rect 43822 15934 43874 15986
rect 3838 15822 3890 15874
rect 9214 15822 9266 15874
rect 9438 15822 9490 15874
rect 10334 15822 10386 15874
rect 10558 15822 10610 15874
rect 14926 15822 14978 15874
rect 16270 15822 16322 15874
rect 19294 15822 19346 15874
rect 20414 15822 20466 15874
rect 20862 15822 20914 15874
rect 21646 15822 21698 15874
rect 21982 15822 22034 15874
rect 24894 15822 24946 15874
rect 27134 15822 27186 15874
rect 27806 15822 27858 15874
rect 30606 15822 30658 15874
rect 33182 15822 33234 15874
rect 42926 15822 42978 15874
rect 45054 15822 45106 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 5070 15486 5122 15538
rect 10222 15486 10274 15538
rect 20078 15486 20130 15538
rect 26910 15486 26962 15538
rect 36206 15486 36258 15538
rect 36318 15486 36370 15538
rect 39006 15486 39058 15538
rect 44830 15486 44882 15538
rect 45838 15486 45890 15538
rect 46622 15486 46674 15538
rect 2158 15374 2210 15426
rect 2494 15374 2546 15426
rect 4286 15374 4338 15426
rect 9662 15374 9714 15426
rect 16494 15374 16546 15426
rect 20414 15374 20466 15426
rect 21422 15374 21474 15426
rect 25902 15374 25954 15426
rect 27022 15374 27074 15426
rect 34974 15374 35026 15426
rect 38782 15374 38834 15426
rect 45502 15374 45554 15426
rect 4622 15262 4674 15314
rect 11678 15262 11730 15314
rect 14926 15262 14978 15314
rect 15374 15262 15426 15314
rect 15598 15262 15650 15314
rect 15822 15262 15874 15314
rect 16046 15262 16098 15314
rect 19630 15262 19682 15314
rect 19854 15262 19906 15314
rect 20638 15262 20690 15314
rect 21982 15262 22034 15314
rect 22206 15262 22258 15314
rect 23550 15262 23602 15314
rect 25342 15262 25394 15314
rect 25566 15262 25618 15314
rect 27806 15262 27858 15314
rect 29934 15262 29986 15314
rect 30494 15262 30546 15314
rect 30942 15262 30994 15314
rect 31502 15262 31554 15314
rect 32286 15262 32338 15314
rect 33182 15262 33234 15314
rect 33406 15262 33458 15314
rect 33742 15262 33794 15314
rect 34414 15262 34466 15314
rect 34638 15262 34690 15314
rect 35758 15262 35810 15314
rect 36094 15262 36146 15314
rect 36654 15262 36706 15314
rect 36990 15262 37042 15314
rect 37550 15262 37602 15314
rect 37886 15262 37938 15314
rect 41694 15262 41746 15314
rect 42478 15262 42530 15314
rect 47294 15262 47346 15314
rect 12350 15150 12402 15202
rect 14478 15150 14530 15202
rect 19742 15150 19794 15202
rect 21870 15150 21922 15202
rect 23214 15150 23266 15202
rect 24670 15150 24722 15202
rect 35310 15150 35362 15202
rect 38110 15150 38162 15202
rect 38334 15150 38386 15202
rect 38446 15150 38498 15202
rect 38894 15150 38946 15202
rect 39566 15150 39618 15202
rect 46958 15150 47010 15202
rect 9886 15038 9938 15090
rect 15262 15038 15314 15090
rect 16382 15038 16434 15090
rect 23438 15038 23490 15090
rect 26014 15038 26066 15090
rect 26126 15038 26178 15090
rect 31726 15038 31778 15090
rect 37214 15038 37266 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 5742 14702 5794 14754
rect 6078 14702 6130 14754
rect 12574 14702 12626 14754
rect 19742 14702 19794 14754
rect 20638 14702 20690 14754
rect 21198 14702 21250 14754
rect 44942 14702 44994 14754
rect 45390 14702 45442 14754
rect 47182 14702 47234 14754
rect 11006 14590 11058 14642
rect 11566 14590 11618 14642
rect 25342 14590 25394 14642
rect 26462 14590 26514 14642
rect 27470 14590 27522 14642
rect 35646 14590 35698 14642
rect 36206 14590 36258 14642
rect 37886 14590 37938 14642
rect 39118 14590 39170 14642
rect 41246 14590 41298 14642
rect 44942 14590 44994 14642
rect 45390 14590 45442 14642
rect 1710 14478 1762 14530
rect 2270 14478 2322 14530
rect 7422 14478 7474 14530
rect 7870 14478 7922 14530
rect 8542 14478 8594 14530
rect 17166 14478 17218 14530
rect 17278 14478 17330 14530
rect 17726 14478 17778 14530
rect 19406 14478 19458 14530
rect 20078 14478 20130 14530
rect 20302 14478 20354 14530
rect 21534 14478 21586 14530
rect 22430 14478 22482 14530
rect 22990 14478 23042 14530
rect 23550 14478 23602 14530
rect 24334 14478 24386 14530
rect 25230 14478 25282 14530
rect 26014 14478 26066 14530
rect 26238 14478 26290 14530
rect 27582 14478 27634 14530
rect 27918 14478 27970 14530
rect 29822 14478 29874 14530
rect 30382 14478 30434 14530
rect 31390 14478 31442 14530
rect 33406 14478 33458 14530
rect 37438 14478 37490 14530
rect 38446 14478 38498 14530
rect 42814 14478 42866 14530
rect 6302 14366 6354 14418
rect 6862 14366 6914 14418
rect 7646 14366 7698 14418
rect 12910 14366 12962 14418
rect 17054 14366 17106 14418
rect 18734 14366 18786 14418
rect 20750 14366 20802 14418
rect 21310 14366 21362 14418
rect 21758 14366 21810 14418
rect 22766 14366 22818 14418
rect 23998 14366 24050 14418
rect 24110 14366 24162 14418
rect 28366 14366 28418 14418
rect 31054 14366 31106 14418
rect 31502 14366 31554 14418
rect 33966 14366 34018 14418
rect 35534 14366 35586 14418
rect 36990 14366 37042 14418
rect 42478 14366 42530 14418
rect 47406 14366 47458 14418
rect 47742 14366 47794 14418
rect 4734 14254 4786 14306
rect 12686 14254 12738 14306
rect 14366 14254 14418 14306
rect 16606 14254 16658 14306
rect 18062 14254 18114 14306
rect 18622 14254 18674 14306
rect 18958 14254 19010 14306
rect 19182 14254 19234 14306
rect 22094 14254 22146 14306
rect 27358 14254 27410 14306
rect 28478 14254 28530 14306
rect 28702 14254 28754 14306
rect 32398 14254 32450 14306
rect 36878 14254 36930 14306
rect 37214 14254 37266 14306
rect 41694 14254 41746 14306
rect 46846 14254 46898 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 6526 13918 6578 13970
rect 6974 13918 7026 13970
rect 7422 13918 7474 13970
rect 15710 13918 15762 13970
rect 21310 13918 21362 13970
rect 25230 13918 25282 13970
rect 28254 13918 28306 13970
rect 34526 13918 34578 13970
rect 36094 13918 36146 13970
rect 36990 13918 37042 13970
rect 37886 13918 37938 13970
rect 41134 13918 41186 13970
rect 45166 13918 45218 13970
rect 45502 13918 45554 13970
rect 48302 13918 48354 13970
rect 7982 13806 8034 13858
rect 8430 13806 8482 13858
rect 12014 13806 12066 13858
rect 15262 13806 15314 13858
rect 15934 13806 15986 13858
rect 17390 13806 17442 13858
rect 17838 13806 17890 13858
rect 19070 13806 19122 13858
rect 20526 13806 20578 13858
rect 21198 13806 21250 13858
rect 25566 13806 25618 13858
rect 26686 13806 26738 13858
rect 29262 13806 29314 13858
rect 31838 13806 31890 13858
rect 34078 13806 34130 13858
rect 34862 13806 34914 13858
rect 35198 13806 35250 13858
rect 46398 13806 46450 13858
rect 3614 13694 3666 13746
rect 4174 13694 4226 13746
rect 7758 13694 7810 13746
rect 11342 13694 11394 13746
rect 16158 13694 16210 13746
rect 17614 13694 17666 13746
rect 19518 13694 19570 13746
rect 20078 13694 20130 13746
rect 21422 13694 21474 13746
rect 21870 13694 21922 13746
rect 26462 13694 26514 13746
rect 27246 13694 27298 13746
rect 27694 13694 27746 13746
rect 28590 13694 28642 13746
rect 29150 13694 29202 13746
rect 30830 13694 30882 13746
rect 31054 13694 31106 13746
rect 33630 13694 33682 13746
rect 35758 13694 35810 13746
rect 37326 13694 37378 13746
rect 38222 13694 38274 13746
rect 45838 13694 45890 13746
rect 46510 13694 46562 13746
rect 14142 13582 14194 13634
rect 15038 13582 15090 13634
rect 15486 13582 15538 13634
rect 17502 13582 17554 13634
rect 19630 13582 19682 13634
rect 22542 13582 22594 13634
rect 24670 13582 24722 13634
rect 26126 13582 26178 13634
rect 33182 13582 33234 13634
rect 36542 13582 36594 13634
rect 38670 13582 38722 13634
rect 15710 13470 15762 13522
rect 27582 13470 27634 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 7982 13134 8034 13186
rect 15374 13134 15426 13186
rect 28254 13134 28306 13186
rect 28590 13134 28642 13186
rect 6190 13022 6242 13074
rect 6750 13022 6802 13074
rect 12798 13022 12850 13074
rect 13470 13022 13522 13074
rect 14366 13022 14418 13074
rect 14814 13022 14866 13074
rect 16382 13022 16434 13074
rect 21646 13022 21698 13074
rect 24558 13022 24610 13074
rect 29598 13022 29650 13074
rect 30270 13022 30322 13074
rect 31166 13022 31218 13074
rect 32286 13022 32338 13074
rect 32734 13022 32786 13074
rect 33182 13022 33234 13074
rect 33742 13022 33794 13074
rect 34078 13022 34130 13074
rect 34974 13022 35026 13074
rect 35198 13022 35250 13074
rect 36318 13022 36370 13074
rect 37998 13022 38050 13074
rect 44270 13022 44322 13074
rect 48302 13022 48354 13074
rect 4174 12910 4226 12962
rect 4958 12910 5010 12962
rect 5742 12910 5794 12962
rect 8430 12910 8482 12962
rect 14142 12910 14194 12962
rect 15038 12910 15090 12962
rect 15710 12910 15762 12962
rect 16942 12910 16994 12962
rect 17390 12910 17442 12962
rect 17838 12910 17890 12962
rect 25006 12910 25058 12962
rect 25678 12910 25730 12962
rect 26462 12910 26514 12962
rect 27358 12910 27410 12962
rect 27918 12910 27970 12962
rect 29262 12910 29314 12962
rect 30718 12910 30770 12962
rect 31950 12910 32002 12962
rect 33854 12910 33906 12962
rect 35534 12910 35586 12962
rect 40798 12910 40850 12962
rect 41134 12910 41186 12962
rect 41918 12910 41970 12962
rect 45166 12910 45218 12962
rect 45950 12910 46002 12962
rect 2606 12798 2658 12850
rect 3838 12798 3890 12850
rect 4846 12798 4898 12850
rect 8766 12798 8818 12850
rect 15934 12798 15986 12850
rect 16494 12798 16546 12850
rect 17726 12798 17778 12850
rect 25454 12798 25506 12850
rect 26126 12798 26178 12850
rect 27694 12798 27746 12850
rect 31726 12798 31778 12850
rect 34190 12798 34242 12850
rect 34414 12798 34466 12850
rect 35870 12798 35922 12850
rect 37326 12798 37378 12850
rect 40126 12798 40178 12850
rect 2270 12686 2322 12738
rect 7646 12686 7698 12738
rect 12126 12686 12178 12738
rect 12350 12686 12402 12738
rect 16158 12686 16210 12738
rect 16270 12686 16322 12738
rect 16718 12686 16770 12738
rect 17614 12686 17666 12738
rect 22094 12686 22146 12738
rect 23886 12686 23938 12738
rect 24222 12686 24274 12738
rect 25902 12686 25954 12738
rect 26238 12686 26290 12738
rect 27806 12686 27858 12738
rect 28366 12686 28418 12738
rect 32622 12686 32674 12738
rect 37662 12686 37714 12738
rect 44942 12686 44994 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4734 12350 4786 12402
rect 5294 12350 5346 12402
rect 5742 12350 5794 12402
rect 13134 12350 13186 12402
rect 15934 12350 15986 12402
rect 17726 12350 17778 12402
rect 18510 12350 18562 12402
rect 22542 12350 22594 12402
rect 25454 12350 25506 12402
rect 26238 12350 26290 12402
rect 30494 12350 30546 12402
rect 35422 12350 35474 12402
rect 38670 12350 38722 12402
rect 39230 12350 39282 12402
rect 42254 12350 42306 12402
rect 46286 12350 46338 12402
rect 7870 12238 7922 12290
rect 8206 12238 8258 12290
rect 14590 12238 14642 12290
rect 16270 12238 16322 12290
rect 17614 12238 17666 12290
rect 18622 12238 18674 12290
rect 21086 12238 21138 12290
rect 21422 12238 21474 12290
rect 21982 12238 22034 12290
rect 22318 12238 22370 12290
rect 27582 12238 27634 12290
rect 28142 12238 28194 12290
rect 31502 12238 31554 12290
rect 32286 12238 32338 12290
rect 44158 12238 44210 12290
rect 46622 12238 46674 12290
rect 1710 12126 1762 12178
rect 2270 12126 2322 12178
rect 14366 12126 14418 12178
rect 15038 12126 15090 12178
rect 17950 12126 18002 12178
rect 20862 12126 20914 12178
rect 21758 12126 21810 12178
rect 22654 12126 22706 12178
rect 23102 12126 23154 12178
rect 25902 12126 25954 12178
rect 26574 12126 26626 12178
rect 27694 12126 27746 12178
rect 29150 12126 29202 12178
rect 29934 12126 29986 12178
rect 30270 12126 30322 12178
rect 30718 12126 30770 12178
rect 31054 12126 31106 12178
rect 32510 12126 32562 12178
rect 33070 12126 33122 12178
rect 33518 12126 33570 12178
rect 34302 12126 34354 12178
rect 34526 12126 34578 12178
rect 34862 12126 34914 12178
rect 35758 12126 35810 12178
rect 36094 12126 36146 12178
rect 37438 12126 37490 12178
rect 37998 12126 38050 12178
rect 42590 12126 42642 12178
rect 43262 12126 43314 12178
rect 44382 12126 44434 12178
rect 14478 12014 14530 12066
rect 15598 12014 15650 12066
rect 21870 12014 21922 12066
rect 23550 12014 23602 12066
rect 27022 12014 27074 12066
rect 30494 12014 30546 12066
rect 32622 12014 32674 12066
rect 38110 12014 38162 12066
rect 38446 12014 38498 12066
rect 38782 12014 38834 12066
rect 41022 12014 41074 12066
rect 43598 12014 43650 12066
rect 18398 11902 18450 11954
rect 22878 11902 22930 11954
rect 28590 11902 28642 11954
rect 29822 11902 29874 11954
rect 36094 11902 36146 11954
rect 36430 11902 36482 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 14926 11566 14978 11618
rect 15374 11566 15426 11618
rect 19182 11566 19234 11618
rect 22878 11566 22930 11618
rect 47406 11566 47458 11618
rect 11006 11454 11058 11506
rect 11454 11454 11506 11506
rect 13918 11454 13970 11506
rect 14702 11454 14754 11506
rect 16046 11454 16098 11506
rect 17614 11454 17666 11506
rect 18398 11454 18450 11506
rect 18958 11454 19010 11506
rect 26462 11454 26514 11506
rect 27022 11454 27074 11506
rect 27806 11454 27858 11506
rect 29934 11454 29986 11506
rect 32174 11454 32226 11506
rect 35422 11454 35474 11506
rect 39006 11454 39058 11506
rect 7870 11342 7922 11394
rect 8542 11342 8594 11394
rect 12910 11342 12962 11394
rect 14254 11342 14306 11394
rect 14478 11342 14530 11394
rect 15934 11342 15986 11394
rect 17838 11342 17890 11394
rect 20302 11342 20354 11394
rect 20526 11342 20578 11394
rect 20862 11342 20914 11394
rect 21422 11342 21474 11394
rect 21534 11342 21586 11394
rect 22094 11342 22146 11394
rect 22654 11342 22706 11394
rect 23102 11342 23154 11394
rect 23662 11342 23714 11394
rect 28478 11342 28530 11394
rect 29598 11342 29650 11394
rect 30606 11342 30658 11394
rect 31614 11342 31666 11394
rect 32622 11342 32674 11394
rect 35086 11342 35138 11394
rect 35534 11342 35586 11394
rect 36990 11342 37042 11394
rect 37214 11342 37266 11394
rect 38110 11342 38162 11394
rect 41918 11342 41970 11394
rect 46958 11342 47010 11394
rect 12350 11230 12402 11282
rect 21646 11230 21698 11282
rect 23214 11230 23266 11282
rect 24334 11230 24386 11282
rect 29374 11230 29426 11282
rect 30382 11230 30434 11282
rect 31838 11230 31890 11282
rect 32510 11230 32562 11282
rect 34526 11230 34578 11282
rect 36206 11230 36258 11282
rect 37774 11230 37826 11282
rect 38222 11230 38274 11282
rect 41134 11230 41186 11282
rect 46622 11230 46674 11282
rect 4958 11118 5010 11170
rect 15710 11118 15762 11170
rect 16158 11118 16210 11170
rect 19518 11118 19570 11170
rect 20750 11118 20802 11170
rect 38446 11118 38498 11170
rect 42366 11118 42418 11170
rect 45502 11118 45554 11170
rect 47742 11118 47794 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4734 10782 4786 10834
rect 8206 10782 8258 10834
rect 15150 10782 15202 10834
rect 15262 10782 15314 10834
rect 15374 10782 15426 10834
rect 18062 10782 18114 10834
rect 18958 10782 19010 10834
rect 19070 10782 19122 10834
rect 21198 10782 21250 10834
rect 22318 10782 22370 10834
rect 22542 10782 22594 10834
rect 22990 10782 23042 10834
rect 27022 10782 27074 10834
rect 33294 10782 33346 10834
rect 38110 10782 38162 10834
rect 39454 10782 39506 10834
rect 45278 10782 45330 10834
rect 14030 10670 14082 10722
rect 19966 10670 20018 10722
rect 20078 10670 20130 10722
rect 20414 10670 20466 10722
rect 31838 10670 31890 10722
rect 33182 10670 33234 10722
rect 35646 10670 35698 10722
rect 37326 10670 37378 10722
rect 37550 10670 37602 10722
rect 38558 10670 38610 10722
rect 38670 10670 38722 10722
rect 38782 10670 38834 10722
rect 39678 10670 39730 10722
rect 45726 10670 45778 10722
rect 46286 10670 46338 10722
rect 47294 10670 47346 10722
rect 47630 10670 47682 10722
rect 1710 10558 1762 10610
rect 2270 10558 2322 10610
rect 5182 10558 5234 10610
rect 5854 10558 5906 10610
rect 8654 10558 8706 10610
rect 9662 10558 9714 10610
rect 13918 10558 13970 10610
rect 14814 10558 14866 10610
rect 17838 10558 17890 10610
rect 19294 10558 19346 10610
rect 19630 10558 19682 10610
rect 19742 10558 19794 10610
rect 20750 10558 20802 10610
rect 21086 10558 21138 10610
rect 21422 10558 21474 10610
rect 21870 10558 21922 10610
rect 23214 10558 23266 10610
rect 27358 10558 27410 10610
rect 27694 10558 27746 10610
rect 28030 10558 28082 10610
rect 29486 10558 29538 10610
rect 30718 10558 30770 10610
rect 31054 10558 31106 10610
rect 34638 10558 34690 10610
rect 35198 10558 35250 10610
rect 37774 10558 37826 10610
rect 37886 10558 37938 10610
rect 39790 10558 39842 10610
rect 42142 10558 42194 10610
rect 42926 10558 42978 10610
rect 46510 10558 46562 10610
rect 10334 10446 10386 10498
rect 12462 10446 12514 10498
rect 14366 10446 14418 10498
rect 14702 10446 14754 10498
rect 15822 10446 15874 10498
rect 22430 10446 22482 10498
rect 22878 10446 22930 10498
rect 31950 10446 32002 10498
rect 12910 10334 12962 10386
rect 13246 10334 13298 10386
rect 20750 10334 20802 10386
rect 39230 10334 39282 10386
rect 46846 10334 46898 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 3838 9998 3890 10050
rect 7982 9998 8034 10050
rect 12350 9998 12402 10050
rect 12574 9998 12626 10050
rect 14030 9998 14082 10050
rect 14366 9998 14418 10050
rect 22430 9998 22482 10050
rect 29150 9998 29202 10050
rect 29486 9998 29538 10050
rect 33630 9998 33682 10050
rect 33854 9998 33906 10050
rect 12686 9886 12738 9938
rect 22654 9886 22706 9938
rect 24894 9886 24946 9938
rect 27022 9886 27074 9938
rect 29710 9886 29762 9938
rect 35086 9886 35138 9938
rect 35870 9886 35922 9938
rect 37998 9886 38050 9938
rect 39118 9886 39170 9938
rect 44942 9886 44994 9938
rect 48302 9886 48354 9938
rect 4510 9774 4562 9826
rect 10894 9774 10946 9826
rect 13582 9774 13634 9826
rect 21310 9774 21362 9826
rect 21534 9774 21586 9826
rect 21982 9774 22034 9826
rect 24110 9774 24162 9826
rect 27918 9774 27970 9826
rect 31054 9774 31106 9826
rect 31390 9774 31442 9826
rect 32398 9774 32450 9826
rect 33070 9774 33122 9826
rect 33182 9774 33234 9826
rect 33406 9774 33458 9826
rect 35534 9774 35586 9826
rect 37102 9774 37154 9826
rect 37662 9774 37714 9826
rect 42030 9774 42082 9826
rect 43486 9774 43538 9826
rect 45166 9774 45218 9826
rect 45950 9774 46002 9826
rect 2158 9662 2210 9714
rect 2494 9662 2546 9714
rect 3502 9662 3554 9714
rect 4622 9662 4674 9714
rect 6078 9662 6130 9714
rect 6414 9662 6466 9714
rect 7646 9662 7698 9714
rect 8318 9662 8370 9714
rect 8542 9662 8594 9714
rect 10558 9662 10610 9714
rect 14142 9662 14194 9714
rect 15486 9662 15538 9714
rect 16606 9662 16658 9714
rect 17166 9662 17218 9714
rect 17502 9662 17554 9714
rect 18398 9662 18450 9714
rect 19294 9662 19346 9714
rect 21758 9662 21810 9714
rect 30382 9662 30434 9714
rect 31950 9662 32002 9714
rect 32846 9662 32898 9714
rect 33966 9662 34018 9714
rect 36094 9662 36146 9714
rect 37214 9662 37266 9714
rect 41246 9662 41298 9714
rect 43150 9662 43202 9714
rect 9438 9550 9490 9602
rect 11902 9550 11954 9602
rect 12350 9550 12402 9602
rect 14926 9550 14978 9602
rect 15262 9550 15314 9602
rect 15374 9550 15426 9602
rect 16046 9550 16098 9602
rect 16718 9550 16770 9602
rect 16942 9550 16994 9602
rect 18062 9550 18114 9602
rect 18286 9550 18338 9602
rect 18846 9550 18898 9602
rect 19406 9550 19458 9602
rect 19854 9550 19906 9602
rect 20638 9550 20690 9602
rect 21646 9550 21698 9602
rect 22654 9550 22706 9602
rect 23774 9550 23826 9602
rect 28142 9550 28194 9602
rect 28590 9550 28642 9602
rect 31502 9550 31554 9602
rect 32622 9550 32674 9602
rect 34302 9550 34354 9602
rect 34638 9550 34690 9602
rect 37438 9550 37490 9602
rect 37886 9550 37938 9602
rect 38110 9550 38162 9602
rect 38334 9550 38386 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 11006 9214 11058 9266
rect 11342 9214 11394 9266
rect 14478 9214 14530 9266
rect 14702 9214 14754 9266
rect 17614 9214 17666 9266
rect 19070 9214 19122 9266
rect 19294 9214 19346 9266
rect 19406 9214 19458 9266
rect 34302 9214 34354 9266
rect 34862 9214 34914 9266
rect 39454 9214 39506 9266
rect 4398 9102 4450 9154
rect 6302 9102 6354 9154
rect 8430 9102 8482 9154
rect 15038 9102 15090 9154
rect 17838 9102 17890 9154
rect 18174 9102 18226 9154
rect 19854 9102 19906 9154
rect 21534 9102 21586 9154
rect 21646 9102 21698 9154
rect 24670 9102 24722 9154
rect 25230 9102 25282 9154
rect 25678 9102 25730 9154
rect 32174 9102 32226 9154
rect 33630 9102 33682 9154
rect 37550 9102 37602 9154
rect 45950 9102 46002 9154
rect 3726 8990 3778 9042
rect 4510 8990 4562 9042
rect 6638 8990 6690 9042
rect 7422 8990 7474 9042
rect 7758 8990 7810 9042
rect 8318 8990 8370 9042
rect 12574 8990 12626 9042
rect 16158 8990 16210 9042
rect 17278 8990 17330 9042
rect 18510 8990 18562 9042
rect 18846 8990 18898 9042
rect 19182 8990 19234 9042
rect 20190 8990 20242 9042
rect 21198 8990 21250 9042
rect 22990 8990 23042 9042
rect 23326 8990 23378 9042
rect 25454 8990 25506 9042
rect 27582 8990 27634 9042
rect 27918 8990 27970 9042
rect 28478 8990 28530 9042
rect 28814 8990 28866 9042
rect 29150 8990 29202 9042
rect 32286 8990 32338 9042
rect 33406 8990 33458 9042
rect 34078 8990 34130 9042
rect 38334 8990 38386 9042
rect 39230 8990 39282 9042
rect 46286 8990 46338 9042
rect 5070 8878 5122 8930
rect 9662 8878 9714 8930
rect 11902 8878 11954 8930
rect 12126 8878 12178 8930
rect 12462 8878 12514 8930
rect 13694 8878 13746 8930
rect 15374 8878 15426 8930
rect 16494 8878 16546 8930
rect 16830 8878 16882 8930
rect 17502 8878 17554 8930
rect 20302 8878 20354 8930
rect 22206 8878 22258 8930
rect 27134 8878 27186 8930
rect 31054 8878 31106 8930
rect 33070 8878 33122 8930
rect 35422 8878 35474 8930
rect 38782 8878 38834 8930
rect 3390 8766 3442 8818
rect 15486 8766 15538 8818
rect 21646 8766 21698 8818
rect 23326 8766 23378 8818
rect 25790 8766 25842 8818
rect 34414 8766 34466 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 16158 8430 16210 8482
rect 16494 8430 16546 8482
rect 37326 8430 37378 8482
rect 4734 8318 4786 8370
rect 8654 8318 8706 8370
rect 11902 8318 11954 8370
rect 13694 8318 13746 8370
rect 14590 8318 14642 8370
rect 17390 8318 17442 8370
rect 18734 8318 18786 8370
rect 24222 8318 24274 8370
rect 25678 8318 25730 8370
rect 27918 8318 27970 8370
rect 28478 8318 28530 8370
rect 29486 8318 29538 8370
rect 34078 8318 34130 8370
rect 35198 8318 35250 8370
rect 37214 8318 37266 8370
rect 38558 8318 38610 8370
rect 44942 8318 44994 8370
rect 1710 8206 1762 8258
rect 2270 8206 2322 8258
rect 5742 8206 5794 8258
rect 6302 8206 6354 8258
rect 8990 8206 9042 8258
rect 17726 8206 17778 8258
rect 18846 8206 18898 8258
rect 19294 8206 19346 8258
rect 21310 8206 21362 8258
rect 24894 8206 24946 8258
rect 29262 8206 29314 8258
rect 29822 8206 29874 8258
rect 31838 8206 31890 8258
rect 34750 8206 34802 8258
rect 35758 8206 35810 8258
rect 41582 8206 41634 8258
rect 45166 8206 45218 8258
rect 45950 8206 46002 8258
rect 9774 8094 9826 8146
rect 12574 8094 12626 8146
rect 12798 8094 12850 8146
rect 13582 8094 13634 8146
rect 15262 8094 15314 8146
rect 16382 8094 16434 8146
rect 18174 8094 18226 8146
rect 18510 8094 18562 8146
rect 19630 8094 19682 8146
rect 20190 8094 20242 8146
rect 22094 8094 22146 8146
rect 30382 8094 30434 8146
rect 32398 8094 32450 8146
rect 40574 8094 40626 8146
rect 12686 7982 12738 8034
rect 14030 7982 14082 8034
rect 15598 7982 15650 8034
rect 20526 7982 20578 8034
rect 29934 7982 29986 8034
rect 36206 7982 36258 8034
rect 37886 7982 37938 8034
rect 41358 7982 41410 8034
rect 42478 7982 42530 8034
rect 48302 7982 48354 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 2158 7646 2210 7698
rect 4286 7646 4338 7698
rect 5630 7646 5682 7698
rect 6078 7646 6130 7698
rect 7758 7646 7810 7698
rect 8206 7646 8258 7698
rect 10110 7646 10162 7698
rect 16382 7646 16434 7698
rect 16718 7646 16770 7698
rect 20414 7646 20466 7698
rect 21310 7646 21362 7698
rect 23662 7646 23714 7698
rect 24110 7646 24162 7698
rect 24558 7646 24610 7698
rect 29822 7646 29874 7698
rect 30830 7646 30882 7698
rect 32510 7646 32562 7698
rect 33294 7646 33346 7698
rect 34638 7646 34690 7698
rect 34974 7646 35026 7698
rect 35534 7646 35586 7698
rect 35870 7646 35922 7698
rect 36654 7646 36706 7698
rect 38110 7646 38162 7698
rect 41246 7646 41298 7698
rect 43822 7646 43874 7698
rect 46510 7646 46562 7698
rect 2494 7534 2546 7586
rect 11230 7534 11282 7586
rect 11342 7534 11394 7586
rect 12798 7534 12850 7586
rect 13582 7534 13634 7586
rect 15598 7534 15650 7586
rect 17950 7534 18002 7586
rect 20638 7534 20690 7586
rect 20974 7534 21026 7586
rect 21982 7534 22034 7586
rect 28142 7534 28194 7586
rect 29262 7534 29314 7586
rect 29710 7534 29762 7586
rect 32174 7534 32226 7586
rect 34078 7534 34130 7586
rect 42366 7534 42418 7586
rect 44270 7534 44322 7586
rect 47182 7534 47234 7586
rect 47630 7534 47682 7586
rect 10446 7422 10498 7474
rect 11006 7422 11058 7474
rect 11790 7422 11842 7474
rect 12126 7422 12178 7474
rect 12910 7422 12962 7474
rect 13918 7422 13970 7474
rect 18174 7422 18226 7474
rect 18510 7422 18562 7474
rect 18846 7422 18898 7474
rect 19182 7422 19234 7474
rect 25678 7422 25730 7474
rect 26462 7422 26514 7474
rect 26910 7422 26962 7474
rect 27470 7422 27522 7474
rect 27694 7422 27746 7474
rect 28366 7422 28418 7474
rect 29038 7422 29090 7474
rect 30718 7422 30770 7474
rect 30942 7422 30994 7474
rect 31502 7422 31554 7474
rect 37550 7422 37602 7474
rect 37886 7422 37938 7474
rect 38782 7422 38834 7474
rect 39342 7422 39394 7474
rect 40238 7422 40290 7474
rect 42030 7422 42082 7474
rect 43150 7422 43202 7474
rect 43598 7422 43650 7474
rect 45054 7422 45106 7474
rect 45950 7422 46002 7474
rect 4734 7310 4786 7362
rect 5070 7310 5122 7362
rect 6526 7310 6578 7362
rect 7198 7310 7250 7362
rect 8542 7310 8594 7362
rect 9102 7310 9154 7362
rect 9774 7310 9826 7362
rect 14590 7310 14642 7362
rect 18398 7310 18450 7362
rect 19742 7310 19794 7362
rect 20414 7310 20466 7362
rect 22990 7310 23042 7362
rect 25902 7310 25954 7362
rect 27918 7310 27970 7362
rect 33630 7310 33682 7362
rect 37102 7310 37154 7362
rect 42814 7310 42866 7362
rect 48190 7310 48242 7362
rect 7870 7198 7922 7250
rect 8430 7198 8482 7250
rect 17390 7198 17442 7250
rect 17726 7198 17778 7250
rect 25566 7198 25618 7250
rect 41582 7198 41634 7250
rect 46846 7198 46898 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 3950 6862 4002 6914
rect 7870 6862 7922 6914
rect 12574 6862 12626 6914
rect 15150 6862 15202 6914
rect 15486 6862 15538 6914
rect 18286 6862 18338 6914
rect 35534 6862 35586 6914
rect 46958 6862 47010 6914
rect 6078 6750 6130 6802
rect 15598 6750 15650 6802
rect 16158 6750 16210 6802
rect 18958 6750 19010 6802
rect 23998 6750 24050 6802
rect 29822 6750 29874 6802
rect 31278 6750 31330 6802
rect 34750 6750 34802 6802
rect 4734 6638 4786 6690
rect 9886 6638 9938 6690
rect 10670 6638 10722 6690
rect 11006 6638 11058 6690
rect 12798 6638 12850 6690
rect 13918 6638 13970 6690
rect 15262 6638 15314 6690
rect 18062 6638 18114 6690
rect 18622 6638 18674 6690
rect 21534 6638 21586 6690
rect 22206 6638 22258 6690
rect 23214 6638 23266 6690
rect 26014 6638 26066 6690
rect 28142 6638 28194 6690
rect 28366 6638 28418 6690
rect 29150 6638 29202 6690
rect 29262 6638 29314 6690
rect 29598 6638 29650 6690
rect 31950 6638 32002 6690
rect 32622 6638 32674 6690
rect 36094 6638 36146 6690
rect 37214 6638 37266 6690
rect 37550 6638 37602 6690
rect 37998 6638 38050 6690
rect 40350 6638 40402 6690
rect 40798 6638 40850 6690
rect 41358 6638 41410 6690
rect 43710 6638 43762 6690
rect 45054 6638 45106 6690
rect 45502 6638 45554 6690
rect 1934 6526 1986 6578
rect 4510 6526 4562 6578
rect 6750 6526 6802 6578
rect 7534 6526 7586 6578
rect 8094 6526 8146 6578
rect 8542 6526 8594 6578
rect 10222 6526 10274 6578
rect 11230 6526 11282 6578
rect 11566 6526 11618 6578
rect 14142 6526 14194 6578
rect 14478 6526 14530 6578
rect 17166 6526 17218 6578
rect 20302 6526 20354 6578
rect 21422 6526 21474 6578
rect 25006 6526 25058 6578
rect 26574 6526 26626 6578
rect 26798 6526 26850 6578
rect 27806 6526 27858 6578
rect 30158 6526 30210 6578
rect 30494 6526 30546 6578
rect 36318 6526 36370 6578
rect 38558 6526 38610 6578
rect 46174 6526 46226 6578
rect 46622 6526 46674 6578
rect 47182 6526 47234 6578
rect 47518 6526 47570 6578
rect 2830 6414 2882 6466
rect 3278 6414 3330 6466
rect 3614 6414 3666 6466
rect 6414 6414 6466 6466
rect 9214 6414 9266 6466
rect 9550 6414 9602 6466
rect 12238 6414 12290 6466
rect 13582 6414 13634 6466
rect 22542 6414 22594 6466
rect 23774 6414 23826 6466
rect 26126 6414 26178 6466
rect 28030 6414 28082 6466
rect 30830 6414 30882 6466
rect 35198 6414 35250 6466
rect 39006 6414 39058 6466
rect 39790 6414 39842 6466
rect 45838 6414 45890 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4734 6078 4786 6130
rect 5182 6078 5234 6130
rect 8654 6078 8706 6130
rect 17726 6078 17778 6130
rect 24222 6078 24274 6130
rect 24446 6078 24498 6130
rect 24670 6078 24722 6130
rect 25342 6078 25394 6130
rect 25566 6078 25618 6130
rect 26350 6078 26402 6130
rect 27246 6078 27298 6130
rect 33742 6078 33794 6130
rect 38222 6078 38274 6130
rect 38670 6078 38722 6130
rect 44942 6078 44994 6130
rect 45390 6078 45442 6130
rect 9774 5966 9826 6018
rect 9998 5966 10050 6018
rect 10670 5966 10722 6018
rect 11790 5966 11842 6018
rect 15038 5966 15090 6018
rect 16382 5966 16434 6018
rect 18398 5966 18450 6018
rect 18734 5966 18786 6018
rect 20526 5966 20578 6018
rect 23550 5966 23602 6018
rect 25230 5966 25282 6018
rect 28254 5966 28306 6018
rect 31726 5966 31778 6018
rect 37438 5966 37490 6018
rect 39678 5966 39730 6018
rect 40238 5966 40290 6018
rect 41470 5966 41522 6018
rect 43150 5966 43202 6018
rect 1710 5854 1762 5906
rect 2270 5854 2322 5906
rect 5742 5854 5794 5906
rect 6302 5854 6354 5906
rect 10446 5854 10498 5906
rect 11006 5854 11058 5906
rect 14814 5854 14866 5906
rect 17390 5854 17442 5906
rect 19742 5854 19794 5906
rect 22990 5854 23042 5906
rect 23214 5854 23266 5906
rect 23438 5854 23490 5906
rect 25790 5854 25842 5906
rect 26910 5854 26962 5906
rect 28366 5854 28418 5906
rect 32510 5854 32562 5906
rect 33518 5854 33570 5906
rect 34078 5854 34130 5906
rect 34638 5854 34690 5906
rect 37662 5854 37714 5906
rect 39454 5854 39506 5906
rect 42926 5854 42978 5906
rect 43710 5854 43762 5906
rect 45726 5854 45778 5906
rect 9662 5742 9714 5794
rect 13918 5742 13970 5794
rect 14366 5742 14418 5794
rect 15374 5742 15426 5794
rect 22654 5742 22706 5794
rect 24558 5742 24610 5794
rect 26014 5742 26066 5794
rect 26686 5742 26738 5794
rect 29598 5742 29650 5794
rect 37102 5742 37154 5794
rect 41022 5742 41074 5794
rect 42142 5742 42194 5794
rect 46846 5742 46898 5794
rect 18958 5630 19010 5682
rect 19294 5630 19346 5682
rect 28814 5630 28866 5682
rect 29150 5630 29202 5682
rect 39118 5630 39170 5682
rect 44046 5630 44098 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 4174 5294 4226 5346
rect 12350 5294 12402 5346
rect 12686 5294 12738 5346
rect 29598 5294 29650 5346
rect 31054 5294 31106 5346
rect 37662 5294 37714 5346
rect 37998 5294 38050 5346
rect 1822 5182 1874 5234
rect 3054 5182 3106 5234
rect 3502 5182 3554 5234
rect 5742 5182 5794 5234
rect 9550 5182 9602 5234
rect 11678 5182 11730 5234
rect 15150 5182 15202 5234
rect 16270 5182 16322 5234
rect 18398 5182 18450 5234
rect 18734 5182 18786 5234
rect 20750 5182 20802 5234
rect 24894 5182 24946 5234
rect 31726 5182 31778 5234
rect 35534 5182 35586 5234
rect 35982 5182 36034 5234
rect 36430 5182 36482 5234
rect 36990 5182 37042 5234
rect 43262 5182 43314 5234
rect 44830 5182 44882 5234
rect 48302 5182 48354 5234
rect 2494 5070 2546 5122
rect 3838 5070 3890 5122
rect 4846 5070 4898 5122
rect 6414 5070 6466 5122
rect 7086 5070 7138 5122
rect 7534 5070 7586 5122
rect 8206 5070 8258 5122
rect 8878 5070 8930 5122
rect 12910 5070 12962 5122
rect 15486 5070 15538 5122
rect 21422 5070 21474 5122
rect 22094 5070 22146 5122
rect 27246 5070 27298 5122
rect 27582 5070 27634 5122
rect 28590 5070 28642 5122
rect 29262 5070 29314 5122
rect 30046 5070 30098 5122
rect 30830 5070 30882 5122
rect 34638 5070 34690 5122
rect 35086 5070 35138 5122
rect 38558 5070 38610 5122
rect 39230 5070 39282 5122
rect 42142 5070 42194 5122
rect 43710 5070 43762 5122
rect 45166 5070 45218 5122
rect 45838 5070 45890 5122
rect 2158 4958 2210 5010
rect 4734 4958 4786 5010
rect 8430 4958 8482 5010
rect 14142 4958 14194 5010
rect 19742 4958 19794 5010
rect 28254 4958 28306 5010
rect 30270 4958 30322 5010
rect 33854 4958 33906 5010
rect 38782 4958 38834 5010
rect 6078 4846 6130 4898
rect 6750 4846 6802 4898
rect 7758 4846 7810 4898
rect 22766 4846 22818 4898
rect 27918 4846 27970 4898
rect 31390 4846 31442 4898
rect 37102 4846 37154 4898
rect 40238 4846 40290 4898
rect 42478 4846 42530 4898
rect 43934 4846 43986 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 4846 4510 4898 4562
rect 5742 4510 5794 4562
rect 18174 4510 18226 4562
rect 20750 4510 20802 4562
rect 34078 4510 34130 4562
rect 39566 4510 39618 4562
rect 40910 4510 40962 4562
rect 47294 4510 47346 4562
rect 6862 4398 6914 4450
rect 10558 4398 10610 4450
rect 13582 4398 13634 4450
rect 14478 4398 14530 4450
rect 17390 4398 17442 4450
rect 17502 4398 17554 4450
rect 17726 4398 17778 4450
rect 18510 4398 18562 4450
rect 19070 4398 19122 4450
rect 21310 4398 21362 4450
rect 22542 4398 22594 4450
rect 25902 4398 25954 4450
rect 26238 4398 26290 4450
rect 33070 4398 33122 4450
rect 33742 4398 33794 4450
rect 34414 4398 34466 4450
rect 34862 4398 34914 4450
rect 35870 4398 35922 4450
rect 40014 4398 40066 4450
rect 40350 4398 40402 4450
rect 1710 4286 1762 4338
rect 2382 4286 2434 4338
rect 5518 4286 5570 4338
rect 6078 4286 6130 4338
rect 10222 4286 10274 4338
rect 11118 4286 11170 4338
rect 17838 4286 17890 4338
rect 18174 4286 18226 4338
rect 21870 4286 21922 4338
rect 26910 4286 26962 4338
rect 31950 4286 32002 4338
rect 33294 4286 33346 4338
rect 36430 4286 36482 4338
rect 37214 4286 37266 4338
rect 43262 4286 43314 4338
rect 43822 4286 43874 4338
rect 44158 4286 44210 4338
rect 44830 4286 44882 4338
rect 8990 4174 9042 4226
rect 10670 4174 10722 4226
rect 16606 4174 16658 4226
rect 20190 4174 20242 4226
rect 24670 4174 24722 4226
rect 25678 4174 25730 4226
rect 11454 4062 11506 4114
rect 25342 4062 25394 4114
rect 27918 4062 27970 4114
rect 30046 4062 30098 4114
rect 35310 4062 35362 4114
rect 35758 4062 35810 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 16830 3726 16882 3778
rect 20750 3726 20802 3778
rect 21086 3726 21138 3778
rect 24558 3726 24610 3778
rect 24894 3726 24946 3778
rect 8206 3614 8258 3666
rect 9326 3614 9378 3666
rect 11118 3614 11170 3666
rect 13470 3614 13522 3666
rect 29374 3614 29426 3666
rect 36990 3614 37042 3666
rect 40798 3614 40850 3666
rect 44606 3614 44658 3666
rect 46510 3614 46562 3666
rect 48190 3614 48242 3666
rect 1822 3502 1874 3554
rect 2494 3502 2546 3554
rect 3166 3502 3218 3554
rect 3726 3502 3778 3554
rect 4398 3502 4450 3554
rect 5966 3502 6018 3554
rect 6078 3502 6130 3554
rect 6974 3502 7026 3554
rect 7646 3502 7698 3554
rect 8766 3502 8818 3554
rect 19966 3502 20018 3554
rect 21422 3502 21474 3554
rect 25230 3502 25282 3554
rect 28366 3502 28418 3554
rect 31278 3502 31330 3554
rect 32622 3502 32674 3554
rect 35198 3502 35250 3554
rect 36430 3502 36482 3554
rect 39790 3502 39842 3554
rect 43598 3502 43650 3554
rect 2718 3390 2770 3442
rect 3390 3390 3442 3442
rect 4062 3390 4114 3442
rect 4958 3390 5010 3442
rect 5518 3390 5570 3442
rect 6190 3390 6242 3442
rect 7198 3390 7250 3442
rect 7870 3390 7922 3442
rect 10670 3390 10722 3442
rect 12462 3390 12514 3442
rect 13582 3390 13634 3442
rect 15710 3390 15762 3442
rect 19294 3390 19346 3442
rect 20190 3390 20242 3442
rect 20974 3390 21026 3442
rect 23214 3390 23266 3442
rect 24782 3390 24834 3442
rect 31614 3390 31666 3442
rect 33742 3390 33794 3442
rect 2046 3278 2098 3330
rect 26238 3278 26290 3330
rect 35422 3278 35474 3330
rect 38894 3278 38946 3330
rect 42702 3278 42754 3330
rect 47406 3278 47458 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 27020 50370 27076 50382
rect 27020 50318 27022 50370
rect 27074 50318 27076 50370
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 27020 50034 27076 50318
rect 27020 49982 27022 50034
rect 27074 49982 27076 50034
rect 27020 49970 27076 49982
rect 27916 50370 27972 50382
rect 27916 50318 27918 50370
rect 27970 50318 27972 50370
rect 26796 49812 26852 49822
rect 26796 49810 27412 49812
rect 26796 49758 26798 49810
rect 26850 49758 27412 49810
rect 26796 49756 27412 49758
rect 26796 49746 26852 49756
rect 21084 49700 21140 49710
rect 21532 49700 21588 49710
rect 21084 49698 21588 49700
rect 21084 49646 21086 49698
rect 21138 49646 21534 49698
rect 21586 49646 21588 49698
rect 21084 49644 21588 49646
rect 21084 49634 21140 49644
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 14476 49028 14532 49038
rect 14476 48934 14532 48972
rect 15036 49026 15092 49038
rect 15036 48974 15038 49026
rect 15090 48974 15092 49026
rect 15036 48804 15092 48974
rect 16828 49028 16884 49038
rect 15036 48738 15092 48748
rect 16268 48804 16324 48814
rect 16268 48466 16324 48748
rect 16268 48414 16270 48466
rect 16322 48414 16324 48466
rect 16268 48402 16324 48414
rect 16604 48244 16660 48254
rect 16604 48150 16660 48188
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 9996 47458 10052 47470
rect 9996 47406 9998 47458
rect 10050 47406 10052 47458
rect 9996 46900 10052 47406
rect 10556 47460 10612 47470
rect 10556 47458 10948 47460
rect 10556 47406 10558 47458
rect 10610 47406 10948 47458
rect 10556 47404 10948 47406
rect 10556 47394 10612 47404
rect 9996 46834 10052 46844
rect 10892 46898 10948 47404
rect 12908 47236 12964 47246
rect 12796 47234 12964 47236
rect 12796 47182 12910 47234
rect 12962 47182 12964 47234
rect 12796 47180 12964 47182
rect 10892 46846 10894 46898
rect 10946 46846 10948 46898
rect 10892 46834 10948 46846
rect 11004 46900 11060 46910
rect 9548 46788 9604 46798
rect 8876 46786 9604 46788
rect 8876 46734 9550 46786
rect 9602 46734 9604 46786
rect 8876 46732 9604 46734
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 8316 45890 8372 45902
rect 8316 45838 8318 45890
rect 8370 45838 8372 45890
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 7532 44322 7588 44334
rect 7532 44270 7534 44322
rect 7586 44270 7588 44322
rect 4732 43540 4788 43550
rect 5292 43540 5348 43550
rect 4732 43538 4900 43540
rect 4732 43486 4734 43538
rect 4786 43486 4900 43538
rect 4732 43484 4900 43486
rect 4732 43474 4788 43484
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 2380 40402 2436 40414
rect 2380 40350 2382 40402
rect 2434 40350 2436 40402
rect 2380 39396 2436 40350
rect 3164 40404 3220 40414
rect 4844 40404 4900 43484
rect 5292 43538 5684 43540
rect 5292 43486 5294 43538
rect 5346 43486 5684 43538
rect 5292 43484 5684 43486
rect 5292 43474 5348 43484
rect 5628 42642 5684 43484
rect 7532 43428 7588 44270
rect 8092 44322 8148 44334
rect 8092 44270 8094 44322
rect 8146 44270 8148 44322
rect 8092 43762 8148 44270
rect 8092 43710 8094 43762
rect 8146 43710 8148 43762
rect 8092 43698 8148 43710
rect 7532 43362 7588 43372
rect 7644 43426 7700 43438
rect 7644 43374 7646 43426
rect 7698 43374 7700 43426
rect 7644 42756 7700 43374
rect 8316 43428 8372 45838
rect 8876 45890 8932 46732
rect 9548 46722 9604 46732
rect 9884 46676 9940 46686
rect 9884 46674 10052 46676
rect 9884 46622 9886 46674
rect 9938 46622 10052 46674
rect 9884 46620 10052 46622
rect 9884 46610 9940 46620
rect 8876 45838 8878 45890
rect 8930 45838 8932 45890
rect 8876 45826 8932 45838
rect 9996 45332 10052 46620
rect 11004 45780 11060 46844
rect 11676 46900 11732 46910
rect 11676 46806 11732 46844
rect 11228 46676 11284 46686
rect 11228 46674 11732 46676
rect 11228 46622 11230 46674
rect 11282 46622 11732 46674
rect 11228 46620 11732 46622
rect 11228 46610 11284 46620
rect 11676 46114 11732 46620
rect 11676 46062 11678 46114
rect 11730 46062 11732 46114
rect 11676 46050 11732 46062
rect 12012 45890 12068 45902
rect 12012 45838 12014 45890
rect 12066 45838 12068 45890
rect 10892 45724 11060 45780
rect 11116 45780 11172 45790
rect 10220 45332 10276 45342
rect 9996 45330 10276 45332
rect 9996 45278 10222 45330
rect 10274 45278 10276 45330
rect 9996 45276 10276 45278
rect 10220 45266 10276 45276
rect 10556 44882 10612 44894
rect 10556 44830 10558 44882
rect 10610 44830 10612 44882
rect 10444 44436 10500 44446
rect 10556 44436 10612 44830
rect 10444 44434 10612 44436
rect 10444 44382 10446 44434
rect 10498 44382 10612 44434
rect 10444 44380 10612 44382
rect 10892 44434 10948 45724
rect 11116 45106 11172 45724
rect 11676 45780 11732 45790
rect 11228 45668 11284 45678
rect 11228 45220 11284 45612
rect 11340 45220 11396 45230
rect 11228 45218 11396 45220
rect 11228 45166 11342 45218
rect 11394 45166 11396 45218
rect 11228 45164 11396 45166
rect 11116 45054 11118 45106
rect 11170 45054 11172 45106
rect 11116 45042 11172 45054
rect 10892 44382 10894 44434
rect 10946 44382 10948 44434
rect 8428 43540 8484 43550
rect 8428 43538 8708 43540
rect 8428 43486 8430 43538
rect 8482 43486 8708 43538
rect 8428 43484 8708 43486
rect 8428 43474 8484 43484
rect 8316 43362 8372 43372
rect 8652 42978 8708 43484
rect 8876 43428 8932 43438
rect 8876 43334 8932 43372
rect 8652 42926 8654 42978
rect 8706 42926 8708 42978
rect 8652 42914 8708 42926
rect 5628 42590 5630 42642
rect 5682 42590 5684 42642
rect 5628 42578 5684 42590
rect 5964 42644 6020 42654
rect 5964 42642 6580 42644
rect 5964 42590 5966 42642
rect 6018 42590 6580 42642
rect 5964 42588 6580 42590
rect 5964 42578 6020 42588
rect 6524 42194 6580 42588
rect 6524 42142 6526 42194
rect 6578 42142 6580 42194
rect 6524 42130 6580 42142
rect 7644 42082 7700 42700
rect 8988 42756 9044 42766
rect 8988 42662 9044 42700
rect 9772 42754 9828 42766
rect 9772 42702 9774 42754
rect 9826 42702 9828 42754
rect 9660 42642 9716 42654
rect 9660 42590 9662 42642
rect 9714 42590 9716 42642
rect 9660 42196 9716 42590
rect 9660 42130 9716 42140
rect 9772 42644 9828 42702
rect 7644 42030 7646 42082
rect 7698 42030 7700 42082
rect 7644 42018 7700 42030
rect 9772 42084 9828 42588
rect 10220 42756 10276 42766
rect 9772 42018 9828 42028
rect 9884 42308 9940 42318
rect 7532 41972 7588 41982
rect 6860 41748 6916 41758
rect 6860 41654 6916 41692
rect 6636 41186 6692 41198
rect 6636 41134 6638 41186
rect 6690 41134 6692 41186
rect 6412 40964 6468 40974
rect 6412 40962 6580 40964
rect 6412 40910 6414 40962
rect 6466 40910 6580 40962
rect 6412 40908 6580 40910
rect 6412 40898 6468 40908
rect 3164 40402 3332 40404
rect 3164 40350 3166 40402
rect 3218 40350 3332 40402
rect 3164 40348 3332 40350
rect 3164 40338 3220 40348
rect 3276 39506 3332 40348
rect 4844 40338 4900 40348
rect 5516 40402 5572 40414
rect 5516 40350 5518 40402
rect 5570 40350 5572 40402
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 3276 39454 3278 39506
rect 3330 39454 3332 39506
rect 3276 39442 3332 39454
rect 3612 39508 3668 39518
rect 3612 39506 3892 39508
rect 3612 39454 3614 39506
rect 3666 39454 3892 39506
rect 3612 39452 3892 39454
rect 3612 39442 3668 39452
rect 2156 39340 2436 39396
rect 1820 38836 1876 38846
rect 2156 38836 2212 39340
rect 1820 38834 2156 38836
rect 1820 38782 1822 38834
rect 1874 38782 2156 38834
rect 1820 38780 2156 38782
rect 1820 37266 1876 38780
rect 2156 38742 2212 38780
rect 2268 38834 2324 38846
rect 2268 38782 2270 38834
rect 2322 38782 2324 38834
rect 2268 37938 2324 38782
rect 3836 38274 3892 39452
rect 5180 38836 5236 38846
rect 4732 38722 4788 38734
rect 4732 38670 4734 38722
rect 4786 38670 4788 38722
rect 4732 38668 4788 38670
rect 4732 38612 4900 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4844 38276 4900 38612
rect 3836 38222 3838 38274
rect 3890 38222 3892 38274
rect 3836 38210 3892 38222
rect 4732 38220 4900 38276
rect 4172 38050 4228 38062
rect 4172 37998 4174 38050
rect 4226 37998 4228 38050
rect 2268 37886 2270 37938
rect 2322 37886 2324 37938
rect 2268 37874 2324 37886
rect 2604 37940 2660 37950
rect 2604 37846 2660 37884
rect 1820 37214 1822 37266
rect 1874 37214 1876 37266
rect 1820 37202 1876 37214
rect 2380 37268 2436 37278
rect 2380 37266 2548 37268
rect 2380 37214 2382 37266
rect 2434 37214 2548 37266
rect 2380 37212 2548 37214
rect 2380 37202 2436 37212
rect 2492 36370 2548 37212
rect 4172 37156 4228 37998
rect 4172 37090 4228 37100
rect 4284 37492 4340 37502
rect 2492 36318 2494 36370
rect 2546 36318 2548 36370
rect 2492 36306 2548 36318
rect 2828 36372 2884 36382
rect 2828 36278 2884 36316
rect 1820 34914 1876 34926
rect 1820 34862 1822 34914
rect 1874 34862 1876 34914
rect 1820 32562 1876 34862
rect 2380 34914 2436 34926
rect 2380 34862 2382 34914
rect 2434 34862 2436 34914
rect 2380 34354 2436 34862
rect 2380 34302 2382 34354
rect 2434 34302 2436 34354
rect 2380 34290 2436 34302
rect 3836 34916 3892 34926
rect 2716 34132 2772 34142
rect 2716 34038 2772 34076
rect 3836 33570 3892 34860
rect 4172 34132 4228 34142
rect 4284 34132 4340 37436
rect 4732 37492 4788 38220
rect 4956 38164 5012 38174
rect 4844 38052 4900 38062
rect 4844 37958 4900 37996
rect 4956 37938 5012 38108
rect 4956 37886 4958 37938
rect 5010 37886 5012 37938
rect 4956 37874 5012 37886
rect 4732 37426 4788 37436
rect 5180 37490 5236 38780
rect 5516 38164 5572 40350
rect 5740 40404 5796 40414
rect 5852 40404 5908 40414
rect 5796 40402 5908 40404
rect 5796 40350 5854 40402
rect 5906 40350 5908 40402
rect 5796 40348 5908 40350
rect 5740 39732 5796 40348
rect 5852 40338 5908 40348
rect 6524 40402 6580 40908
rect 6524 40350 6526 40402
rect 6578 40350 6580 40402
rect 6524 40338 6580 40350
rect 6636 39844 6692 41134
rect 6748 39844 6804 39854
rect 6636 39842 6804 39844
rect 6636 39790 6750 39842
rect 6802 39790 6804 39842
rect 6636 39788 6804 39790
rect 6748 39778 6804 39788
rect 7084 39844 7140 39854
rect 7084 39750 7140 39788
rect 5740 39394 5796 39676
rect 7532 39618 7588 41916
rect 9660 41970 9716 41982
rect 9660 41918 9662 41970
rect 9714 41918 9716 41970
rect 7532 39566 7534 39618
rect 7586 39566 7588 39618
rect 7532 39554 7588 39566
rect 7644 41748 7700 41758
rect 7644 40404 7700 41692
rect 9324 41186 9380 41198
rect 9324 41134 9326 41186
rect 9378 41134 9380 41186
rect 8988 40516 9044 40526
rect 8988 40422 9044 40460
rect 7644 39506 7700 40348
rect 9212 40180 9268 40190
rect 7644 39454 7646 39506
rect 7698 39454 7700 39506
rect 7644 39442 7700 39454
rect 8988 40124 9212 40180
rect 5740 39342 5742 39394
rect 5794 39342 5796 39394
rect 5740 38836 5796 39342
rect 8988 39058 9044 40124
rect 9212 40114 9268 40124
rect 9324 39732 9380 41134
rect 9660 40626 9716 41918
rect 9660 40574 9662 40626
rect 9714 40574 9716 40626
rect 9660 40562 9716 40574
rect 8988 39006 8990 39058
rect 9042 39006 9044 39058
rect 5852 38836 5908 38846
rect 5796 38834 5908 38836
rect 5796 38782 5854 38834
rect 5906 38782 5908 38834
rect 5796 38780 5908 38782
rect 5740 38770 5796 38780
rect 5852 38770 5908 38780
rect 6636 38834 6692 38846
rect 6636 38782 6638 38834
rect 6690 38782 6692 38834
rect 6636 38276 6692 38782
rect 6636 38210 6692 38220
rect 7420 38276 7476 38286
rect 5516 38098 5572 38108
rect 6076 38164 6132 38174
rect 6076 38070 6132 38108
rect 5180 37438 5182 37490
rect 5234 37438 5236 37490
rect 5180 37426 5236 37438
rect 5292 38052 5348 38062
rect 4732 37156 4788 37166
rect 4732 37062 4788 37100
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4732 34916 4788 34926
rect 4732 34822 4788 34860
rect 5068 34916 5124 34926
rect 5068 34242 5124 34860
rect 5068 34190 5070 34242
rect 5122 34190 5124 34242
rect 5068 34178 5124 34190
rect 5292 34244 5348 37996
rect 6300 38052 6356 38062
rect 5740 37940 5796 37950
rect 5740 37846 5796 37884
rect 6300 37938 6356 37996
rect 6300 37886 6302 37938
rect 6354 37886 6356 37938
rect 6076 36482 6132 36494
rect 6076 36430 6078 36482
rect 6130 36430 6132 36482
rect 5740 36372 5796 36382
rect 5740 36278 5796 36316
rect 4508 34132 4564 34142
rect 4284 34130 4564 34132
rect 4284 34078 4510 34130
rect 4562 34078 4564 34130
rect 4284 34076 4564 34078
rect 4172 34038 4228 34076
rect 4508 34066 4564 34076
rect 5292 34130 5348 34188
rect 5292 34078 5294 34130
rect 5346 34078 5348 34130
rect 5292 34066 5348 34078
rect 5628 35698 5684 35710
rect 5628 35646 5630 35698
rect 5682 35646 5684 35698
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 3836 33518 3838 33570
rect 3890 33518 3892 33570
rect 3836 33506 3892 33518
rect 4396 33346 4452 33358
rect 4396 33294 4398 33346
rect 4450 33294 4452 33346
rect 4396 33236 4452 33294
rect 5628 33348 5684 35646
rect 5740 34244 5796 34254
rect 5740 34150 5796 34188
rect 6076 33572 6132 36430
rect 6300 36370 6356 37886
rect 6860 37938 6916 37950
rect 6860 37886 6862 37938
rect 6914 37886 6916 37938
rect 6860 37492 6916 37886
rect 7420 37938 7476 38220
rect 7420 37886 7422 37938
rect 7474 37886 7476 37938
rect 7420 37874 7476 37886
rect 7756 37940 7812 37950
rect 7756 37938 8260 37940
rect 7756 37886 7758 37938
rect 7810 37886 8260 37938
rect 7756 37884 8260 37886
rect 7756 37874 7812 37884
rect 6860 37426 6916 37436
rect 6300 36318 6302 36370
rect 6354 36318 6356 36370
rect 6300 36306 6356 36318
rect 6860 37156 6916 37166
rect 6860 36370 6916 37100
rect 8204 36706 8260 37884
rect 8204 36654 8206 36706
rect 8258 36654 8260 36706
rect 8204 36642 8260 36654
rect 6860 36318 6862 36370
rect 6914 36318 6916 36370
rect 6860 36306 6916 36318
rect 8540 36482 8596 36494
rect 8540 36430 8542 36482
rect 8594 36430 8596 36482
rect 8540 35924 8596 36430
rect 8540 35830 8596 35868
rect 8764 36370 8820 36382
rect 8764 36318 8766 36370
rect 8818 36318 8820 36370
rect 6188 35700 6244 35710
rect 8428 35700 8484 35710
rect 6188 35698 6468 35700
rect 6188 35646 6190 35698
rect 6242 35646 6468 35698
rect 6188 35644 6468 35646
rect 6188 35634 6244 35644
rect 6412 34802 6468 35644
rect 8316 34914 8372 34926
rect 8316 34862 8318 34914
rect 8370 34862 8372 34914
rect 6412 34750 6414 34802
rect 6466 34750 6468 34802
rect 6412 34738 6468 34750
rect 6748 34804 6804 34814
rect 6748 34710 6804 34748
rect 7980 34804 8036 34814
rect 7980 34710 8036 34748
rect 8316 34692 8372 34862
rect 8316 34626 8372 34636
rect 6076 33506 6132 33516
rect 6188 34130 6244 34142
rect 6188 34078 6190 34130
rect 6242 34078 6244 34130
rect 6188 34020 6244 34078
rect 6748 34020 6804 34030
rect 6188 34018 6804 34020
rect 6188 33966 6750 34018
rect 6802 33966 6804 34018
rect 6188 33964 6804 33966
rect 6076 33348 6132 33358
rect 5628 33346 6132 33348
rect 5628 33294 6078 33346
rect 6130 33294 6132 33346
rect 5628 33292 6132 33294
rect 4396 33170 4452 33180
rect 4620 33234 4676 33246
rect 4620 33182 4622 33234
rect 4674 33182 4676 33234
rect 2492 33124 2548 33134
rect 1820 32510 1822 32562
rect 1874 32510 1876 32562
rect 1820 32004 1876 32510
rect 2268 32562 2324 32574
rect 2268 32510 2270 32562
rect 2322 32510 2324 32562
rect 2268 31948 2324 32510
rect 1820 30210 1876 31948
rect 2156 31892 2324 31948
rect 2156 31666 2212 31892
rect 2492 31778 2548 33068
rect 3500 33124 3556 33134
rect 3500 33030 3556 33068
rect 2492 31726 2494 31778
rect 2546 31726 2548 31778
rect 2492 31714 2548 31726
rect 3948 32788 4004 32798
rect 4620 32788 4676 33182
rect 5068 33236 5124 33246
rect 4732 32788 4788 32798
rect 4620 32732 4732 32788
rect 3948 32002 4004 32732
rect 4732 32694 4788 32732
rect 5068 32452 5124 33180
rect 5740 32562 5796 32574
rect 5740 32510 5742 32562
rect 5794 32510 5796 32562
rect 5180 32452 5236 32462
rect 5068 32450 5236 32452
rect 5068 32398 5182 32450
rect 5234 32398 5236 32450
rect 5068 32396 5236 32398
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 3948 31950 3950 32002
rect 4002 31950 4004 32002
rect 2156 31614 2158 31666
rect 2210 31614 2212 31666
rect 2156 31602 2212 31614
rect 2492 31556 2548 31566
rect 1820 30158 1822 30210
rect 1874 30158 1876 30210
rect 1820 28642 1876 30158
rect 2156 31106 2212 31118
rect 2156 31054 2158 31106
rect 2210 31054 2212 31106
rect 2156 30212 2212 31054
rect 2492 31106 2548 31500
rect 3612 31556 3668 31566
rect 3612 31462 3668 31500
rect 2492 31054 2494 31106
rect 2546 31054 2548 31106
rect 2492 31042 2548 31054
rect 3948 30996 4004 31950
rect 5068 31892 5124 32396
rect 5180 32386 5236 32396
rect 5740 32340 5796 32510
rect 5964 32340 6020 32350
rect 5740 32338 6020 32340
rect 5740 32286 5966 32338
rect 6018 32286 6020 32338
rect 5740 32284 6020 32286
rect 5964 32274 6020 32284
rect 6076 32004 6132 33292
rect 4956 31836 5124 31892
rect 5740 31892 5796 31902
rect 4732 31780 4788 31790
rect 4956 31780 5012 31836
rect 4732 31778 5012 31780
rect 4732 31726 4734 31778
rect 4786 31726 5012 31778
rect 4732 31724 5012 31726
rect 4508 31668 4564 31678
rect 3948 30930 4004 30940
rect 4396 31666 4564 31668
rect 4396 31614 4510 31666
rect 4562 31614 4564 31666
rect 4396 31612 4564 31614
rect 4396 31106 4452 31612
rect 4508 31602 4564 31612
rect 4396 31054 4398 31106
rect 4450 31054 4452 31106
rect 4396 30772 4452 31054
rect 4284 30716 4452 30772
rect 4732 30772 4788 31724
rect 5404 31668 5460 31678
rect 5404 31218 5460 31612
rect 5404 31166 5406 31218
rect 5458 31166 5460 31218
rect 5404 31154 5460 31166
rect 4844 31108 4900 31118
rect 4844 31014 4900 31052
rect 5740 31108 5796 31836
rect 5068 30996 5124 31006
rect 5068 30902 5124 30940
rect 4732 30716 4900 30772
rect 2268 30212 2324 30222
rect 2156 30210 2324 30212
rect 2156 30158 2270 30210
rect 2322 30158 2324 30210
rect 2156 30156 2324 30158
rect 2268 30146 2324 30156
rect 4284 29876 4340 30716
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4732 29986 4788 29998
rect 4732 29934 4734 29986
rect 4786 29934 4788 29986
rect 4732 29876 4788 29934
rect 4284 29820 4788 29876
rect 1820 28590 1822 28642
rect 1874 28590 1876 28642
rect 1820 28578 1876 28590
rect 2492 28642 2548 28654
rect 2492 28590 2494 28642
rect 2546 28590 2548 28642
rect 2492 28082 2548 28590
rect 2492 28030 2494 28082
rect 2546 28030 2548 28082
rect 2492 28018 2548 28030
rect 2828 27860 2884 27870
rect 2828 27766 2884 27804
rect 4060 27860 4116 27870
rect 4284 27860 4340 29820
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4844 28868 4900 30716
rect 5740 30210 5796 31052
rect 5964 30996 6020 31006
rect 6076 30996 6132 31948
rect 5964 30994 6076 30996
rect 5964 30942 5966 30994
rect 6018 30942 6076 30994
rect 5964 30940 6076 30942
rect 5964 30930 6020 30940
rect 5740 30158 5742 30210
rect 5794 30158 5796 30210
rect 5740 30146 5796 30158
rect 4732 28812 4900 28868
rect 4396 27860 4452 27870
rect 4284 27858 4452 27860
rect 4284 27806 4398 27858
rect 4450 27806 4452 27858
rect 4284 27804 4452 27806
rect 4732 27860 4788 28812
rect 4844 28642 4900 28654
rect 4844 28590 4846 28642
rect 4898 28590 4900 28642
rect 4844 28084 4900 28590
rect 5180 28084 5236 28094
rect 4844 28028 5180 28084
rect 5180 27970 5236 28028
rect 5180 27918 5182 27970
rect 5234 27918 5236 27970
rect 5180 27906 5236 27918
rect 4844 27860 4900 27870
rect 4732 27858 4900 27860
rect 4732 27806 4846 27858
rect 4898 27806 4900 27858
rect 4732 27804 4900 27806
rect 4060 27766 4116 27804
rect 4396 27794 4452 27804
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4172 27076 4228 27086
rect 2604 26964 2660 26974
rect 2604 26870 2660 26908
rect 3836 26964 3892 27002
rect 4172 26982 4228 27020
rect 4844 27074 4900 27804
rect 6076 27858 6132 30940
rect 6076 27806 6078 27858
rect 6130 27806 6132 27858
rect 6076 27794 6132 27806
rect 6188 32450 6244 33964
rect 6748 33954 6804 33964
rect 6636 33348 6692 33358
rect 6636 33346 7028 33348
rect 6636 33294 6638 33346
rect 6690 33294 7028 33346
rect 6636 33292 7028 33294
rect 6636 33282 6692 33292
rect 6972 32786 7028 33292
rect 6972 32734 6974 32786
rect 7026 32734 7028 32786
rect 6972 32722 7028 32734
rect 8092 32676 8148 32686
rect 7308 32564 7364 32574
rect 7756 32564 7812 32574
rect 7308 32562 7812 32564
rect 7308 32510 7310 32562
rect 7362 32510 7758 32562
rect 7810 32510 7812 32562
rect 7308 32508 7812 32510
rect 7308 32498 7364 32508
rect 7756 32498 7812 32508
rect 8092 32562 8148 32620
rect 8092 32510 8094 32562
rect 8146 32510 8148 32562
rect 8092 32498 8148 32510
rect 6188 32398 6190 32450
rect 6242 32398 6244 32450
rect 6188 32338 6244 32398
rect 6188 32286 6190 32338
rect 6242 32286 6244 32338
rect 4844 27022 4846 27074
rect 4898 27022 4900 27074
rect 4844 27010 4900 27022
rect 5628 27076 5684 27086
rect 5628 26982 5684 27020
rect 3836 26898 3892 26908
rect 4732 26962 4788 26974
rect 4732 26910 4734 26962
rect 4786 26910 4788 26962
rect 2268 26850 2324 26862
rect 2268 26798 2270 26850
rect 2322 26798 2324 26850
rect 1820 26292 1876 26302
rect 1820 26290 1988 26292
rect 1820 26238 1822 26290
rect 1874 26238 1988 26290
rect 1820 26236 1988 26238
rect 1820 26226 1876 26236
rect 1932 24722 1988 26236
rect 2268 26290 2324 26798
rect 2268 26238 2270 26290
rect 2322 26238 2324 26290
rect 2268 26226 2324 26238
rect 4732 26178 4788 26910
rect 5180 26292 5236 26302
rect 5180 26198 5236 26236
rect 5740 26292 5796 26302
rect 4732 26126 4734 26178
rect 4786 26126 4788 26178
rect 1932 24670 1934 24722
rect 1986 24670 1988 24722
rect 1820 23156 1876 23166
rect 1932 23156 1988 24670
rect 1820 23154 1988 23156
rect 1820 23102 1822 23154
rect 1874 23102 1988 23154
rect 1820 23100 1988 23102
rect 1820 23090 1876 23100
rect 1932 22484 1988 23100
rect 1932 21586 1988 22428
rect 1932 21534 1934 21586
rect 1986 21534 1988 21586
rect 1820 19236 1876 19246
rect 1932 19236 1988 21534
rect 1820 19234 1988 19236
rect 1820 19182 1822 19234
rect 1874 19182 1988 19234
rect 1820 19180 1988 19182
rect 2044 26068 2100 26078
rect 4732 26068 4788 26126
rect 1820 19170 1876 19180
rect 1708 16882 1764 16894
rect 1708 16830 1710 16882
rect 1762 16830 1764 16882
rect 1708 14530 1764 16830
rect 1708 14478 1710 14530
rect 1762 14478 1764 14530
rect 1708 13748 1764 14478
rect 1708 12178 1764 13692
rect 1708 12126 1710 12178
rect 1762 12126 1764 12178
rect 1708 10610 1764 12126
rect 1708 10558 1710 10610
rect 1762 10558 1764 10610
rect 1708 8258 1764 10558
rect 2044 8428 2100 26012
rect 4284 26012 4788 26068
rect 2604 24722 2660 24734
rect 2604 24670 2606 24722
rect 2658 24670 2660 24722
rect 2604 23826 2660 24670
rect 4172 23940 4228 23950
rect 4284 23940 4340 26012
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4956 24612 5012 24622
rect 4844 24610 5012 24612
rect 4844 24558 4958 24610
rect 5010 24558 5012 24610
rect 4844 24556 5012 24558
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4228 23884 4340 23940
rect 4172 23846 4228 23884
rect 2604 23774 2606 23826
rect 2658 23774 2660 23826
rect 2604 23762 2660 23774
rect 2940 23828 2996 23838
rect 2940 23734 2996 23772
rect 3836 23828 3892 23838
rect 3836 23734 3892 23772
rect 4844 23828 4900 24556
rect 4956 24546 5012 24556
rect 5516 24612 5572 24622
rect 5628 24612 5684 24622
rect 5516 24610 5628 24612
rect 5516 24558 5518 24610
rect 5570 24558 5628 24610
rect 5516 24556 5628 24558
rect 5516 24546 5572 24556
rect 4844 23734 4900 23772
rect 4956 23938 5012 23950
rect 4956 23886 4958 23938
rect 5010 23886 5012 23938
rect 4956 23268 5012 23886
rect 4956 23202 5012 23212
rect 2268 23154 2324 23166
rect 2268 23102 2270 23154
rect 2322 23102 2324 23154
rect 2268 22258 2324 23102
rect 4732 23156 4788 23166
rect 4732 23062 4788 23100
rect 5516 23156 5572 23166
rect 2604 22932 2660 22942
rect 2604 22370 2660 22876
rect 5292 22932 5348 22942
rect 5292 22838 5348 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 2604 22318 2606 22370
rect 2658 22318 2660 22370
rect 2604 22306 2660 22318
rect 4956 22372 5012 22382
rect 5012 22316 5124 22372
rect 4956 22278 5012 22316
rect 2268 22206 2270 22258
rect 2322 22206 2324 22258
rect 2268 22194 2324 22206
rect 2492 21586 2548 21598
rect 2492 21534 2494 21586
rect 2546 21534 2548 21586
rect 2492 20692 2548 21534
rect 4844 21588 4900 21598
rect 4844 21494 4900 21532
rect 2940 21364 2996 21374
rect 2940 20802 2996 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 2940 20750 2942 20802
rect 2994 20750 2996 20802
rect 2940 20738 2996 20750
rect 5068 20914 5124 22316
rect 5516 21588 5572 23100
rect 5628 23154 5684 24556
rect 5628 23102 5630 23154
rect 5682 23102 5684 23154
rect 5628 23090 5684 23102
rect 5740 24050 5796 26236
rect 5740 23998 5742 24050
rect 5794 23998 5796 24050
rect 5740 22372 5796 23998
rect 5852 23268 5908 23278
rect 5852 23174 5908 23212
rect 5740 22306 5796 22316
rect 5740 22148 5796 22158
rect 5740 22054 5796 22092
rect 6188 22148 6244 32286
rect 8428 31892 8484 35644
rect 8428 31826 8484 31836
rect 8540 34804 8596 34814
rect 8764 34804 8820 36318
rect 8988 36372 9044 39006
rect 9212 39396 9268 39406
rect 9324 39396 9380 39676
rect 9212 39394 9380 39396
rect 9212 39342 9214 39394
rect 9266 39342 9380 39394
rect 9212 39340 9380 39342
rect 9212 38836 9268 39340
rect 9660 38836 9716 38846
rect 9212 38780 9660 38836
rect 9660 38742 9716 38780
rect 9884 38668 9940 42252
rect 9996 42082 10052 42094
rect 9996 42030 9998 42082
rect 10050 42030 10052 42082
rect 9996 41186 10052 42030
rect 9996 41134 9998 41186
rect 10050 41134 10052 41186
rect 9996 41122 10052 41134
rect 9996 40180 10052 40190
rect 9996 40086 10052 40124
rect 9772 38612 9940 38668
rect 10108 38612 10164 38622
rect 9660 38164 9716 38174
rect 9660 38070 9716 38108
rect 9436 37940 9492 37950
rect 9436 37846 9492 37884
rect 9100 37268 9156 37278
rect 9100 37174 9156 37212
rect 9100 36372 9156 36382
rect 8988 36370 9268 36372
rect 8988 36318 9102 36370
rect 9154 36318 9268 36370
rect 8988 36316 9268 36318
rect 9100 36306 9156 36316
rect 9212 36260 9268 36316
rect 9212 36204 9716 36260
rect 8540 34802 8820 34804
rect 8540 34750 8542 34802
rect 8594 34750 8820 34802
rect 8540 34748 8820 34750
rect 8876 35924 8932 35934
rect 8876 35588 8932 35868
rect 9660 35810 9716 36204
rect 9660 35758 9662 35810
rect 9714 35758 9716 35810
rect 9660 35746 9716 35758
rect 8876 34802 8932 35532
rect 9772 35308 9828 38612
rect 9996 37826 10052 37838
rect 9996 37774 9998 37826
rect 10050 37774 10052 37826
rect 9996 37380 10052 37774
rect 9996 37314 10052 37324
rect 10108 37378 10164 38556
rect 10220 37490 10276 42700
rect 10444 42196 10500 44380
rect 10892 43764 10948 44382
rect 10892 43428 10948 43708
rect 10892 43362 10948 43372
rect 10220 37438 10222 37490
rect 10274 37438 10276 37490
rect 10220 37426 10276 37438
rect 10332 37940 10388 37950
rect 10108 37326 10110 37378
rect 10162 37326 10164 37378
rect 10108 37268 10164 37326
rect 9884 37154 9940 37166
rect 9884 37102 9886 37154
rect 9938 37102 9940 37154
rect 9884 35476 9940 37102
rect 10108 37044 10164 37212
rect 9884 35410 9940 35420
rect 9996 36988 10164 37044
rect 8876 34750 8878 34802
rect 8930 34750 8932 34802
rect 6524 30996 6580 31006
rect 6524 30994 6916 30996
rect 6524 30942 6526 30994
rect 6578 30942 6916 30994
rect 6524 30940 6916 30942
rect 6524 30930 6580 30940
rect 6860 30098 6916 30940
rect 8428 30324 8484 30334
rect 8428 30230 8484 30268
rect 6860 30046 6862 30098
rect 6914 30046 6916 30098
rect 6860 30034 6916 30046
rect 7196 30100 7252 30110
rect 8092 30100 8148 30110
rect 7196 30098 8148 30100
rect 7196 30046 7198 30098
rect 7250 30046 8094 30098
rect 8146 30046 8148 30098
rect 7196 30044 8148 30046
rect 7196 30034 7252 30044
rect 8092 30034 8148 30044
rect 8316 28756 8372 28766
rect 6636 28644 6692 28654
rect 6636 27858 6692 28588
rect 8204 28644 8260 28654
rect 8204 28550 8260 28588
rect 8316 28642 8372 28700
rect 8316 28590 8318 28642
rect 8370 28590 8372 28642
rect 8316 28578 8372 28590
rect 8540 28532 8596 34748
rect 8876 34738 8932 34750
rect 9548 35252 9828 35308
rect 8652 33572 8708 33582
rect 8652 32674 8708 33516
rect 8988 33572 9044 33582
rect 8988 33458 9044 33516
rect 8988 33406 8990 33458
rect 9042 33406 9044 33458
rect 8988 33394 9044 33406
rect 8652 32622 8654 32674
rect 8706 32622 8708 32674
rect 8652 32610 8708 32622
rect 8876 32676 8932 32686
rect 8764 32562 8820 32574
rect 8764 32510 8766 32562
rect 8818 32510 8820 32562
rect 8764 30100 8820 32510
rect 8876 31218 8932 32620
rect 8876 31166 8878 31218
rect 8930 31166 8932 31218
rect 8876 30100 8932 31166
rect 8988 30100 9044 30110
rect 8876 30098 9044 30100
rect 8876 30046 8990 30098
rect 9042 30046 9044 30098
rect 8876 30044 9044 30046
rect 8764 30006 8820 30044
rect 8988 30034 9044 30044
rect 8764 28644 8820 28654
rect 8988 28644 9044 28654
rect 8764 28642 8932 28644
rect 8764 28590 8766 28642
rect 8818 28590 8932 28642
rect 8764 28588 8932 28590
rect 8764 28578 8820 28588
rect 8652 28532 8708 28542
rect 8540 28476 8652 28532
rect 8652 28466 8708 28476
rect 8092 28420 8148 28430
rect 8092 28418 8260 28420
rect 8092 28366 8094 28418
rect 8146 28366 8260 28418
rect 8092 28364 8260 28366
rect 8092 28354 8148 28364
rect 6636 27806 6638 27858
rect 6690 27806 6692 27858
rect 6636 27794 6692 27806
rect 7868 27524 7924 27534
rect 7644 27188 7700 27198
rect 7644 23716 7700 27132
rect 7756 24052 7812 24062
rect 7756 23958 7812 23996
rect 7868 23938 7924 27468
rect 8204 27188 8260 28364
rect 8876 27860 8932 28588
rect 8988 28082 9044 28588
rect 9548 28308 9604 35252
rect 9660 34692 9716 34702
rect 9660 34020 9716 34636
rect 9996 34132 10052 36988
rect 10108 36258 10164 36270
rect 10108 36206 10110 36258
rect 10162 36206 10164 36258
rect 10108 35812 10164 36206
rect 10332 36036 10388 37884
rect 10444 37492 10500 42140
rect 10668 42866 10724 42878
rect 10668 42814 10670 42866
rect 10722 42814 10724 42866
rect 10668 42644 10724 42814
rect 11116 42756 11172 42766
rect 11116 42662 11172 42700
rect 10556 40514 10612 40526
rect 10556 40462 10558 40514
rect 10610 40462 10612 40514
rect 10556 39844 10612 40462
rect 10668 40402 10724 42588
rect 11340 42084 11396 45164
rect 11676 44434 11732 45724
rect 12012 45668 12068 45838
rect 12684 45890 12740 45902
rect 12684 45838 12686 45890
rect 12738 45838 12740 45890
rect 12684 45780 12740 45838
rect 12684 45714 12740 45724
rect 12796 45778 12852 47180
rect 12908 47170 12964 47180
rect 13580 47234 13636 47246
rect 13580 47182 13582 47234
rect 13634 47182 13636 47234
rect 12908 46900 12964 46910
rect 13580 46900 13636 47182
rect 12964 46844 13636 46900
rect 12908 46806 12964 46844
rect 13132 46674 13188 46844
rect 13132 46622 13134 46674
rect 13186 46622 13188 46674
rect 13132 46610 13188 46622
rect 13916 46674 13972 46686
rect 13916 46622 13918 46674
rect 13970 46622 13972 46674
rect 12796 45726 12798 45778
rect 12850 45726 12852 45778
rect 12012 45602 12068 45612
rect 11676 44382 11678 44434
rect 11730 44382 11732 44434
rect 11676 44370 11732 44382
rect 12124 44098 12180 44110
rect 12124 44046 12126 44098
rect 12178 44046 12180 44098
rect 12012 43540 12068 43550
rect 12012 43446 12068 43484
rect 11564 43428 11620 43438
rect 11564 43334 11620 43372
rect 12124 43428 12180 44046
rect 12348 43764 12404 43774
rect 12236 43652 12292 43662
rect 12348 43652 12740 43708
rect 12236 43558 12292 43596
rect 11452 42754 11508 42766
rect 11452 42702 11454 42754
rect 11506 42702 11508 42754
rect 11452 42308 11508 42702
rect 12012 42756 12068 42766
rect 12124 42756 12180 43372
rect 12068 42700 12180 42756
rect 12684 43538 12740 43652
rect 12684 43486 12686 43538
rect 12738 43486 12740 43538
rect 12012 42662 12068 42700
rect 11452 42242 11508 42252
rect 11340 42028 12068 42084
rect 10668 40350 10670 40402
rect 10722 40350 10724 40402
rect 10668 40338 10724 40350
rect 11564 40964 11620 40974
rect 10556 39778 10612 39788
rect 11564 39844 11620 40908
rect 10556 39396 10612 39406
rect 10556 38274 10612 39340
rect 11564 39058 11620 39788
rect 11564 39006 11566 39058
rect 11618 39006 11620 39058
rect 11564 38994 11620 39006
rect 11676 39394 11732 39406
rect 11676 39342 11678 39394
rect 11730 39342 11732 39394
rect 10780 38836 10836 38846
rect 10780 38742 10836 38780
rect 11340 38722 11396 38734
rect 11340 38670 11342 38722
rect 11394 38670 11396 38722
rect 11340 38668 11396 38670
rect 10556 38222 10558 38274
rect 10610 38222 10612 38274
rect 10556 38210 10612 38222
rect 10780 38612 11396 38668
rect 11676 38724 11732 39342
rect 11900 39394 11956 39406
rect 11900 39342 11902 39394
rect 11954 39342 11956 39394
rect 11788 39284 11844 39294
rect 11788 39058 11844 39228
rect 11788 39006 11790 39058
rect 11842 39006 11844 39058
rect 11788 38994 11844 39006
rect 11900 38946 11956 39342
rect 11900 38894 11902 38946
rect 11954 38894 11956 38946
rect 11900 38882 11956 38894
rect 11676 38658 11732 38668
rect 10780 37604 10836 38612
rect 12012 38164 12068 42028
rect 12460 40964 12516 40974
rect 12684 40964 12740 43486
rect 12796 41188 12852 45726
rect 13692 45666 13748 45678
rect 13692 45614 13694 45666
rect 13746 45614 13748 45666
rect 13692 45106 13748 45614
rect 13916 45330 13972 46622
rect 16268 46564 16324 46574
rect 16156 46562 16324 46564
rect 16156 46510 16270 46562
rect 16322 46510 16324 46562
rect 16156 46508 16324 46510
rect 13916 45278 13918 45330
rect 13970 45278 13972 45330
rect 13916 45266 13972 45278
rect 14028 45890 14084 45902
rect 14028 45838 14030 45890
rect 14082 45838 14084 45890
rect 13692 45054 13694 45106
rect 13746 45054 13748 45106
rect 13692 45042 13748 45054
rect 13132 43652 13188 43662
rect 13132 43538 13188 43596
rect 13132 43486 13134 43538
rect 13186 43486 13188 43538
rect 13132 43474 13188 43486
rect 13580 43540 13636 43550
rect 13580 42978 13636 43484
rect 13580 42926 13582 42978
rect 13634 42926 13636 42978
rect 13580 42914 13636 42926
rect 13916 42756 13972 42766
rect 13916 42662 13972 42700
rect 14028 42308 14084 45838
rect 14364 45780 14420 45790
rect 14364 42754 14420 45724
rect 14812 45780 14868 45790
rect 14812 45686 14868 45724
rect 15708 45780 15764 45790
rect 15596 43426 15652 43438
rect 15596 43374 15598 43426
rect 15650 43374 15652 43426
rect 14364 42702 14366 42754
rect 14418 42702 14420 42754
rect 14364 42690 14420 42702
rect 15484 42754 15540 42766
rect 15484 42702 15486 42754
rect 15538 42702 15540 42754
rect 14028 42242 14084 42252
rect 14700 42642 14756 42654
rect 14700 42590 14702 42642
rect 14754 42590 14756 42642
rect 14700 42308 14756 42590
rect 14700 42242 14756 42252
rect 15484 41972 15540 42702
rect 15596 42084 15652 43374
rect 15596 42018 15652 42028
rect 15484 41906 15540 41916
rect 12796 41132 13188 41188
rect 12908 40964 12964 40974
rect 12684 40962 12964 40964
rect 12684 40910 12910 40962
rect 12962 40910 12964 40962
rect 12684 40908 12964 40910
rect 12460 40870 12516 40908
rect 12796 40628 12852 40638
rect 12236 40516 12292 40526
rect 12124 40404 12180 40414
rect 12124 38836 12180 40348
rect 12236 39842 12292 40460
rect 12796 40402 12852 40572
rect 12796 40350 12798 40402
rect 12850 40350 12852 40402
rect 12796 40338 12852 40350
rect 12908 40404 12964 40908
rect 12908 40338 12964 40348
rect 12236 39790 12238 39842
rect 12290 39790 12292 39842
rect 12236 39778 12292 39790
rect 12460 39508 12516 39518
rect 12460 39414 12516 39452
rect 13020 39396 13076 39406
rect 12908 39394 13076 39396
rect 12908 39342 13022 39394
rect 13074 39342 13076 39394
rect 12908 39340 13076 39342
rect 12908 39284 12964 39340
rect 13020 39330 13076 39340
rect 13132 39396 13188 41132
rect 15036 41186 15092 41198
rect 15036 41134 15038 41186
rect 15090 41134 15092 41186
rect 14364 40962 14420 40974
rect 14364 40910 14366 40962
rect 14418 40910 14420 40962
rect 14364 39732 14420 40910
rect 14476 40962 14532 40974
rect 14476 40910 14478 40962
rect 14530 40910 14532 40962
rect 14476 40628 14532 40910
rect 14588 40962 14644 40974
rect 14588 40910 14590 40962
rect 14642 40910 14644 40962
rect 14588 40740 14644 40910
rect 14588 40674 14644 40684
rect 14476 40562 14532 40572
rect 15036 40628 15092 41134
rect 15036 40562 15092 40572
rect 15260 41074 15316 41086
rect 15260 41022 15262 41074
rect 15314 41022 15316 41074
rect 15260 40626 15316 41022
rect 15372 40964 15428 40974
rect 15372 40870 15428 40908
rect 15260 40574 15262 40626
rect 15314 40574 15316 40626
rect 15260 40562 15316 40574
rect 15484 40628 15540 40638
rect 15484 40534 15540 40572
rect 15708 40516 15764 45724
rect 16156 45780 16212 46508
rect 16268 46498 16324 46508
rect 16828 46116 16884 48972
rect 17612 49028 17668 49038
rect 18284 49028 18340 49038
rect 17388 48802 17444 48814
rect 17388 48750 17390 48802
rect 17442 48750 17444 48802
rect 17276 48244 17332 48254
rect 17276 47682 17332 48188
rect 17276 47630 17278 47682
rect 17330 47630 17332 47682
rect 17276 47618 17332 47630
rect 17388 47348 17444 48750
rect 17612 48466 17668 48972
rect 17612 48414 17614 48466
rect 17666 48414 17668 48466
rect 17612 48402 17668 48414
rect 18172 49026 18340 49028
rect 18172 48974 18286 49026
rect 18338 48974 18340 49026
rect 18172 48972 18340 48974
rect 18172 48466 18228 48972
rect 18284 48962 18340 48972
rect 21420 49026 21476 49644
rect 21532 49634 21588 49644
rect 21868 49028 21924 49038
rect 21420 48974 21422 49026
rect 21474 48974 21476 49026
rect 20748 48802 20804 48814
rect 20748 48750 20750 48802
rect 20802 48750 20804 48802
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 18172 48414 18174 48466
rect 18226 48414 18228 48466
rect 18172 48402 18228 48414
rect 18396 48356 18452 48366
rect 17612 47460 17668 47470
rect 18396 47460 18452 48300
rect 19852 48354 19908 48366
rect 19852 48302 19854 48354
rect 19906 48302 19908 48354
rect 18508 48244 18564 48254
rect 18956 48244 19012 48254
rect 18508 48242 19012 48244
rect 18508 48190 18510 48242
rect 18562 48190 18958 48242
rect 19010 48190 19012 48242
rect 18508 48188 19012 48190
rect 18508 48178 18564 48188
rect 18956 48178 19012 48188
rect 17612 47458 17780 47460
rect 17612 47406 17614 47458
rect 17666 47406 17780 47458
rect 17612 47404 17780 47406
rect 17612 47394 17668 47404
rect 17388 47282 17444 47292
rect 17388 46788 17444 46798
rect 16268 46060 16828 46116
rect 16268 45890 16324 46060
rect 16828 46022 16884 46060
rect 16940 46786 17444 46788
rect 16940 46734 17390 46786
rect 17442 46734 17444 46786
rect 16940 46732 17444 46734
rect 16268 45838 16270 45890
rect 16322 45838 16324 45890
rect 16268 45826 16324 45838
rect 16716 45892 16772 45902
rect 16716 45890 16884 45892
rect 16716 45838 16718 45890
rect 16770 45838 16884 45890
rect 16716 45836 16884 45838
rect 16716 45826 16772 45836
rect 16828 45780 16884 45836
rect 16940 45780 16996 46732
rect 17388 46722 17444 46732
rect 16828 45724 16996 45780
rect 17612 46674 17668 46686
rect 17612 46622 17614 46674
rect 17666 46622 17668 46674
rect 16156 45714 16212 45724
rect 17500 45332 17556 45342
rect 17612 45332 17668 46622
rect 17724 45444 17780 47404
rect 18284 47458 18452 47460
rect 18284 47406 18398 47458
rect 18450 47406 18452 47458
rect 18284 47404 18452 47406
rect 18172 47348 18228 47358
rect 18172 47254 18228 47292
rect 17724 45378 17780 45388
rect 17500 45330 17668 45332
rect 17500 45278 17502 45330
rect 17554 45278 17668 45330
rect 17500 45276 17668 45278
rect 17500 45266 17556 45276
rect 18284 45106 18340 47404
rect 18396 47394 18452 47404
rect 19292 48018 19348 48030
rect 19292 47966 19294 48018
rect 19346 47966 19348 48018
rect 18620 47348 18676 47358
rect 18508 45444 18564 45454
rect 18508 45218 18564 45388
rect 18508 45166 18510 45218
rect 18562 45166 18564 45218
rect 18508 45154 18564 45166
rect 18284 45054 18286 45106
rect 18338 45054 18340 45106
rect 17836 44884 17892 44894
rect 17836 44790 17892 44828
rect 18284 44436 18340 45054
rect 18396 44436 18452 44446
rect 18284 44434 18452 44436
rect 18284 44382 18398 44434
rect 18450 44382 18452 44434
rect 18284 44380 18452 44382
rect 18396 44370 18452 44380
rect 17948 44098 18004 44110
rect 17948 44046 17950 44098
rect 18002 44046 18004 44098
rect 17948 43650 18004 44046
rect 17948 43598 17950 43650
rect 18002 43598 18004 43650
rect 17612 43428 17668 43438
rect 17948 43428 18004 43598
rect 17612 43426 17780 43428
rect 17612 43374 17614 43426
rect 17666 43374 17780 43426
rect 17612 43372 17780 43374
rect 17612 43362 17668 43372
rect 17724 43204 17780 43372
rect 17948 43362 18004 43372
rect 18172 43538 18228 43550
rect 18172 43486 18174 43538
rect 18226 43486 18228 43538
rect 18172 43204 18228 43486
rect 17724 43148 18228 43204
rect 16044 42756 16100 42766
rect 16044 42754 16436 42756
rect 16044 42702 16046 42754
rect 16098 42702 16436 42754
rect 16044 42700 16436 42702
rect 16044 42690 16100 42700
rect 16268 41972 16324 41982
rect 16268 41186 16324 41916
rect 16268 41134 16270 41186
rect 16322 41134 16324 41186
rect 16268 41122 16324 41134
rect 15708 40422 15764 40460
rect 15820 40402 15876 40414
rect 15820 40350 15822 40402
rect 15874 40350 15876 40402
rect 14364 39676 14980 39732
rect 13132 39330 13188 39340
rect 13244 39508 13300 39518
rect 12124 38770 12180 38780
rect 12236 38834 12292 38846
rect 12236 38782 12238 38834
rect 12290 38782 12292 38834
rect 12236 38724 12292 38782
rect 12684 38836 12740 38846
rect 12236 38658 12292 38668
rect 12348 38724 12404 38734
rect 12348 38722 12628 38724
rect 12348 38670 12350 38722
rect 12402 38670 12628 38722
rect 12348 38668 12628 38670
rect 12348 38658 12404 38668
rect 12236 38164 12292 38174
rect 12012 38162 12292 38164
rect 12012 38110 12238 38162
rect 12290 38110 12292 38162
rect 12012 38108 12292 38110
rect 12236 38098 12292 38108
rect 11452 38052 11508 38062
rect 11340 38050 11508 38052
rect 11340 37998 11454 38050
rect 11506 37998 11508 38050
rect 11340 37996 11508 37998
rect 11228 37938 11284 37950
rect 11228 37886 11230 37938
rect 11282 37886 11284 37938
rect 10892 37828 10948 37838
rect 11228 37828 11284 37886
rect 10892 37826 11284 37828
rect 10892 37774 10894 37826
rect 10946 37774 11284 37826
rect 10892 37772 11284 37774
rect 10892 37762 10948 37772
rect 10780 37548 11172 37604
rect 10444 37436 10612 37492
rect 10444 37268 10500 37278
rect 10444 37174 10500 37212
rect 10556 36484 10612 37436
rect 10892 37378 10948 37390
rect 10892 37326 10894 37378
rect 10946 37326 10948 37378
rect 10668 37266 10724 37278
rect 10668 37214 10670 37266
rect 10722 37214 10724 37266
rect 10668 37156 10724 37214
rect 10668 37090 10724 37100
rect 10780 37044 10836 37054
rect 10668 36484 10724 36494
rect 10556 36482 10724 36484
rect 10556 36430 10670 36482
rect 10722 36430 10724 36482
rect 10556 36428 10724 36430
rect 10668 36418 10724 36428
rect 10556 36258 10612 36270
rect 10556 36206 10558 36258
rect 10610 36206 10612 36258
rect 10556 36148 10612 36206
rect 10668 36148 10724 36158
rect 10556 36092 10668 36148
rect 10668 36082 10724 36092
rect 10332 35980 10612 36036
rect 10220 35812 10276 35822
rect 10108 35810 10276 35812
rect 10108 35758 10222 35810
rect 10274 35758 10276 35810
rect 10108 35756 10276 35758
rect 10220 35700 10276 35756
rect 10220 35634 10276 35644
rect 10444 35588 10500 35598
rect 10444 35494 10500 35532
rect 10332 35028 10388 35038
rect 10332 34934 10388 34972
rect 10556 35026 10612 35980
rect 10780 35922 10836 36988
rect 10780 35870 10782 35922
rect 10834 35870 10836 35922
rect 10780 35858 10836 35870
rect 10556 34974 10558 35026
rect 10610 34974 10612 35026
rect 10444 34356 10500 34366
rect 10556 34356 10612 34974
rect 10444 34354 10612 34356
rect 10444 34302 10446 34354
rect 10498 34302 10612 34354
rect 10444 34300 10612 34302
rect 10668 35476 10724 35486
rect 10444 34290 10500 34300
rect 10668 34244 10724 35420
rect 10892 35140 10948 37326
rect 11004 37380 11060 37418
rect 11004 37314 11060 37324
rect 10892 35074 10948 35084
rect 11004 36260 11060 36270
rect 11116 36260 11172 37548
rect 11228 37380 11284 37390
rect 11228 36594 11284 37324
rect 11228 36542 11230 36594
rect 11282 36542 11284 36594
rect 11228 36530 11284 36542
rect 11340 37266 11396 37996
rect 11452 37986 11508 37996
rect 12348 38050 12404 38062
rect 12348 37998 12350 38050
rect 12402 37998 12404 38050
rect 11340 37214 11342 37266
rect 11394 37214 11396 37266
rect 11004 36258 11172 36260
rect 11004 36206 11006 36258
rect 11058 36206 11172 36258
rect 11004 36204 11172 36206
rect 11228 36258 11284 36270
rect 11228 36206 11230 36258
rect 11282 36206 11284 36258
rect 10780 34916 10836 34926
rect 10780 34822 10836 34860
rect 11004 34692 11060 36204
rect 11228 35476 11284 36206
rect 11228 35410 11284 35420
rect 11340 35364 11396 37214
rect 11564 37940 11620 37950
rect 11340 35298 11396 35308
rect 11452 37154 11508 37166
rect 11452 37102 11454 37154
rect 11506 37102 11508 37154
rect 11116 35026 11172 35038
rect 11452 35028 11508 37102
rect 11564 36370 11620 37884
rect 12124 37940 12180 37950
rect 11564 36318 11566 36370
rect 11618 36318 11620 36370
rect 11564 36306 11620 36318
rect 11676 37492 11732 37502
rect 11676 35476 11732 37436
rect 12012 37380 12068 37390
rect 12012 37286 12068 37324
rect 11788 37268 11844 37278
rect 11788 37174 11844 37212
rect 11900 36370 11956 36382
rect 11900 36318 11902 36370
rect 11954 36318 11956 36370
rect 11900 36260 11956 36318
rect 11900 36194 11956 36204
rect 11116 34974 11118 35026
rect 11170 34974 11172 35026
rect 11116 34916 11172 34974
rect 11116 34850 11172 34860
rect 11228 34972 11508 35028
rect 11564 35420 11732 35476
rect 11900 35700 11956 35710
rect 10556 34188 10724 34244
rect 10780 34636 11060 34692
rect 9996 34076 10164 34132
rect 9660 33954 9716 33964
rect 9884 34018 9940 34030
rect 9884 33966 9886 34018
rect 9938 33966 9940 34018
rect 9660 32788 9716 32798
rect 9660 32694 9716 32732
rect 9660 30996 9716 31006
rect 9660 30902 9716 30940
rect 9884 29428 9940 33966
rect 10108 33796 10164 34076
rect 9996 33740 10164 33796
rect 9996 32788 10052 33740
rect 10332 33572 10388 33582
rect 10332 33346 10388 33516
rect 10332 33294 10334 33346
rect 10386 33294 10388 33346
rect 10332 33282 10388 33294
rect 10220 33236 10276 33246
rect 10220 33142 10276 33180
rect 10556 33012 10612 34188
rect 10668 33236 10724 33246
rect 10780 33236 10836 34636
rect 10724 33180 10836 33236
rect 11116 34018 11172 34030
rect 11116 33966 11118 34018
rect 11170 33966 11172 34018
rect 10668 33142 10724 33180
rect 10892 33122 10948 33134
rect 10892 33070 10894 33122
rect 10946 33070 10948 33122
rect 10892 33012 10948 33070
rect 10556 32956 10948 33012
rect 10892 32900 10948 32956
rect 10892 32834 10948 32844
rect 11004 33122 11060 33134
rect 11004 33070 11006 33122
rect 11058 33070 11060 33122
rect 9996 32674 10052 32732
rect 11004 32786 11060 33070
rect 11004 32734 11006 32786
rect 11058 32734 11060 32786
rect 11004 32722 11060 32734
rect 9996 32622 9998 32674
rect 10050 32622 10052 32674
rect 9996 32610 10052 32622
rect 10108 32676 10164 32686
rect 10108 32582 10164 32620
rect 10332 32564 10388 32574
rect 10780 32564 10836 32574
rect 10332 32562 10836 32564
rect 10332 32510 10334 32562
rect 10386 32510 10782 32562
rect 10834 32510 10836 32562
rect 10332 32508 10836 32510
rect 10332 32498 10388 32508
rect 10780 32498 10836 32508
rect 10220 30996 10276 31006
rect 11116 30996 11172 33966
rect 11228 32786 11284 34972
rect 11452 34692 11508 34702
rect 11564 34692 11620 35420
rect 11676 35140 11732 35150
rect 11676 34802 11732 35084
rect 11676 34750 11678 34802
rect 11730 34750 11732 34802
rect 11676 34738 11732 34750
rect 11788 34916 11844 34926
rect 11788 34802 11844 34860
rect 11788 34750 11790 34802
rect 11842 34750 11844 34802
rect 11788 34738 11844 34750
rect 11452 34690 11620 34692
rect 11452 34638 11454 34690
rect 11506 34638 11620 34690
rect 11452 34636 11620 34638
rect 11452 34626 11508 34636
rect 11900 34580 11956 35644
rect 12124 35308 12180 37884
rect 12348 37604 12404 37998
rect 12348 37538 12404 37548
rect 12460 37938 12516 37950
rect 12460 37886 12462 37938
rect 12514 37886 12516 37938
rect 12348 37380 12404 37390
rect 12348 36484 12404 37324
rect 12460 37266 12516 37886
rect 12460 37214 12462 37266
rect 12514 37214 12516 37266
rect 12460 37202 12516 37214
rect 12348 36482 12516 36484
rect 12348 36430 12350 36482
rect 12402 36430 12516 36482
rect 12348 36428 12516 36430
rect 12348 36418 12404 36428
rect 12012 35252 12180 35308
rect 12012 35028 12068 35252
rect 12012 34802 12068 34972
rect 12012 34750 12014 34802
rect 12066 34750 12068 34802
rect 12012 34738 12068 34750
rect 12124 35140 12180 35150
rect 12124 34804 12180 35084
rect 12236 35028 12292 35038
rect 12236 34934 12292 34972
rect 11900 34524 12068 34580
rect 11788 33122 11844 33134
rect 11788 33070 11790 33122
rect 11842 33070 11844 33122
rect 11788 32788 11844 33070
rect 11228 32734 11230 32786
rect 11282 32734 11284 32786
rect 11228 32722 11284 32734
rect 11452 32732 11844 32788
rect 12012 32788 12068 34524
rect 12124 33234 12180 34748
rect 12460 33348 12516 36428
rect 12572 36482 12628 38668
rect 12572 36430 12574 36482
rect 12626 36430 12628 36482
rect 12572 36418 12628 36430
rect 12684 35586 12740 38780
rect 12908 37604 12964 39228
rect 13244 38724 13300 39452
rect 14028 39508 14084 39518
rect 14028 39414 14084 39452
rect 14700 39506 14756 39518
rect 14700 39454 14702 39506
rect 14754 39454 14756 39506
rect 13692 39394 13748 39406
rect 13692 39342 13694 39394
rect 13746 39342 13748 39394
rect 13692 39284 13748 39342
rect 13692 39218 13748 39228
rect 14364 39394 14420 39406
rect 14364 39342 14366 39394
rect 14418 39342 14420 39394
rect 13020 38668 13300 38724
rect 13356 38834 13412 38846
rect 13356 38782 13358 38834
rect 13410 38782 13412 38834
rect 13020 38612 13188 38668
rect 13020 37604 13076 37614
rect 12908 37548 13020 37604
rect 13020 37538 13076 37548
rect 12908 37156 12964 37166
rect 12796 36484 12852 36494
rect 12796 36390 12852 36428
rect 12908 36482 12964 37100
rect 12908 36430 12910 36482
rect 12962 36430 12964 36482
rect 12908 36418 12964 36430
rect 12684 35534 12686 35586
rect 12738 35534 12740 35586
rect 12684 35522 12740 35534
rect 13132 35364 13188 38612
rect 13244 38500 13300 38510
rect 13244 37266 13300 38444
rect 13356 38164 13412 38782
rect 13356 38098 13412 38108
rect 13580 38724 13636 38734
rect 13580 38388 13636 38668
rect 13244 37214 13246 37266
rect 13298 37214 13300 37266
rect 13244 37202 13300 37214
rect 13468 37266 13524 37278
rect 13468 37214 13470 37266
rect 13522 37214 13524 37266
rect 13356 37042 13412 37054
rect 13356 36990 13358 37042
rect 13410 36990 13412 37042
rect 13356 36372 13412 36990
rect 13468 37044 13524 37214
rect 13468 36978 13524 36988
rect 13580 36932 13636 38332
rect 14140 38500 14196 38510
rect 14140 38162 14196 38444
rect 14140 38110 14142 38162
rect 14194 38110 14196 38162
rect 14140 38098 14196 38110
rect 13692 38052 13748 38062
rect 13692 37380 13748 37996
rect 14364 38050 14420 39342
rect 14588 39396 14644 39406
rect 14588 39302 14644 39340
rect 14700 39060 14756 39454
rect 14700 38994 14756 39004
rect 14924 38836 14980 39676
rect 15820 39060 15876 40350
rect 16268 40404 16324 40414
rect 16268 40310 16324 40348
rect 15820 38994 15876 39004
rect 14812 38164 14868 38174
rect 14812 38070 14868 38108
rect 14364 37998 14366 38050
rect 14418 37998 14420 38050
rect 14364 37986 14420 37998
rect 14700 37828 14756 37838
rect 14924 37828 14980 38780
rect 15708 38724 15764 38734
rect 16044 38724 16100 38734
rect 15708 38722 16100 38724
rect 15708 38670 15710 38722
rect 15762 38670 16046 38722
rect 16098 38670 16100 38722
rect 15708 38668 16100 38670
rect 15708 38658 15764 38668
rect 16044 38658 16100 38668
rect 16156 38722 16212 38734
rect 16156 38670 16158 38722
rect 16210 38670 16212 38722
rect 15484 37828 15540 37838
rect 14700 37734 14756 37772
rect 14812 37826 14980 37828
rect 14812 37774 14926 37826
rect 14978 37774 14980 37826
rect 14812 37772 14980 37774
rect 13692 37314 13748 37324
rect 13916 37380 13972 37390
rect 13916 37286 13972 37324
rect 14140 37268 14196 37278
rect 14140 37174 14196 37212
rect 13692 37156 13748 37166
rect 14700 37156 14756 37166
rect 13692 37062 13748 37100
rect 14588 37154 14756 37156
rect 14588 37102 14702 37154
rect 14754 37102 14756 37154
rect 14588 37100 14756 37102
rect 13580 36876 14196 36932
rect 14028 36484 14084 36494
rect 14028 36390 14084 36428
rect 13356 36306 13412 36316
rect 13692 36260 13748 36270
rect 13692 35588 13748 36204
rect 13916 35924 13972 35934
rect 14140 35924 14196 36876
rect 14364 36596 14420 36606
rect 14252 36372 14308 36382
rect 14252 36278 14308 36316
rect 14252 35924 14308 35934
rect 14140 35922 14308 35924
rect 14140 35870 14254 35922
rect 14306 35870 14308 35922
rect 14140 35868 14308 35870
rect 13916 35700 13972 35868
rect 14252 35858 14308 35868
rect 13916 35698 14196 35700
rect 13916 35646 13918 35698
rect 13970 35646 14196 35698
rect 13916 35644 14196 35646
rect 13916 35634 13972 35644
rect 12572 35308 13188 35364
rect 13244 35532 13748 35588
rect 12572 34802 12628 35308
rect 12572 34750 12574 34802
rect 12626 34750 12628 34802
rect 12572 34738 12628 34750
rect 12908 34804 12964 34814
rect 13244 34804 13300 35532
rect 13468 35364 13524 35374
rect 12908 34802 13300 34804
rect 12908 34750 12910 34802
rect 12962 34750 13300 34802
rect 12908 34748 13300 34750
rect 13356 35028 13412 35038
rect 12908 34738 12964 34748
rect 12124 33182 12126 33234
rect 12178 33182 12180 33234
rect 12124 33170 12180 33182
rect 12236 33292 12852 33348
rect 11452 32562 11508 32732
rect 12012 32722 12068 32732
rect 12124 32788 12180 32798
rect 12236 32788 12292 33292
rect 12460 33122 12516 33134
rect 12460 33070 12462 33122
rect 12514 33070 12516 33122
rect 12460 33012 12516 33070
rect 12460 32946 12516 32956
rect 12124 32786 12292 32788
rect 12124 32734 12126 32786
rect 12178 32734 12292 32786
rect 12124 32732 12292 32734
rect 12572 32788 12628 32798
rect 12572 32786 12740 32788
rect 12572 32734 12574 32786
rect 12626 32734 12740 32786
rect 12572 32732 12740 32734
rect 12124 32722 12180 32732
rect 12572 32722 12628 32732
rect 12460 32676 12516 32686
rect 11452 32510 11454 32562
rect 11506 32510 11508 32562
rect 11452 31444 11508 32510
rect 11564 32564 11620 32574
rect 12236 32564 12292 32574
rect 11564 32470 11620 32508
rect 11676 32562 12292 32564
rect 11676 32510 12238 32562
rect 12290 32510 12292 32562
rect 11676 32508 12292 32510
rect 12460 32564 12516 32620
rect 12684 32676 12740 32732
rect 12796 32676 12852 33292
rect 12908 33122 12964 33134
rect 12908 33070 12910 33122
rect 12962 33070 12964 33122
rect 12908 33012 12964 33070
rect 12908 32946 12964 32956
rect 12908 32676 12964 32686
rect 12796 32674 12964 32676
rect 12796 32622 12910 32674
rect 12962 32622 12964 32674
rect 12796 32620 12964 32622
rect 12684 32610 12740 32620
rect 12908 32610 12964 32620
rect 12572 32564 12628 32574
rect 12460 32562 12628 32564
rect 12460 32510 12574 32562
rect 12626 32510 12628 32562
rect 12460 32508 12628 32510
rect 11676 31890 11732 32508
rect 12236 32498 12292 32508
rect 12572 32498 12628 32508
rect 11676 31838 11678 31890
rect 11730 31838 11732 31890
rect 11676 31826 11732 31838
rect 11564 31668 11620 31678
rect 11564 31574 11620 31612
rect 11900 31668 11956 31678
rect 11900 31574 11956 31612
rect 12124 31666 12180 31678
rect 12124 31614 12126 31666
rect 12178 31614 12180 31666
rect 12124 31556 12180 31614
rect 12684 31556 12740 31566
rect 12124 31554 12740 31556
rect 12124 31502 12686 31554
rect 12738 31502 12740 31554
rect 12124 31500 12740 31502
rect 11452 31388 11844 31444
rect 10220 30994 10388 30996
rect 10220 30942 10222 30994
rect 10274 30942 10388 30994
rect 10220 30940 10388 30942
rect 10220 30930 10276 30940
rect 10332 30098 10388 30940
rect 10892 30940 11116 30996
rect 10668 30212 10724 30222
rect 10668 30118 10724 30156
rect 10332 30046 10334 30098
rect 10386 30046 10388 30098
rect 10332 30034 10388 30046
rect 9884 29372 10052 29428
rect 9884 28756 9940 28794
rect 9884 28690 9940 28700
rect 9772 28644 9828 28654
rect 9772 28550 9828 28588
rect 9548 28252 9828 28308
rect 8988 28030 8990 28082
rect 9042 28030 9044 28082
rect 8988 28018 9044 28030
rect 9660 28084 9716 28094
rect 9660 27990 9716 28028
rect 9772 27972 9828 28252
rect 9996 28196 10052 29372
rect 10332 28532 10388 28542
rect 9996 28140 10276 28196
rect 9772 27970 10052 27972
rect 9772 27918 9774 27970
rect 9826 27918 10052 27970
rect 9772 27916 10052 27918
rect 9772 27906 9828 27916
rect 9436 27860 9492 27870
rect 8876 27858 9492 27860
rect 8876 27806 9438 27858
rect 9490 27806 9492 27858
rect 8876 27804 9492 27806
rect 9436 27794 9492 27804
rect 8204 27122 8260 27132
rect 9212 27524 9268 27534
rect 8092 27076 8148 27086
rect 8092 26982 8148 27020
rect 8764 27074 8820 27086
rect 8764 27022 8766 27074
rect 8818 27022 8820 27074
rect 8764 26292 8820 27022
rect 8876 26964 8932 26974
rect 8876 26514 8932 26908
rect 8876 26462 8878 26514
rect 8930 26462 8932 26514
rect 8876 26450 8932 26462
rect 8988 26962 9044 26974
rect 8988 26910 8990 26962
rect 9042 26910 9044 26962
rect 8652 26066 8708 26078
rect 8652 26014 8654 26066
rect 8706 26014 8708 26066
rect 8652 25730 8708 26014
rect 8652 25678 8654 25730
rect 8706 25678 8708 25730
rect 8316 25506 8372 25518
rect 8316 25454 8318 25506
rect 8370 25454 8372 25506
rect 7980 24722 8036 24734
rect 7980 24670 7982 24722
rect 8034 24670 8036 24722
rect 7980 24052 8036 24670
rect 8316 24612 8372 25454
rect 8540 25282 8596 25294
rect 8540 25230 8542 25282
rect 8594 25230 8596 25282
rect 8540 24948 8596 25230
rect 8652 25284 8708 25678
rect 8652 25218 8708 25228
rect 8316 24546 8372 24556
rect 8428 24892 8596 24948
rect 8092 24052 8148 24062
rect 7980 24050 8148 24052
rect 7980 23998 8094 24050
rect 8146 23998 8148 24050
rect 7980 23996 8148 23998
rect 8092 23986 8148 23996
rect 7868 23886 7870 23938
rect 7922 23886 7924 23938
rect 7868 23874 7924 23886
rect 8204 23938 8260 23950
rect 8204 23886 8206 23938
rect 8258 23886 8260 23938
rect 7644 23660 8036 23716
rect 7980 23378 8036 23660
rect 7980 23326 7982 23378
rect 8034 23326 8036 23378
rect 7980 23314 8036 23326
rect 6188 22082 6244 22092
rect 6300 23268 6356 23278
rect 6300 22482 6356 23212
rect 6412 23266 6468 23278
rect 6412 23214 6414 23266
rect 6466 23214 6468 23266
rect 6412 23156 6468 23214
rect 6412 23090 6468 23100
rect 8204 23154 8260 23886
rect 8428 23938 8484 24892
rect 8540 24724 8596 24734
rect 8764 24724 8820 26236
rect 8988 26178 9044 26910
rect 9212 26908 9268 27468
rect 9324 27412 9380 27422
rect 9324 27074 9380 27356
rect 9996 27188 10052 27916
rect 10108 27970 10164 27982
rect 10108 27918 10110 27970
rect 10162 27918 10164 27970
rect 10108 27524 10164 27918
rect 10108 27300 10164 27468
rect 10108 27234 10164 27244
rect 9884 27186 10052 27188
rect 9884 27134 9998 27186
rect 10050 27134 10052 27186
rect 9884 27132 10052 27134
rect 9324 27022 9326 27074
rect 9378 27022 9380 27074
rect 9324 27010 9380 27022
rect 9436 27076 9492 27086
rect 9436 26982 9492 27020
rect 9548 26962 9604 26974
rect 9548 26910 9550 26962
rect 9602 26910 9604 26962
rect 9548 26908 9604 26910
rect 9212 26852 9604 26908
rect 9548 26404 9604 26414
rect 8988 26126 8990 26178
rect 9042 26126 9044 26178
rect 8988 26114 9044 26126
rect 9436 26348 9548 26404
rect 9212 25508 9268 25518
rect 9212 25414 9268 25452
rect 9436 24946 9492 26348
rect 9548 26338 9604 26348
rect 9660 26180 9716 26190
rect 9436 24894 9438 24946
rect 9490 24894 9492 24946
rect 9436 24882 9492 24894
rect 9548 26178 9716 26180
rect 9548 26126 9662 26178
rect 9714 26126 9716 26178
rect 9548 26124 9716 26126
rect 9100 24836 9156 24846
rect 8988 24724 9044 24734
rect 8764 24668 8988 24724
rect 8540 24630 8596 24668
rect 8428 23886 8430 23938
rect 8482 23886 8484 23938
rect 8428 23874 8484 23886
rect 8764 23716 8820 23726
rect 8204 23102 8206 23154
rect 8258 23102 8260 23154
rect 8092 23042 8148 23054
rect 8092 22990 8094 23042
rect 8146 22990 8148 23042
rect 8092 22708 8148 22990
rect 6300 22430 6302 22482
rect 6354 22430 6356 22482
rect 5628 21588 5684 21598
rect 5516 21586 5684 21588
rect 5516 21534 5630 21586
rect 5682 21534 5684 21586
rect 5516 21532 5684 21534
rect 5628 21522 5684 21532
rect 6300 21586 6356 22430
rect 7308 22652 8148 22708
rect 6524 22372 6580 22382
rect 6524 22278 6580 22316
rect 7308 22370 7364 22652
rect 8204 22596 8260 23102
rect 8652 23714 8820 23716
rect 8652 23662 8766 23714
rect 8818 23662 8820 23714
rect 8652 23660 8820 23662
rect 8652 23154 8708 23660
rect 8764 23650 8820 23660
rect 8652 23102 8654 23154
rect 8706 23102 8708 23154
rect 8652 23090 8708 23102
rect 8204 22530 8260 22540
rect 7308 22318 7310 22370
rect 7362 22318 7364 22370
rect 7308 22306 7364 22318
rect 6972 22148 7028 22158
rect 6300 21534 6302 21586
rect 6354 21534 6356 21586
rect 5292 21364 5348 21374
rect 5292 21270 5348 21308
rect 5068 20862 5070 20914
rect 5122 20862 5124 20914
rect 2604 20692 2660 20702
rect 2492 20690 2660 20692
rect 2492 20638 2606 20690
rect 2658 20638 2660 20690
rect 2492 20636 2660 20638
rect 2604 20626 2660 20636
rect 5068 20132 5124 20862
rect 6300 20804 6356 21534
rect 6412 21698 6468 21710
rect 6412 21646 6414 21698
rect 6466 21646 6468 21698
rect 6412 21588 6468 21646
rect 6412 21026 6468 21532
rect 6972 21476 7028 22092
rect 8876 21588 8932 24668
rect 8988 24630 9044 24668
rect 9100 24276 9156 24780
rect 9548 24724 9604 26124
rect 9660 26114 9716 26124
rect 9884 26180 9940 27132
rect 9996 27122 10052 27132
rect 9996 26964 10052 26974
rect 10220 26908 10276 28140
rect 10332 27858 10388 28476
rect 10668 28530 10724 28542
rect 10668 28478 10670 28530
rect 10722 28478 10724 28530
rect 10444 28420 10500 28430
rect 10668 28420 10724 28478
rect 10444 28418 10724 28420
rect 10444 28366 10446 28418
rect 10498 28366 10724 28418
rect 10444 28364 10724 28366
rect 10444 28354 10500 28364
rect 10332 27806 10334 27858
rect 10386 27806 10388 27858
rect 10332 27794 10388 27806
rect 9996 26402 10052 26908
rect 9996 26350 9998 26402
rect 10050 26350 10052 26402
rect 9996 26338 10052 26350
rect 10108 26852 10276 26908
rect 10668 26908 10724 28364
rect 10780 28418 10836 28430
rect 10780 28366 10782 28418
rect 10834 28366 10836 28418
rect 10780 28084 10836 28366
rect 10780 28018 10836 28028
rect 10892 27858 10948 30940
rect 11116 30930 11172 30940
rect 11676 30212 11732 30222
rect 11676 30118 11732 30156
rect 11004 28644 11060 28654
rect 11004 28642 11396 28644
rect 11004 28590 11006 28642
rect 11058 28590 11396 28642
rect 11004 28588 11396 28590
rect 11004 28578 11060 28588
rect 10892 27806 10894 27858
rect 10946 27806 10948 27858
rect 10892 27794 10948 27806
rect 10780 27412 10836 27422
rect 10780 27074 10836 27356
rect 10780 27022 10782 27074
rect 10834 27022 10836 27074
rect 10780 27010 10836 27022
rect 11116 27186 11172 27198
rect 11116 27134 11118 27186
rect 11170 27134 11172 27186
rect 11116 26964 11172 27134
rect 11340 27076 11396 28588
rect 11564 28418 11620 28430
rect 11564 28366 11566 28418
rect 11618 28366 11620 28418
rect 11452 27860 11508 27870
rect 11564 27860 11620 28366
rect 11452 27858 11620 27860
rect 11452 27806 11454 27858
rect 11506 27806 11620 27858
rect 11452 27804 11620 27806
rect 11452 27794 11508 27804
rect 11676 27186 11732 27198
rect 11676 27134 11678 27186
rect 11730 27134 11732 27186
rect 11564 27076 11620 27086
rect 11340 27074 11620 27076
rect 11340 27022 11566 27074
rect 11618 27022 11620 27074
rect 11340 27020 11620 27022
rect 11564 27010 11620 27020
rect 10668 26852 10836 26908
rect 10108 26404 10164 26852
rect 10108 26310 10164 26348
rect 10668 26404 10724 26414
rect 10668 26310 10724 26348
rect 10332 26292 10388 26302
rect 10332 26290 10500 26292
rect 10332 26238 10334 26290
rect 10386 26238 10500 26290
rect 10332 26236 10500 26238
rect 10332 26226 10388 26236
rect 9884 26114 9940 26124
rect 10444 26066 10500 26236
rect 10444 26014 10446 26066
rect 10498 26014 10500 26066
rect 10444 26002 10500 26014
rect 9660 25956 9716 25966
rect 9660 25618 9716 25900
rect 9660 25566 9662 25618
rect 9714 25566 9716 25618
rect 9660 25554 9716 25566
rect 10332 25506 10388 25518
rect 10332 25454 10334 25506
rect 10386 25454 10388 25506
rect 9884 25394 9940 25406
rect 9884 25342 9886 25394
rect 9938 25342 9940 25394
rect 9884 25060 9940 25342
rect 9884 24994 9940 25004
rect 9996 25394 10052 25406
rect 9996 25342 9998 25394
rect 10050 25342 10052 25394
rect 9884 24836 9940 24846
rect 9884 24742 9940 24780
rect 9660 24724 9716 24734
rect 9548 24668 9660 24724
rect 9660 24658 9716 24668
rect 9772 24722 9828 24734
rect 9772 24670 9774 24722
rect 9826 24670 9828 24722
rect 8988 24220 9156 24276
rect 9436 24500 9492 24510
rect 8988 23828 9044 24220
rect 9436 23938 9492 24444
rect 9436 23886 9438 23938
rect 9490 23886 9492 23938
rect 9436 23874 9492 23886
rect 9548 24498 9604 24510
rect 9548 24446 9550 24498
rect 9602 24446 9604 24498
rect 8988 23734 9044 23772
rect 9100 23828 9156 23838
rect 9324 23828 9380 23838
rect 9100 23826 9324 23828
rect 9100 23774 9102 23826
rect 9154 23774 9324 23826
rect 9100 23772 9324 23774
rect 9100 23762 9156 23772
rect 9324 23762 9380 23772
rect 9548 23826 9604 24446
rect 9772 24276 9828 24670
rect 9884 24500 9940 24510
rect 9996 24500 10052 25342
rect 10332 25060 10388 25454
rect 10780 25284 10836 26852
rect 11116 26178 11172 26908
rect 11676 26908 11732 27134
rect 11788 27076 11844 31388
rect 12012 30436 12068 30446
rect 12012 30342 12068 30380
rect 12012 29204 12068 29214
rect 11900 29148 12012 29204
rect 11900 28642 11956 29148
rect 12012 29138 12068 29148
rect 11900 28590 11902 28642
rect 11954 28590 11956 28642
rect 11900 28578 11956 28590
rect 12012 27076 12068 27086
rect 11788 27020 12012 27076
rect 12012 26982 12068 27020
rect 11676 26852 11844 26908
rect 11116 26126 11118 26178
rect 11170 26126 11172 26178
rect 10892 26066 10948 26078
rect 10892 26014 10894 26066
rect 10946 26014 10948 26066
rect 10892 25506 10948 26014
rect 11116 25956 11172 26126
rect 11116 25890 11172 25900
rect 10892 25454 10894 25506
rect 10946 25454 10948 25506
rect 10892 25442 10948 25454
rect 11340 25394 11396 25406
rect 11340 25342 11342 25394
rect 11394 25342 11396 25394
rect 10780 25228 11172 25284
rect 9884 24498 10052 24500
rect 9884 24446 9886 24498
rect 9938 24446 10052 24498
rect 9884 24444 10052 24446
rect 10220 25004 10948 25060
rect 9884 24434 9940 24444
rect 9548 23774 9550 23826
rect 9602 23774 9604 23826
rect 9212 23604 9268 23614
rect 9100 23380 9156 23390
rect 9100 23286 9156 23324
rect 9212 22596 9268 23548
rect 9548 23380 9604 23774
rect 9548 23314 9604 23324
rect 9660 24220 9772 24276
rect 9212 22530 9268 22540
rect 9660 22484 9716 24220
rect 9772 24210 9828 24220
rect 9996 23940 10052 23950
rect 9996 23846 10052 23884
rect 9772 23714 9828 23726
rect 9772 23662 9774 23714
rect 9826 23662 9828 23714
rect 9772 23268 9828 23662
rect 10108 23714 10164 23726
rect 10108 23662 10110 23714
rect 10162 23662 10164 23714
rect 10108 23380 10164 23662
rect 10220 23716 10276 25004
rect 10892 24946 10948 25004
rect 10892 24894 10894 24946
rect 10946 24894 10948 24946
rect 10892 24882 10948 24894
rect 11004 24948 11060 24958
rect 10556 24836 10612 24846
rect 10444 24610 10500 24622
rect 10444 24558 10446 24610
rect 10498 24558 10500 24610
rect 10332 24498 10388 24510
rect 10332 24446 10334 24498
rect 10386 24446 10388 24498
rect 10332 23938 10388 24446
rect 10444 24276 10500 24558
rect 10444 24210 10500 24220
rect 10332 23886 10334 23938
rect 10386 23886 10388 23938
rect 10332 23874 10388 23886
rect 10556 23938 10612 24780
rect 11004 24498 11060 24892
rect 11004 24446 11006 24498
rect 11058 24446 11060 24498
rect 11004 24434 11060 24446
rect 10556 23886 10558 23938
rect 10610 23886 10612 23938
rect 10556 23874 10612 23886
rect 10780 23938 10836 23950
rect 10780 23886 10782 23938
rect 10834 23886 10836 23938
rect 10220 23660 10388 23716
rect 9772 23202 9828 23212
rect 9996 23324 10164 23380
rect 10220 23492 10276 23502
rect 10220 23378 10276 23436
rect 10220 23326 10222 23378
rect 10274 23326 10276 23378
rect 9548 22428 9716 22484
rect 9772 23044 9828 23054
rect 9996 23044 10052 23324
rect 10220 23314 10276 23326
rect 10108 23156 10164 23166
rect 10108 23062 10164 23100
rect 9772 23042 10052 23044
rect 9772 22990 9774 23042
rect 9826 22990 10052 23042
rect 9772 22988 10052 22990
rect 9548 21924 9604 22428
rect 9660 22260 9716 22270
rect 9660 22166 9716 22204
rect 9100 21868 9604 21924
rect 9772 21924 9828 22988
rect 9996 22596 10052 22606
rect 9996 22502 10052 22540
rect 10220 22484 10276 22494
rect 10108 22260 10164 22270
rect 10108 22166 10164 22204
rect 9884 21924 9940 21934
rect 9772 21868 9884 21924
rect 9100 21810 9156 21868
rect 9100 21758 9102 21810
rect 9154 21758 9156 21810
rect 9100 21746 9156 21758
rect 9548 21700 9604 21868
rect 9660 21700 9716 21710
rect 9548 21698 9716 21700
rect 9548 21646 9662 21698
rect 9714 21646 9716 21698
rect 9548 21644 9716 21646
rect 9660 21634 9716 21644
rect 9772 21588 9828 21598
rect 8876 21532 9380 21588
rect 6972 21382 7028 21420
rect 7308 21476 7364 21486
rect 6412 20974 6414 21026
rect 6466 20974 6468 21026
rect 6412 20962 6468 20974
rect 6300 20748 6692 20804
rect 6636 20690 6692 20748
rect 6636 20638 6638 20690
rect 6690 20638 6692 20690
rect 6636 20626 6692 20638
rect 6972 20690 7028 20702
rect 6972 20638 6974 20690
rect 7026 20638 7028 20690
rect 6076 20580 6132 20590
rect 5964 20578 6132 20580
rect 5964 20526 6078 20578
rect 6130 20526 6132 20578
rect 5964 20524 6132 20526
rect 5964 20356 6020 20524
rect 6076 20514 6132 20524
rect 5068 20066 5124 20076
rect 5404 20300 6020 20356
rect 5404 20018 5460 20300
rect 5404 19966 5406 20018
rect 5458 19966 5460 20018
rect 5404 19954 5460 19966
rect 5628 20130 5684 20142
rect 5628 20078 5630 20130
rect 5682 20078 5684 20130
rect 5628 20020 5684 20078
rect 5852 20132 5908 20142
rect 5852 20020 5908 20076
rect 6972 20132 7028 20638
rect 5628 19954 5684 19964
rect 5740 20018 5908 20020
rect 5740 19966 5854 20018
rect 5906 19966 5908 20018
rect 5740 19964 5908 19966
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4396 19460 4452 19470
rect 2268 19234 2324 19246
rect 2268 19182 2270 19234
rect 2322 19182 2324 19234
rect 2268 18674 2324 19182
rect 2268 18622 2270 18674
rect 2322 18622 2324 18674
rect 2268 18610 2324 18622
rect 4172 19012 4228 19022
rect 2604 18452 2660 18462
rect 2604 18358 2660 18396
rect 4060 18452 4116 18462
rect 4060 18358 4116 18396
rect 4172 17890 4228 18956
rect 4396 18450 4452 19404
rect 5740 19346 5796 19964
rect 5852 19954 5908 19964
rect 6524 20020 6580 20030
rect 6524 19926 6580 19964
rect 6972 19460 7028 20076
rect 6972 19394 7028 19404
rect 7308 19348 7364 21420
rect 8988 20916 9044 20926
rect 8988 20822 9044 20860
rect 9324 20914 9380 21532
rect 9772 21494 9828 21532
rect 9324 20862 9326 20914
rect 9378 20862 9380 20914
rect 9324 20850 9380 20862
rect 8204 20804 8260 20814
rect 5740 19294 5742 19346
rect 5794 19294 5796 19346
rect 4732 19012 4788 19022
rect 4732 18918 4788 18956
rect 5180 19012 5236 19022
rect 5180 18562 5236 18956
rect 5180 18510 5182 18562
rect 5234 18510 5236 18562
rect 5180 18498 5236 18510
rect 4396 18398 4398 18450
rect 4450 18398 4452 18450
rect 4396 18386 4452 18398
rect 4844 18450 4900 18462
rect 4844 18398 4846 18450
rect 4898 18398 4900 18450
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4172 17838 4174 17890
rect 4226 17838 4228 17890
rect 4172 17826 4228 17838
rect 4620 17668 4676 17678
rect 4844 17668 4900 18398
rect 4620 17666 4900 17668
rect 4620 17614 4622 17666
rect 4674 17614 4900 17666
rect 4620 17612 4900 17614
rect 4956 17668 5012 17678
rect 2492 17556 2548 17566
rect 2492 17462 2548 17500
rect 3836 17556 3892 17566
rect 3836 17462 3892 17500
rect 4620 17556 4676 17612
rect 4956 17556 5012 17612
rect 2156 17442 2212 17454
rect 2156 17390 2158 17442
rect 2210 17390 2212 17442
rect 2156 16884 2212 17390
rect 4172 16996 4228 17006
rect 2268 16884 2324 16894
rect 2156 16882 2324 16884
rect 2156 16830 2270 16882
rect 2322 16830 2324 16882
rect 2156 16828 2324 16830
rect 2268 16818 2324 16828
rect 4172 16322 4228 16940
rect 4620 16884 4676 17500
rect 4732 17554 5012 17556
rect 4732 17502 4958 17554
rect 5010 17502 5012 17554
rect 4732 17500 5012 17502
rect 4732 17106 4788 17500
rect 4956 17490 5012 17500
rect 4732 17054 4734 17106
rect 4786 17054 4788 17106
rect 4732 17042 4788 17054
rect 4956 16884 5012 16894
rect 4620 16828 4900 16884
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4172 16270 4174 16322
rect 4226 16270 4228 16322
rect 4172 16258 4228 16270
rect 4844 16098 4900 16828
rect 4844 16046 4846 16098
rect 4898 16046 4900 16098
rect 4844 16034 4900 16046
rect 5740 16884 5796 19294
rect 7084 19346 7364 19348
rect 7084 19294 7310 19346
rect 7362 19294 7364 19346
rect 7084 19292 7364 19294
rect 6860 19236 6916 19246
rect 7084 19236 7140 19292
rect 7308 19282 7364 19292
rect 7532 20580 7588 20590
rect 6860 19234 7140 19236
rect 6860 19182 6862 19234
rect 6914 19182 7140 19234
rect 6860 19180 7140 19182
rect 6860 19170 6916 19180
rect 6300 19122 6356 19134
rect 6300 19070 6302 19122
rect 6354 19070 6356 19122
rect 6300 18564 6356 19070
rect 6076 18508 6356 18564
rect 6748 18562 6804 18574
rect 6748 18510 6750 18562
rect 6802 18510 6804 18562
rect 6076 17556 6132 18508
rect 6412 18452 6468 18462
rect 6188 18450 6468 18452
rect 6188 18398 6414 18450
rect 6466 18398 6468 18450
rect 6188 18396 6468 18398
rect 6188 17890 6244 18396
rect 6412 18386 6468 18396
rect 6188 17838 6190 17890
rect 6242 17838 6244 17890
rect 6188 17826 6244 17838
rect 6748 17780 6804 18510
rect 6636 17724 6804 17780
rect 6524 17668 6580 17678
rect 6524 17574 6580 17612
rect 6076 17490 6132 17500
rect 5852 16884 5908 16894
rect 5740 16882 6132 16884
rect 5740 16830 5854 16882
rect 5906 16830 6132 16882
rect 5740 16828 6132 16830
rect 4956 15986 5012 16828
rect 5852 16818 5908 16828
rect 4956 15934 4958 15986
rect 5010 15934 5012 15986
rect 2492 15876 2548 15886
rect 2156 15426 2212 15438
rect 2156 15374 2158 15426
rect 2210 15374 2212 15426
rect 2156 14532 2212 15374
rect 2492 15426 2548 15820
rect 3836 15876 3892 15886
rect 3836 15782 3892 15820
rect 2492 15374 2494 15426
rect 2546 15374 2548 15426
rect 2492 15362 2548 15374
rect 4284 15426 4340 15438
rect 4284 15374 4286 15426
rect 4338 15374 4340 15426
rect 4284 15148 4340 15374
rect 4172 15092 4340 15148
rect 4620 15314 4676 15326
rect 4620 15262 4622 15314
rect 4674 15262 4676 15314
rect 4620 15092 4676 15262
rect 2268 14532 2324 14542
rect 2156 14530 2324 14532
rect 2156 14478 2270 14530
rect 2322 14478 2324 14530
rect 2156 14476 2324 14478
rect 2268 14466 2324 14476
rect 3612 14308 3668 14318
rect 3612 13748 3668 14252
rect 3612 13654 3668 13692
rect 4172 13746 4228 15092
rect 4620 15026 4676 15036
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4172 13694 4174 13746
rect 4226 13694 4228 13746
rect 4172 13682 4228 13694
rect 4732 14308 4788 14318
rect 4956 14308 5012 15934
rect 5180 16770 5236 16782
rect 5180 16718 5182 16770
rect 5234 16718 5236 16770
rect 4732 14306 5012 14308
rect 4732 14254 4734 14306
rect 4786 14254 5012 14306
rect 4732 14252 5012 14254
rect 5068 15540 5124 15550
rect 5180 15540 5236 16718
rect 5068 15538 5236 15540
rect 5068 15486 5070 15538
rect 5122 15486 5236 15538
rect 5068 15484 5236 15486
rect 5068 14308 5124 15484
rect 5740 15092 5796 15102
rect 4732 13524 4788 14252
rect 5068 14242 5124 14252
rect 5180 14756 5236 14766
rect 5180 13636 5236 14700
rect 5740 14754 5796 15036
rect 6076 15092 6132 16828
rect 6636 16882 6692 17724
rect 6748 17556 6804 17566
rect 6748 17462 6804 17500
rect 7084 17554 7140 17566
rect 7084 17502 7086 17554
rect 7138 17502 7140 17554
rect 7084 16996 7140 17502
rect 7084 16930 7140 16940
rect 6636 16830 6638 16882
rect 6690 16830 6692 16882
rect 6636 16818 6692 16830
rect 6076 15026 6132 15036
rect 7084 16100 7140 16110
rect 5740 14702 5742 14754
rect 5794 14702 5796 14754
rect 5740 14690 5796 14702
rect 6076 14756 6132 14766
rect 6076 14662 6132 14700
rect 6300 14418 6356 14430
rect 6300 14366 6302 14418
rect 6354 14366 6356 14418
rect 5964 14308 6020 14318
rect 4284 13468 4788 13524
rect 4844 13580 5236 13636
rect 5852 14252 5964 14308
rect 4172 12962 4228 12974
rect 4172 12910 4174 12962
rect 4226 12910 4228 12962
rect 2604 12852 2660 12862
rect 2604 12758 2660 12796
rect 3836 12852 3892 12862
rect 3836 12758 3892 12796
rect 2268 12738 2324 12750
rect 2268 12686 2270 12738
rect 2322 12686 2324 12738
rect 2268 12178 2324 12686
rect 2268 12126 2270 12178
rect 2322 12126 2324 12178
rect 2268 12114 2324 12126
rect 3612 12404 3668 12414
rect 2268 10612 2324 10622
rect 2156 10610 2324 10612
rect 2156 10558 2270 10610
rect 2322 10558 2324 10610
rect 2156 10556 2324 10558
rect 2156 9714 2212 10556
rect 2268 10546 2324 10556
rect 2156 9662 2158 9714
rect 2210 9662 2212 9714
rect 2156 9650 2212 9662
rect 2492 9716 2548 9726
rect 2492 9622 2548 9660
rect 3500 9716 3556 9726
rect 3500 9622 3556 9660
rect 1708 8206 1710 8258
rect 1762 8206 1764 8258
rect 1708 7700 1764 8206
rect 1708 5906 1764 7644
rect 1932 8372 2100 8428
rect 2492 8820 2548 8830
rect 1932 6804 1988 8372
rect 2268 8260 2324 8270
rect 2156 8258 2324 8260
rect 2156 8206 2270 8258
rect 2322 8206 2324 8258
rect 2156 8204 2324 8206
rect 2156 7698 2212 8204
rect 2268 8194 2324 8204
rect 2156 7646 2158 7698
rect 2210 7646 2212 7698
rect 2156 7634 2212 7646
rect 2492 7586 2548 8764
rect 3388 8820 3444 8830
rect 3388 8726 3444 8764
rect 2492 7534 2494 7586
rect 2546 7534 2548 7586
rect 2492 7522 2548 7534
rect 1708 5854 1710 5906
rect 1762 5854 1764 5906
rect 1708 5236 1764 5854
rect 1820 6748 1988 6804
rect 1820 5460 1876 6748
rect 3612 6692 3668 12348
rect 4172 12404 4228 12910
rect 4172 12338 4228 12348
rect 3836 10052 3892 10062
rect 4284 10052 4340 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4844 12850 4900 13580
rect 4956 13412 5012 13422
rect 4956 13188 5012 13356
rect 5740 13412 5796 13422
rect 4956 13132 5124 13188
rect 4956 12964 5012 12974
rect 4956 12870 5012 12908
rect 4844 12798 4846 12850
rect 4898 12798 4900 12850
rect 4732 12404 4788 12414
rect 4844 12404 4900 12798
rect 5068 12740 5124 13132
rect 5740 12964 5796 13356
rect 4732 12402 4900 12404
rect 4732 12350 4734 12402
rect 4786 12350 4900 12402
rect 4732 12348 4900 12350
rect 4956 12684 5124 12740
rect 5628 12962 5796 12964
rect 5628 12910 5742 12962
rect 5794 12910 5796 12962
rect 5628 12908 5796 12910
rect 4732 12338 4788 12348
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4956 11396 5012 12684
rect 5292 12404 5348 12414
rect 5292 12310 5348 12348
rect 4732 11340 5012 11396
rect 4732 10836 4788 11340
rect 4956 11172 5012 11182
rect 4732 10834 4900 10836
rect 4732 10782 4734 10834
rect 4786 10782 4900 10834
rect 4732 10780 4900 10782
rect 4732 10770 4788 10780
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4844 10052 4900 10780
rect 4956 10612 5012 11116
rect 5180 10612 5236 10622
rect 4956 10610 5236 10612
rect 4956 10558 5182 10610
rect 5234 10558 5236 10610
rect 4956 10556 5236 10558
rect 3836 10050 4340 10052
rect 3836 9998 3838 10050
rect 3890 9998 4340 10050
rect 3836 9996 4340 9998
rect 4396 9996 4900 10052
rect 3836 9986 3892 9996
rect 4396 9828 4452 9996
rect 3724 9772 4452 9828
rect 4508 9826 4564 9838
rect 4508 9774 4510 9826
rect 4562 9774 4564 9826
rect 3724 9042 3780 9772
rect 4396 9156 4452 9166
rect 3724 8990 3726 9042
rect 3778 8990 3780 9042
rect 3724 8978 3780 8990
rect 4284 9100 4396 9156
rect 4284 8484 4340 9100
rect 4396 9062 4452 9100
rect 4508 9042 4564 9774
rect 4620 9714 4676 9996
rect 4620 9662 4622 9714
rect 4674 9662 4676 9714
rect 4620 9650 4676 9662
rect 4508 8990 4510 9042
rect 4562 8990 4564 9042
rect 4508 8820 4564 8990
rect 5068 8932 5124 8942
rect 5180 8932 5236 10556
rect 5068 8930 5236 8932
rect 5068 8878 5070 8930
rect 5122 8878 5236 8930
rect 5068 8876 5236 8878
rect 5068 8866 5124 8876
rect 4508 8764 4900 8820
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 3948 8428 4788 8484
rect 3948 6914 4004 8428
rect 4732 8370 4788 8428
rect 4732 8318 4734 8370
rect 4786 8318 4788 8370
rect 4732 8306 4788 8318
rect 3948 6862 3950 6914
rect 4002 6862 4004 6914
rect 3948 6850 4004 6862
rect 4284 7700 4340 7710
rect 3612 6636 3780 6692
rect 1932 6580 1988 6590
rect 1932 6578 2436 6580
rect 1932 6526 1934 6578
rect 1986 6526 2436 6578
rect 1932 6524 2436 6526
rect 1932 6514 1988 6524
rect 2268 5908 2324 5918
rect 2156 5906 2324 5908
rect 2156 5854 2270 5906
rect 2322 5854 2324 5906
rect 2156 5852 2324 5854
rect 1820 5404 2100 5460
rect 1820 5236 1876 5246
rect 1708 5234 1876 5236
rect 1708 5182 1822 5234
rect 1874 5182 1876 5234
rect 1708 5180 1876 5182
rect 1708 4338 1764 5180
rect 1820 5170 1876 5180
rect 1708 4286 1710 4338
rect 1762 4286 1764 4338
rect 1708 4274 1764 4286
rect 1932 5124 1988 5134
rect 1932 4116 1988 5068
rect 1820 4060 1988 4116
rect 1820 3554 1876 4060
rect 2044 3556 2100 5404
rect 2156 5010 2212 5852
rect 2268 5842 2324 5852
rect 2156 4958 2158 5010
rect 2210 4958 2212 5010
rect 2156 4946 2212 4958
rect 2380 4900 2436 6524
rect 2492 6468 2548 6478
rect 2492 5122 2548 6412
rect 2492 5070 2494 5122
rect 2546 5070 2548 5122
rect 2492 5058 2548 5070
rect 2828 6466 2884 6478
rect 2828 6414 2830 6466
rect 2882 6414 2884 6466
rect 2716 5012 2772 5022
rect 2380 4844 2548 4900
rect 2380 4340 2436 4350
rect 1820 3502 1822 3554
rect 1874 3502 1876 3554
rect 1820 3490 1876 3502
rect 1932 3500 2100 3556
rect 2156 4338 2436 4340
rect 2156 4286 2382 4338
rect 2434 4286 2436 4338
rect 2156 4284 2436 4286
rect 1932 3108 1988 3500
rect 2156 3444 2212 4284
rect 2380 4274 2436 4284
rect 2044 3388 2212 3444
rect 2492 3554 2548 4844
rect 2492 3502 2494 3554
rect 2546 3502 2548 3554
rect 2044 3330 2100 3388
rect 2044 3278 2046 3330
rect 2098 3278 2100 3330
rect 2044 3266 2100 3278
rect 1932 3052 2100 3108
rect 2044 800 2100 3052
rect 2016 0 2128 800
rect 2492 756 2548 3502
rect 2716 3442 2772 4956
rect 2828 3668 2884 6414
rect 3276 6466 3332 6478
rect 3276 6414 3278 6466
rect 3330 6414 3332 6466
rect 3052 5684 3108 5694
rect 3052 5234 3108 5628
rect 3052 5182 3054 5234
rect 3106 5182 3108 5234
rect 3052 5170 3108 5182
rect 3276 3780 3332 6414
rect 3612 6468 3668 6478
rect 3612 6374 3668 6412
rect 3724 5684 3780 6636
rect 4284 6580 4340 7644
rect 4732 7364 4788 7374
rect 4844 7364 4900 8764
rect 5068 7364 5124 7374
rect 4844 7362 5124 7364
rect 4844 7310 5070 7362
rect 5122 7310 5124 7362
rect 4844 7308 5124 7310
rect 4732 7270 4788 7308
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4732 6692 4788 6702
rect 4956 6692 5012 7308
rect 5068 7298 5124 7308
rect 5180 7364 5236 8876
rect 5628 8484 5684 12908
rect 5740 12898 5796 12908
rect 5740 12404 5796 12414
rect 5852 12404 5908 14252
rect 5964 14242 6020 14252
rect 6300 13860 6356 14366
rect 6860 14418 6916 14430
rect 6860 14366 6862 14418
rect 6914 14366 6916 14418
rect 6524 13972 6580 13982
rect 6860 13972 6916 14366
rect 6524 13970 6916 13972
rect 6524 13918 6526 13970
rect 6578 13918 6916 13970
rect 6524 13916 6916 13918
rect 6524 13906 6580 13916
rect 6188 13076 6244 13086
rect 6300 13076 6356 13804
rect 6860 13748 6916 13916
rect 6972 14308 7028 14318
rect 6972 13970 7028 14252
rect 6972 13918 6974 13970
rect 7026 13918 7028 13970
rect 6972 13906 7028 13918
rect 6860 13682 6916 13692
rect 6188 13074 6356 13076
rect 6188 13022 6190 13074
rect 6242 13022 6356 13074
rect 6188 13020 6356 13022
rect 6748 13412 6804 13422
rect 6748 13074 6804 13356
rect 6748 13022 6750 13074
rect 6802 13022 6804 13074
rect 6188 12964 6244 13020
rect 6748 13010 6804 13022
rect 6188 12898 6244 12908
rect 5740 12402 5908 12404
rect 5740 12350 5742 12402
rect 5794 12350 5908 12402
rect 5740 12348 5908 12350
rect 5740 12338 5796 12348
rect 5852 10612 5908 10622
rect 5852 10610 6132 10612
rect 5852 10558 5854 10610
rect 5906 10558 6132 10610
rect 5852 10556 6132 10558
rect 5852 10546 5908 10556
rect 6076 9714 6132 10556
rect 6076 9662 6078 9714
rect 6130 9662 6132 9714
rect 6076 9650 6132 9662
rect 6412 9716 6468 9726
rect 6412 9622 6468 9660
rect 6300 9154 6356 9166
rect 6300 9102 6302 9154
rect 6354 9102 6356 9154
rect 5628 8428 6132 8484
rect 5628 7698 5684 8428
rect 5628 7646 5630 7698
rect 5682 7646 5684 7698
rect 5628 7634 5684 7646
rect 5740 8258 5796 8270
rect 5740 8206 5742 8258
rect 5794 8206 5796 8258
rect 5180 7298 5236 7308
rect 4732 6690 5012 6692
rect 4732 6638 4734 6690
rect 4786 6638 5012 6690
rect 4732 6636 5012 6638
rect 5740 6804 5796 8206
rect 6076 7698 6132 8428
rect 6300 8258 6356 9102
rect 7084 9156 7140 16044
rect 7420 14868 7476 14878
rect 7308 14812 7420 14868
rect 7308 12404 7364 14812
rect 7420 14802 7476 14812
rect 7420 14530 7476 14542
rect 7420 14478 7422 14530
rect 7474 14478 7476 14530
rect 7420 13970 7476 14478
rect 7420 13918 7422 13970
rect 7474 13918 7476 13970
rect 7420 13906 7476 13918
rect 7308 12338 7364 12348
rect 7084 9090 7140 9100
rect 6636 9044 6692 9054
rect 6636 8950 6692 8988
rect 7420 9044 7476 9054
rect 7420 8950 7476 8988
rect 6300 8206 6302 8258
rect 6354 8206 6356 8258
rect 6300 8194 6356 8206
rect 6076 7646 6078 7698
rect 6130 7646 6132 7698
rect 6076 7634 6132 7646
rect 7420 7812 7476 7822
rect 6076 7364 6132 7374
rect 6076 6804 6132 7308
rect 5740 6802 6132 6804
rect 5740 6750 6078 6802
rect 6130 6750 6132 6802
rect 5740 6748 6132 6750
rect 4732 6626 4788 6636
rect 4508 6580 4564 6590
rect 3724 5348 3780 5628
rect 3724 5282 3780 5292
rect 4172 6578 4676 6580
rect 4172 6526 4510 6578
rect 4562 6526 4676 6578
rect 4172 6524 4676 6526
rect 4172 5346 4228 6524
rect 4508 6514 4564 6524
rect 4620 6132 4676 6524
rect 4732 6132 4788 6142
rect 4620 6076 4732 6132
rect 4732 6038 4788 6076
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4172 5294 4174 5346
rect 4226 5294 4228 5346
rect 4172 5282 4228 5294
rect 4732 5348 4788 5358
rect 3500 5236 3556 5246
rect 3500 5142 3556 5180
rect 3836 5124 3892 5134
rect 3836 5030 3892 5068
rect 4732 5010 4788 5292
rect 4844 5122 4900 6636
rect 5180 6132 5236 6142
rect 5180 6038 5236 6076
rect 5740 5906 5796 6748
rect 6076 6738 6132 6748
rect 6524 7362 6580 7374
rect 6524 7310 6526 7362
rect 6578 7310 6580 7362
rect 6412 6466 6468 6478
rect 6412 6414 6414 6466
rect 6466 6414 6468 6466
rect 5740 5854 5742 5906
rect 5794 5854 5796 5906
rect 5740 5236 5796 5854
rect 6300 5908 6356 5918
rect 6412 5908 6468 6414
rect 6300 5906 6468 5908
rect 6300 5854 6302 5906
rect 6354 5854 6468 5906
rect 6300 5852 6468 5854
rect 6300 5842 6356 5852
rect 5740 5234 6020 5236
rect 5740 5182 5742 5234
rect 5794 5182 6020 5234
rect 5740 5180 6020 5182
rect 5740 5170 5796 5180
rect 4844 5070 4846 5122
rect 4898 5070 4900 5122
rect 4844 5058 4900 5070
rect 4732 4958 4734 5010
rect 4786 4958 4788 5010
rect 4732 4564 4788 4958
rect 4844 4564 4900 4574
rect 4732 4562 4900 4564
rect 4732 4510 4846 4562
rect 4898 4510 4900 4562
rect 4732 4508 4900 4510
rect 4844 4498 4900 4508
rect 5740 4564 5796 4574
rect 5740 4470 5796 4508
rect 5516 4338 5572 4350
rect 5516 4286 5518 4338
rect 5570 4286 5572 4338
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 5516 3892 5572 4286
rect 5964 4340 6020 5180
rect 6412 5124 6468 5134
rect 6524 5124 6580 7310
rect 7196 7364 7252 7374
rect 7196 7270 7252 7308
rect 6748 6580 6804 6590
rect 6748 6486 6804 6524
rect 6412 5122 6580 5124
rect 6412 5070 6414 5122
rect 6466 5070 6580 5122
rect 6412 5068 6580 5070
rect 6412 5058 6468 5068
rect 6076 4900 6132 4910
rect 6076 4898 6244 4900
rect 6076 4846 6078 4898
rect 6130 4846 6244 4898
rect 6076 4844 6244 4846
rect 6076 4834 6132 4844
rect 6076 4340 6132 4350
rect 5964 4338 6132 4340
rect 5964 4286 6078 4338
rect 6130 4286 6132 4338
rect 5964 4284 6132 4286
rect 6076 4274 6132 4284
rect 6188 4116 6244 4844
rect 5516 3826 5572 3836
rect 6076 4060 6244 4116
rect 3276 3714 3332 3724
rect 3724 3780 3780 3790
rect 3164 3668 3220 3678
rect 2828 3612 3164 3668
rect 3164 3554 3220 3612
rect 3164 3502 3166 3554
rect 3218 3502 3220 3554
rect 3164 3490 3220 3502
rect 3388 3556 3444 3566
rect 2716 3390 2718 3442
rect 2770 3390 2772 3442
rect 2716 3378 2772 3390
rect 3388 3442 3444 3500
rect 3724 3554 3780 3724
rect 5628 3780 5684 3790
rect 3724 3502 3726 3554
rect 3778 3502 3780 3554
rect 3724 3490 3780 3502
rect 4284 3668 4340 3678
rect 3388 3390 3390 3442
rect 3442 3390 3444 3442
rect 3388 3378 3444 3390
rect 4060 3444 4116 3482
rect 4060 3378 4116 3388
rect 2828 924 3220 980
rect 2828 756 2884 924
rect 3164 800 3220 924
rect 4284 800 4340 3612
rect 4396 3554 4452 3566
rect 4396 3502 4398 3554
rect 4450 3502 4452 3554
rect 4396 3332 4452 3502
rect 4956 3444 5012 3454
rect 5516 3444 5572 3454
rect 4956 3442 5572 3444
rect 4956 3390 4958 3442
rect 5010 3390 5518 3442
rect 5570 3390 5572 3442
rect 4956 3388 5572 3390
rect 4956 3378 5012 3388
rect 5516 3378 5572 3388
rect 4396 3266 4452 3276
rect 5628 1764 5684 3724
rect 5964 3556 6020 3566
rect 5964 3462 6020 3500
rect 6076 3554 6132 4060
rect 6076 3502 6078 3554
rect 6130 3502 6132 3554
rect 6076 3490 6132 3502
rect 6188 3444 6244 3482
rect 6188 3378 6244 3388
rect 5404 1708 5684 1764
rect 5404 800 5460 1708
rect 6524 800 6580 5068
rect 7084 6468 7140 6478
rect 7084 5122 7140 6412
rect 7084 5070 7086 5122
rect 7138 5070 7140 5122
rect 7084 5058 7140 5070
rect 7420 5012 7476 7756
rect 7532 7700 7588 20524
rect 8092 20580 8148 20590
rect 8204 20580 8260 20748
rect 8540 20692 8596 20702
rect 8092 20578 8260 20580
rect 8092 20526 8094 20578
rect 8146 20526 8260 20578
rect 8092 20524 8260 20526
rect 8092 20514 8148 20524
rect 7868 17444 7924 17454
rect 7868 15148 7924 17388
rect 7756 15092 7812 15102
rect 7868 15092 8036 15148
rect 7644 14532 7700 14542
rect 7756 14532 7812 15036
rect 7868 14532 7924 14542
rect 7756 14530 7924 14532
rect 7756 14478 7870 14530
rect 7922 14478 7924 14530
rect 7756 14476 7924 14478
rect 7644 14418 7700 14476
rect 7868 14466 7924 14476
rect 7644 14366 7646 14418
rect 7698 14366 7700 14418
rect 7644 14354 7700 14366
rect 7980 14308 8036 15092
rect 8204 14868 8260 20524
rect 8428 20580 8484 20590
rect 8428 20486 8484 20524
rect 8428 19348 8484 19358
rect 8428 19254 8484 19292
rect 8540 17780 8596 20636
rect 9660 20692 9716 20702
rect 9660 20598 9716 20636
rect 9884 20356 9940 21868
rect 10220 21812 10276 22428
rect 9996 21756 10276 21812
rect 9996 20916 10052 21756
rect 10332 21700 10388 23660
rect 10668 23492 10724 23502
rect 10444 23268 10500 23278
rect 10444 23266 10612 23268
rect 10444 23214 10446 23266
rect 10498 23214 10612 23266
rect 10444 23212 10612 23214
rect 10444 23202 10500 23212
rect 10556 23154 10612 23212
rect 10556 23102 10558 23154
rect 10610 23102 10612 23154
rect 10556 23090 10612 23102
rect 10668 22482 10724 23436
rect 10780 23378 10836 23886
rect 10780 23326 10782 23378
rect 10834 23326 10836 23378
rect 10780 23314 10836 23326
rect 10892 23268 10948 23278
rect 10892 23154 10948 23212
rect 10892 23102 10894 23154
rect 10946 23102 10948 23154
rect 10892 23090 10948 23102
rect 10668 22430 10670 22482
rect 10722 22430 10724 22482
rect 10668 22418 10724 22430
rect 11004 22260 11060 22270
rect 10780 22258 11060 22260
rect 10780 22206 11006 22258
rect 11058 22206 11060 22258
rect 10780 22204 11060 22206
rect 10780 22036 10836 22204
rect 11004 22194 11060 22204
rect 10332 21606 10388 21644
rect 10444 21980 10836 22036
rect 9996 20802 10052 20860
rect 9996 20750 9998 20802
rect 10050 20750 10052 20802
rect 9996 20738 10052 20750
rect 10444 20356 10500 21980
rect 10668 21810 10724 21822
rect 10668 21758 10670 21810
rect 10722 21758 10724 21810
rect 10556 20802 10612 20814
rect 10556 20750 10558 20802
rect 10610 20750 10612 20802
rect 10556 20580 10612 20750
rect 10556 20514 10612 20524
rect 9436 20300 9940 20356
rect 10108 20300 10500 20356
rect 8988 20132 9044 20142
rect 8988 20038 9044 20076
rect 8988 19348 9044 19358
rect 9436 19348 9492 20300
rect 9996 20020 10052 20030
rect 10108 20020 10164 20300
rect 9996 20018 10164 20020
rect 9996 19966 9998 20018
rect 10050 19966 10164 20018
rect 9996 19964 10164 19966
rect 9996 19954 10052 19964
rect 8988 19346 9492 19348
rect 8988 19294 8990 19346
rect 9042 19294 9492 19346
rect 8988 19292 9492 19294
rect 8988 19282 9044 19292
rect 9436 19122 9492 19292
rect 9884 19348 9940 19358
rect 9436 19070 9438 19122
rect 9490 19070 9492 19122
rect 9436 19058 9492 19070
rect 9548 19122 9604 19134
rect 9548 19070 9550 19122
rect 9602 19070 9604 19122
rect 9212 19012 9268 19022
rect 9212 18918 9268 18956
rect 9324 19010 9380 19022
rect 9324 18958 9326 19010
rect 9378 18958 9380 19010
rect 8428 17778 8596 17780
rect 8428 17726 8542 17778
rect 8594 17726 8596 17778
rect 8428 17724 8596 17726
rect 8316 16212 8372 16222
rect 8428 16212 8484 17724
rect 8540 17714 8596 17724
rect 8876 18900 8932 18910
rect 8764 17668 8820 17678
rect 8764 17574 8820 17612
rect 8876 16772 8932 18844
rect 9324 18452 9380 18958
rect 9324 18386 9380 18396
rect 9548 18116 9604 19070
rect 9100 18060 9604 18116
rect 9660 18340 9716 18350
rect 9100 17890 9156 18060
rect 9100 17838 9102 17890
rect 9154 17838 9156 17890
rect 9100 17826 9156 17838
rect 9324 17666 9380 17678
rect 9324 17614 9326 17666
rect 9378 17614 9380 17666
rect 8988 16996 9044 17006
rect 8988 16902 9044 16940
rect 9324 16884 9380 17614
rect 9660 17666 9716 18284
rect 9772 18338 9828 18350
rect 9772 18286 9774 18338
rect 9826 18286 9828 18338
rect 9772 18116 9828 18286
rect 9772 18050 9828 18060
rect 9884 17892 9940 19292
rect 9996 19234 10052 19246
rect 9996 19182 9998 19234
rect 10050 19182 10052 19234
rect 9996 19012 10052 19182
rect 9996 18946 10052 18956
rect 9660 17614 9662 17666
rect 9714 17614 9716 17666
rect 9660 17602 9716 17614
rect 9772 17836 9940 17892
rect 9996 18450 10052 18462
rect 9996 18398 9998 18450
rect 10050 18398 10052 18450
rect 9660 17108 9716 17118
rect 9772 17108 9828 17836
rect 9884 17668 9940 17678
rect 9884 17574 9940 17612
rect 9884 17444 9940 17454
rect 9996 17444 10052 18398
rect 10108 18340 10164 19964
rect 10444 20020 10500 20030
rect 10444 19926 10500 19964
rect 10556 19348 10612 19358
rect 10556 19254 10612 19292
rect 10108 18274 10164 18284
rect 10332 18450 10388 18462
rect 10332 18398 10334 18450
rect 10386 18398 10388 18450
rect 10332 17780 10388 18398
rect 10668 18450 10724 21758
rect 10780 21586 10836 21980
rect 11116 21924 11172 25228
rect 11228 25282 11284 25294
rect 11228 25230 11230 25282
rect 11282 25230 11284 25282
rect 11228 23940 11284 25230
rect 11340 24948 11396 25342
rect 11340 24882 11396 24892
rect 11564 25396 11620 25406
rect 11340 24724 11396 24734
rect 11340 24630 11396 24668
rect 11228 23874 11284 23884
rect 11564 23380 11620 25340
rect 11788 24500 11844 26852
rect 12012 25620 12068 25630
rect 12012 25526 12068 25564
rect 12124 25284 12180 31500
rect 12684 30996 12740 31500
rect 13020 31220 13076 34748
rect 13356 34130 13412 34972
rect 13356 34078 13358 34130
rect 13410 34078 13412 34130
rect 13356 34066 13412 34078
rect 13468 34690 13524 35308
rect 13468 34638 13470 34690
rect 13522 34638 13524 34690
rect 13468 34020 13524 34638
rect 13804 35140 13860 35150
rect 13804 34914 13860 35084
rect 14140 35028 14196 35644
rect 14252 35028 14308 35038
rect 14196 35026 14308 35028
rect 14196 34974 14254 35026
rect 14306 34974 14308 35026
rect 14196 34972 14308 34974
rect 14140 34934 14196 34972
rect 14252 34962 14308 34972
rect 13804 34862 13806 34914
rect 13858 34862 13860 34914
rect 13468 33964 13748 34020
rect 13468 33122 13524 33134
rect 13468 33070 13470 33122
rect 13522 33070 13524 33122
rect 13468 32900 13524 33070
rect 13468 32834 13524 32844
rect 13132 32676 13188 32686
rect 13132 32562 13188 32620
rect 13132 32510 13134 32562
rect 13186 32510 13188 32562
rect 13132 32498 13188 32510
rect 13468 32564 13524 32574
rect 13468 32470 13524 32508
rect 13356 32452 13412 32462
rect 13356 32358 13412 32396
rect 13692 32340 13748 33964
rect 13804 33234 13860 34862
rect 14364 34468 14420 36540
rect 14588 35922 14644 37100
rect 14700 37090 14756 37100
rect 14588 35870 14590 35922
rect 14642 35870 14644 35922
rect 14588 35140 14644 35870
rect 14252 34412 14420 34468
rect 14476 35084 14588 35140
rect 14476 34468 14532 35084
rect 14588 35074 14644 35084
rect 14700 36260 14756 36270
rect 14812 36260 14868 37772
rect 14924 37762 14980 37772
rect 15372 37826 15540 37828
rect 15372 37774 15486 37826
rect 15538 37774 15540 37826
rect 15372 37772 15540 37774
rect 15036 37380 15092 37390
rect 15036 37156 15092 37324
rect 15372 37268 15428 37772
rect 15484 37762 15540 37772
rect 16156 37828 16212 38670
rect 16268 37940 16324 37950
rect 16268 37846 16324 37884
rect 15484 37492 15540 37502
rect 15484 37398 15540 37436
rect 15372 37202 15428 37212
rect 15596 37268 15652 37278
rect 16044 37268 16100 37278
rect 15596 37266 16100 37268
rect 15596 37214 15598 37266
rect 15650 37214 16046 37266
rect 16098 37214 16100 37266
rect 15596 37212 16100 37214
rect 15596 37202 15652 37212
rect 16044 37202 16100 37212
rect 15036 37100 15316 37156
rect 15148 36596 15204 36606
rect 15148 36482 15204 36540
rect 15148 36430 15150 36482
rect 15202 36430 15204 36482
rect 15148 36418 15204 36430
rect 14756 36204 14868 36260
rect 15036 36258 15092 36270
rect 15036 36206 15038 36258
rect 15090 36206 15092 36258
rect 14588 34804 14644 34814
rect 14700 34804 14756 36204
rect 15036 35364 15092 36206
rect 15260 35812 15316 37100
rect 15708 37044 15764 37054
rect 16156 37044 16212 37772
rect 16380 37490 16436 42700
rect 16828 41186 16884 41198
rect 16828 41134 16830 41186
rect 16882 41134 16884 41186
rect 16828 38668 16884 41134
rect 17052 40964 17108 40974
rect 16940 39620 16996 39630
rect 16940 39526 16996 39564
rect 17052 39396 17108 40908
rect 17612 40516 17668 40526
rect 17612 40422 17668 40460
rect 17500 40404 17556 40414
rect 17500 39844 17556 40348
rect 16716 38612 16884 38668
rect 16940 39340 17108 39396
rect 17276 39788 17556 39844
rect 16716 38162 16772 38612
rect 16716 38110 16718 38162
rect 16770 38110 16772 38162
rect 16716 38098 16772 38110
rect 16604 37940 16660 37950
rect 16604 37938 16772 37940
rect 16604 37886 16606 37938
rect 16658 37886 16772 37938
rect 16604 37884 16772 37886
rect 16604 37874 16660 37884
rect 16380 37438 16382 37490
rect 16434 37438 16436 37490
rect 16380 37426 16436 37438
rect 15708 36950 15764 36988
rect 15932 36988 16212 37044
rect 16380 37266 16436 37278
rect 16380 37214 16382 37266
rect 16434 37214 16436 37266
rect 15372 36596 15428 36606
rect 15372 35922 15428 36540
rect 15372 35870 15374 35922
rect 15426 35870 15428 35922
rect 15372 35858 15428 35870
rect 15596 36482 15652 36494
rect 15596 36430 15598 36482
rect 15650 36430 15652 36482
rect 15260 35746 15316 35756
rect 15596 35588 15652 36430
rect 15820 35924 15876 35934
rect 15820 35830 15876 35868
rect 15596 35522 15652 35532
rect 15036 35308 15316 35364
rect 14588 34802 14756 34804
rect 14588 34750 14590 34802
rect 14642 34750 14756 34802
rect 14588 34748 14756 34750
rect 14588 34738 14644 34748
rect 13916 34132 13972 34142
rect 13916 34130 14084 34132
rect 13916 34078 13918 34130
rect 13970 34078 14084 34130
rect 13916 34076 14084 34078
rect 13916 34066 13972 34076
rect 13804 33182 13806 33234
rect 13858 33182 13860 33234
rect 13804 33170 13860 33182
rect 14028 33236 14084 34076
rect 14028 33170 14084 33180
rect 14252 32788 14308 34412
rect 14476 34402 14532 34412
rect 14924 34690 14980 34702
rect 14924 34638 14926 34690
rect 14978 34638 14980 34690
rect 14924 34356 14980 34638
rect 15036 34356 15092 34366
rect 14924 34300 15036 34356
rect 15092 34300 15204 34356
rect 15036 34262 15092 34300
rect 14476 34130 14532 34142
rect 14476 34078 14478 34130
rect 14530 34078 14532 34130
rect 14476 33460 14532 34078
rect 14476 33394 14532 33404
rect 14364 33122 14420 33134
rect 14364 33070 14366 33122
rect 14418 33070 14420 33122
rect 14364 32900 14420 33070
rect 14364 32834 14420 32844
rect 13804 32786 14308 32788
rect 13804 32734 14254 32786
rect 14306 32734 14308 32786
rect 13804 32732 14308 32734
rect 13804 32674 13860 32732
rect 14252 32722 14308 32732
rect 15148 32786 15204 34300
rect 15260 34244 15316 35308
rect 15372 34692 15428 34702
rect 15372 34468 15428 34636
rect 15372 34402 15428 34412
rect 15372 34244 15428 34254
rect 15260 34188 15372 34244
rect 15372 34178 15428 34188
rect 15596 33460 15652 33470
rect 15596 33366 15652 33404
rect 15820 33348 15876 33358
rect 15932 33348 15988 36988
rect 16156 36484 16212 36494
rect 16156 36482 16324 36484
rect 16156 36430 16158 36482
rect 16210 36430 16324 36482
rect 16156 36428 16324 36430
rect 16156 36418 16212 36428
rect 16156 36260 16212 36270
rect 16156 35922 16212 36204
rect 16156 35870 16158 35922
rect 16210 35870 16212 35922
rect 16156 35858 16212 35870
rect 16268 35922 16324 36428
rect 16268 35870 16270 35922
rect 16322 35870 16324 35922
rect 16268 35858 16324 35870
rect 16380 36260 16436 37214
rect 16716 37266 16772 37884
rect 16716 37214 16718 37266
rect 16770 37214 16772 37266
rect 16380 35922 16436 36204
rect 16380 35870 16382 35922
rect 16434 35870 16436 35922
rect 16380 35858 16436 35870
rect 16492 37044 16548 37054
rect 15876 33292 15988 33348
rect 16380 33572 16436 33582
rect 16492 33572 16548 36988
rect 16604 35810 16660 35822
rect 16604 35758 16606 35810
rect 16658 35758 16660 35810
rect 16604 34914 16660 35758
rect 16604 34862 16606 34914
rect 16658 34862 16660 34914
rect 16604 34850 16660 34862
rect 16716 34468 16772 37214
rect 16940 37938 16996 39340
rect 17276 38668 17332 39788
rect 17500 39618 17556 39630
rect 17500 39566 17502 39618
rect 17554 39566 17556 39618
rect 17500 39058 17556 39566
rect 17500 39006 17502 39058
rect 17554 39006 17556 39058
rect 17500 38994 17556 39006
rect 17612 38948 17668 38958
rect 17612 38854 17668 38892
rect 17388 38836 17444 38846
rect 17388 38742 17444 38780
rect 16940 37886 16942 37938
rect 16994 37886 16996 37938
rect 16940 36932 16996 37886
rect 16940 36866 16996 36876
rect 17052 38612 17332 38668
rect 17724 38668 17780 43148
rect 18396 42756 18452 42766
rect 18172 42700 18396 42756
rect 17948 39060 18004 39070
rect 17724 38612 17892 38668
rect 16940 35028 16996 35038
rect 16940 34914 16996 34972
rect 16940 34862 16942 34914
rect 16994 34862 16996 34914
rect 16940 34850 16996 34862
rect 16380 33570 16548 33572
rect 16380 33518 16382 33570
rect 16434 33518 16548 33570
rect 16380 33516 16548 33518
rect 16604 34412 16772 34468
rect 16828 34690 16884 34702
rect 16828 34638 16830 34690
rect 16882 34638 16884 34690
rect 15820 33254 15876 33292
rect 15148 32734 15150 32786
rect 15202 32734 15204 32786
rect 13804 32622 13806 32674
rect 13858 32622 13860 32674
rect 13804 32610 13860 32622
rect 12684 30930 12740 30940
rect 12796 31164 13076 31220
rect 13580 32284 13748 32340
rect 13580 31668 13636 32284
rect 15148 31948 15204 32734
rect 12572 30884 12628 30894
rect 12572 30324 12628 30828
rect 12236 30100 12292 30110
rect 12236 30006 12292 30044
rect 12572 30098 12628 30268
rect 12572 30046 12574 30098
rect 12626 30046 12628 30098
rect 12572 30034 12628 30046
rect 12348 27300 12404 27310
rect 12348 26292 12404 27244
rect 12572 27300 12628 27310
rect 12572 27076 12628 27244
rect 12572 26908 12628 27020
rect 12460 26852 12628 26908
rect 12684 26964 12740 27002
rect 12684 26898 12740 26908
rect 12460 26514 12516 26852
rect 12460 26462 12462 26514
rect 12514 26462 12516 26514
rect 12460 26450 12516 26462
rect 12348 25506 12404 26236
rect 12348 25454 12350 25506
rect 12402 25454 12404 25506
rect 12348 25442 12404 25454
rect 12684 25394 12740 25406
rect 12684 25342 12686 25394
rect 12738 25342 12740 25394
rect 12124 25228 12404 25284
rect 11900 24948 11956 24958
rect 11900 24722 11956 24892
rect 11900 24670 11902 24722
rect 11954 24670 11956 24722
rect 11900 24658 11956 24670
rect 11788 24444 12292 24500
rect 12124 24164 12180 24202
rect 12124 24098 12180 24108
rect 11676 23938 11732 23950
rect 11676 23886 11678 23938
rect 11730 23886 11732 23938
rect 11676 23604 11732 23886
rect 12124 23940 12180 23950
rect 12124 23846 12180 23884
rect 12236 23938 12292 24444
rect 12236 23886 12238 23938
rect 12290 23886 12292 23938
rect 12236 23874 12292 23886
rect 11676 23548 11844 23604
rect 11676 23380 11732 23390
rect 11228 23378 11732 23380
rect 11228 23326 11678 23378
rect 11730 23326 11732 23378
rect 11228 23324 11732 23326
rect 11228 23266 11284 23324
rect 11676 23314 11732 23324
rect 11228 23214 11230 23266
rect 11282 23214 11284 23266
rect 11228 23202 11284 23214
rect 11676 23156 11732 23166
rect 11340 23044 11396 23054
rect 10780 21534 10782 21586
rect 10834 21534 10836 21586
rect 10780 21522 10836 21534
rect 10892 21868 11172 21924
rect 11228 22988 11340 23044
rect 10780 20692 10836 20702
rect 10892 20692 10948 21868
rect 10780 20690 10948 20692
rect 10780 20638 10782 20690
rect 10834 20638 10948 20690
rect 10780 20636 10948 20638
rect 10780 20626 10836 20636
rect 10892 20244 10948 20636
rect 11116 21700 11172 21710
rect 11116 20690 11172 21644
rect 11116 20638 11118 20690
rect 11170 20638 11172 20690
rect 11116 20626 11172 20638
rect 10892 20178 10948 20188
rect 11004 19906 11060 19918
rect 11004 19854 11006 19906
rect 11058 19854 11060 19906
rect 10668 18398 10670 18450
rect 10722 18398 10724 18450
rect 10668 18386 10724 18398
rect 10892 18452 10948 18462
rect 10892 18358 10948 18396
rect 10780 18338 10836 18350
rect 10780 18286 10782 18338
rect 10834 18286 10836 18338
rect 10444 18226 10500 18238
rect 10444 18174 10446 18226
rect 10498 18174 10500 18226
rect 10444 18116 10500 18174
rect 10780 18228 10836 18286
rect 10780 18162 10836 18172
rect 10444 18050 10500 18060
rect 10332 17724 10500 17780
rect 9884 17442 10052 17444
rect 9884 17390 9886 17442
rect 9938 17390 10052 17442
rect 9884 17388 10052 17390
rect 10108 17666 10164 17678
rect 10108 17614 10110 17666
rect 10162 17614 10164 17666
rect 9884 17378 9940 17388
rect 10108 17332 10164 17614
rect 10108 17266 10164 17276
rect 10332 17554 10388 17566
rect 10332 17502 10334 17554
rect 10386 17502 10388 17554
rect 9660 17106 10052 17108
rect 9660 17054 9662 17106
rect 9714 17054 10052 17106
rect 9660 17052 10052 17054
rect 9660 17042 9716 17052
rect 9996 16996 10052 17052
rect 10332 16996 10388 17502
rect 9996 16940 10164 16996
rect 9324 16818 9380 16828
rect 9884 16884 9940 16894
rect 9940 16828 10052 16884
rect 9884 16818 9940 16828
rect 8876 16706 8932 16716
rect 9660 16772 9716 16782
rect 8316 16210 8484 16212
rect 8316 16158 8318 16210
rect 8370 16158 8484 16210
rect 8316 16156 8484 16158
rect 8316 16146 8372 16156
rect 8428 15428 8484 16156
rect 8764 16660 8820 16670
rect 8540 16100 8596 16110
rect 8540 16006 8596 16044
rect 8428 15362 8484 15372
rect 8764 15148 8820 16604
rect 8876 16212 8932 16222
rect 8876 16210 9604 16212
rect 8876 16158 8878 16210
rect 8930 16158 9604 16210
rect 8876 16156 9604 16158
rect 8876 16146 8932 16156
rect 9548 15986 9604 16156
rect 9548 15934 9550 15986
rect 9602 15934 9604 15986
rect 9548 15922 9604 15934
rect 9660 16100 9716 16716
rect 9996 16210 10052 16828
rect 9996 16158 9998 16210
rect 10050 16158 10052 16210
rect 9996 16146 10052 16158
rect 9660 15986 9716 16044
rect 9660 15934 9662 15986
rect 9714 15934 9716 15986
rect 9660 15922 9716 15934
rect 8204 14802 8260 14812
rect 8652 15092 8820 15148
rect 9212 15874 9268 15886
rect 9212 15822 9214 15874
rect 9266 15822 9268 15874
rect 7756 14252 8036 14308
rect 8428 14644 8484 14654
rect 7756 13972 7812 14252
rect 8428 14084 8484 14588
rect 8540 14532 8596 14542
rect 8540 14438 8596 14476
rect 7644 13916 7812 13972
rect 7868 14028 8484 14084
rect 7644 12964 7700 13916
rect 7756 13748 7812 13758
rect 7756 13654 7812 13692
rect 7868 13188 7924 14028
rect 7980 13860 8036 13870
rect 8036 13804 8260 13860
rect 7980 13766 8036 13804
rect 8204 13524 8260 13804
rect 8428 13858 8484 14028
rect 8428 13806 8430 13858
rect 8482 13806 8484 13858
rect 8428 13794 8484 13806
rect 8204 13468 8484 13524
rect 7980 13188 8036 13198
rect 7868 13186 8036 13188
rect 7868 13134 7982 13186
rect 8034 13134 8036 13186
rect 7868 13132 8036 13134
rect 7980 13122 8036 13132
rect 7644 12908 8148 12964
rect 7644 12740 7700 12750
rect 7644 12738 7924 12740
rect 7644 12686 7646 12738
rect 7698 12686 7924 12738
rect 7644 12684 7924 12686
rect 7644 12674 7700 12684
rect 7868 12290 7924 12684
rect 7868 12238 7870 12290
rect 7922 12238 7924 12290
rect 7868 12226 7924 12238
rect 7980 11732 8036 11742
rect 7868 11394 7924 11406
rect 7868 11342 7870 11394
rect 7922 11342 7924 11394
rect 7868 11172 7924 11342
rect 7868 11106 7924 11116
rect 7980 10050 8036 11676
rect 8092 10836 8148 12908
rect 8428 12962 8484 13468
rect 8428 12910 8430 12962
rect 8482 12910 8484 12962
rect 8428 12898 8484 12910
rect 8204 12290 8260 12302
rect 8204 12238 8206 12290
rect 8258 12238 8260 12290
rect 8204 11396 8260 12238
rect 8540 11396 8596 11406
rect 8204 11394 8596 11396
rect 8204 11342 8542 11394
rect 8594 11342 8596 11394
rect 8204 11340 8596 11342
rect 8540 11330 8596 11340
rect 8204 10836 8260 10846
rect 8652 10836 8708 15092
rect 9212 13524 9268 15822
rect 9436 15876 9492 15886
rect 9436 15782 9492 15820
rect 9660 15428 9716 15438
rect 9660 15334 9716 15372
rect 9884 15090 9940 15102
rect 9884 15038 9886 15090
rect 9938 15038 9940 15090
rect 9884 13748 9940 15038
rect 10108 15092 10164 16940
rect 10332 16930 10388 16940
rect 10444 16884 10500 17724
rect 10892 17220 10948 17230
rect 10892 17106 10948 17164
rect 10892 17054 10894 17106
rect 10946 17054 10948 17106
rect 10892 17042 10948 17054
rect 10444 16818 10500 16828
rect 10220 16770 10276 16782
rect 10220 16718 10222 16770
rect 10274 16718 10276 16770
rect 10220 16658 10276 16718
rect 10220 16606 10222 16658
rect 10274 16606 10276 16658
rect 10220 16594 10276 16606
rect 10780 16100 10836 16110
rect 10220 16044 10724 16100
rect 10220 15538 10276 16044
rect 10668 15986 10724 16044
rect 10668 15934 10670 15986
rect 10722 15934 10724 15986
rect 10668 15922 10724 15934
rect 10780 15986 10836 16044
rect 10780 15934 10782 15986
rect 10834 15934 10836 15986
rect 10780 15922 10836 15934
rect 10220 15486 10222 15538
rect 10274 15486 10276 15538
rect 10220 15474 10276 15486
rect 10332 15874 10388 15886
rect 10332 15822 10334 15874
rect 10386 15822 10388 15874
rect 10108 15026 10164 15036
rect 10332 14756 10388 15822
rect 10556 15876 10612 15886
rect 10556 15782 10612 15820
rect 11004 15148 11060 19854
rect 11228 18116 11284 22988
rect 11340 22978 11396 22988
rect 11564 22484 11620 22494
rect 11564 22370 11620 22428
rect 11676 22482 11732 23100
rect 11788 23044 11844 23548
rect 12124 23156 12180 23194
rect 12180 23100 12292 23156
rect 12124 23090 12180 23100
rect 11788 22978 11844 22988
rect 11676 22430 11678 22482
rect 11730 22430 11732 22482
rect 11676 22418 11732 22430
rect 12124 22930 12180 22942
rect 12124 22878 12126 22930
rect 12178 22878 12180 22930
rect 11564 22318 11566 22370
rect 11618 22318 11620 22370
rect 11564 22306 11620 22318
rect 12124 22260 12180 22878
rect 11900 22258 12180 22260
rect 11900 22206 12126 22258
rect 12178 22206 12180 22258
rect 11900 22204 12180 22206
rect 11340 21586 11396 21598
rect 11340 21534 11342 21586
rect 11394 21534 11396 21586
rect 11340 20132 11396 21534
rect 11564 20802 11620 20814
rect 11564 20750 11566 20802
rect 11618 20750 11620 20802
rect 11340 20066 11396 20076
rect 11452 20578 11508 20590
rect 11452 20526 11454 20578
rect 11506 20526 11508 20578
rect 11228 18050 11284 18060
rect 11340 18452 11396 18462
rect 11116 17892 11172 17902
rect 11116 17778 11172 17836
rect 11116 17726 11118 17778
rect 11170 17726 11172 17778
rect 11116 17714 11172 17726
rect 11228 17666 11284 17678
rect 11228 17614 11230 17666
rect 11282 17614 11284 17666
rect 11116 17556 11172 17566
rect 11116 16210 11172 17500
rect 11116 16158 11118 16210
rect 11170 16158 11172 16210
rect 11116 16146 11172 16158
rect 11004 15092 11172 15148
rect 10332 14690 10388 14700
rect 11004 14644 11060 14654
rect 11004 14550 11060 14588
rect 11116 14308 11172 15092
rect 11116 14242 11172 14252
rect 9884 13682 9940 13692
rect 9212 13458 9268 13468
rect 8764 12852 8820 12862
rect 8764 11732 8820 12796
rect 11228 12852 11284 17614
rect 11340 17668 11396 18396
rect 11452 18450 11508 20526
rect 11564 20020 11620 20750
rect 11564 19954 11620 19964
rect 11788 18452 11844 18462
rect 11452 18398 11454 18450
rect 11506 18398 11508 18450
rect 11452 18386 11508 18398
rect 11676 18450 11844 18452
rect 11676 18398 11790 18450
rect 11842 18398 11844 18450
rect 11676 18396 11844 18398
rect 11340 17106 11396 17612
rect 11564 18340 11620 18350
rect 11564 17666 11620 18284
rect 11564 17614 11566 17666
rect 11618 17614 11620 17666
rect 11564 17602 11620 17614
rect 11676 17668 11732 18396
rect 11788 18386 11844 18396
rect 11788 17892 11844 17902
rect 11788 17798 11844 17836
rect 11676 17602 11732 17612
rect 11900 17444 11956 22204
rect 12124 22194 12180 22204
rect 12236 21586 12292 23100
rect 12236 21534 12238 21586
rect 12290 21534 12292 21586
rect 12236 21522 12292 21534
rect 12124 20804 12180 20814
rect 12124 20710 12180 20748
rect 12348 18788 12404 25228
rect 12460 25282 12516 25294
rect 12460 25230 12462 25282
rect 12514 25230 12516 25282
rect 12460 24948 12516 25230
rect 12460 24882 12516 24892
rect 12460 24612 12516 24622
rect 12460 22372 12516 24556
rect 12684 24388 12740 25342
rect 12684 24322 12740 24332
rect 12684 23940 12740 23950
rect 12572 23044 12628 23054
rect 12572 22950 12628 22988
rect 12684 22930 12740 23884
rect 12684 22878 12686 22930
rect 12738 22878 12740 22930
rect 12684 22866 12740 22878
rect 12796 22820 12852 31164
rect 13468 30436 13524 30446
rect 13356 29204 13412 29214
rect 13356 29110 13412 29148
rect 12908 25508 12964 25518
rect 12908 25414 12964 25452
rect 13468 25506 13524 30380
rect 13580 28642 13636 31612
rect 14924 31892 15204 31948
rect 15260 33236 15316 33246
rect 14588 31106 14644 31118
rect 14588 31054 14590 31106
rect 14642 31054 14644 31106
rect 14588 30884 14644 31054
rect 14588 30818 14644 30828
rect 14812 30994 14868 31006
rect 14812 30942 14814 30994
rect 14866 30942 14868 30994
rect 13692 30772 13748 30782
rect 13692 30770 13860 30772
rect 13692 30718 13694 30770
rect 13746 30718 13860 30770
rect 13692 30716 13860 30718
rect 13692 30706 13748 30716
rect 13692 29204 13748 29214
rect 13692 29110 13748 29148
rect 13580 28590 13582 28642
rect 13634 28590 13636 28642
rect 13580 28578 13636 28590
rect 13804 28642 13860 30716
rect 14028 30770 14084 30782
rect 14028 30718 14030 30770
rect 14082 30718 14084 30770
rect 14028 30436 14084 30718
rect 14812 30660 14868 30942
rect 14812 30594 14868 30604
rect 14028 30370 14084 30380
rect 13916 30100 13972 30110
rect 13916 29540 13972 30044
rect 13916 29446 13972 29484
rect 14476 29538 14532 29550
rect 14476 29486 14478 29538
rect 14530 29486 14532 29538
rect 14476 28980 14532 29486
rect 13804 28590 13806 28642
rect 13858 28590 13860 28642
rect 13804 28578 13860 28590
rect 13916 28924 14532 28980
rect 13804 28084 13860 28094
rect 13916 28084 13972 28924
rect 14252 28754 14308 28766
rect 14252 28702 14254 28754
rect 14306 28702 14308 28754
rect 13804 28082 13972 28084
rect 13804 28030 13806 28082
rect 13858 28030 13972 28082
rect 13804 28028 13972 28030
rect 13804 28018 13860 28028
rect 13580 27972 13636 27982
rect 13580 27188 13636 27916
rect 13580 27122 13636 27132
rect 13692 27074 13748 27086
rect 13692 27022 13694 27074
rect 13746 27022 13748 27074
rect 13468 25454 13470 25506
rect 13522 25454 13524 25506
rect 13468 24948 13524 25454
rect 13580 25618 13636 25630
rect 13580 25566 13582 25618
rect 13634 25566 13636 25618
rect 13580 25508 13636 25566
rect 13692 25620 13748 27022
rect 13804 26292 13860 26302
rect 13804 26198 13860 26236
rect 13916 25732 13972 28028
rect 14028 28642 14084 28654
rect 14028 28590 14030 28642
rect 14082 28590 14084 28642
rect 14028 25956 14084 28590
rect 14252 28644 14308 28702
rect 14364 28644 14420 28654
rect 14252 28588 14364 28644
rect 14364 28578 14420 28588
rect 14476 28530 14532 28924
rect 14924 28868 14980 31892
rect 15260 31780 15316 33180
rect 15260 31686 15316 31724
rect 15484 33234 15540 33246
rect 15484 33182 15486 33234
rect 15538 33182 15540 33234
rect 15484 32674 15540 33182
rect 16044 33236 16100 33246
rect 16044 33142 16100 33180
rect 15484 32622 15486 32674
rect 15538 32622 15540 32674
rect 15372 31444 15428 31454
rect 15372 30882 15428 31388
rect 15484 31108 15540 32622
rect 15932 32452 15988 32462
rect 15820 31778 15876 31790
rect 15820 31726 15822 31778
rect 15874 31726 15876 31778
rect 15820 31220 15876 31726
rect 15820 31154 15876 31164
rect 15484 31042 15540 31052
rect 15372 30830 15374 30882
rect 15426 30830 15428 30882
rect 15372 30660 15428 30830
rect 15372 30594 15428 30604
rect 15708 29652 15764 29662
rect 15708 29428 15764 29596
rect 15148 29426 15764 29428
rect 15148 29374 15710 29426
rect 15762 29374 15764 29426
rect 15148 29372 15764 29374
rect 15148 28980 15204 29372
rect 15708 29362 15764 29372
rect 14476 28478 14478 28530
rect 14530 28478 14532 28530
rect 14476 28466 14532 28478
rect 14812 28812 14980 28868
rect 15036 28924 15204 28980
rect 15260 29204 15316 29214
rect 14588 28418 14644 28430
rect 14588 28366 14590 28418
rect 14642 28366 14644 28418
rect 14140 27972 14196 27982
rect 14140 27878 14196 27916
rect 14476 27972 14532 27982
rect 14476 27878 14532 27916
rect 14588 27524 14644 28366
rect 14812 28308 14868 28812
rect 14812 28242 14868 28252
rect 14924 28644 14980 28654
rect 14588 27458 14644 27468
rect 14812 27970 14868 27982
rect 14812 27918 14814 27970
rect 14866 27918 14868 27970
rect 14476 27188 14532 27198
rect 14532 27132 14644 27188
rect 14476 27122 14532 27132
rect 14140 27086 14196 27098
rect 14140 27034 14142 27086
rect 14194 27076 14196 27086
rect 14194 27034 14420 27076
rect 14140 27020 14420 27034
rect 14364 26628 14420 27020
rect 14140 26572 14420 26628
rect 14140 26514 14196 26572
rect 14140 26462 14142 26514
rect 14194 26462 14196 26514
rect 14140 26450 14196 26462
rect 14252 26292 14308 26302
rect 14476 26292 14532 26302
rect 14252 26290 14420 26292
rect 14252 26238 14254 26290
rect 14306 26238 14420 26290
rect 14252 26236 14420 26238
rect 14252 26226 14308 26236
rect 14028 25890 14084 25900
rect 13916 25676 14084 25732
rect 13692 25564 13972 25620
rect 13580 25442 13636 25452
rect 13804 25394 13860 25406
rect 13804 25342 13806 25394
rect 13858 25342 13860 25394
rect 13804 25284 13860 25342
rect 13804 25218 13860 25228
rect 13468 24882 13524 24892
rect 13468 24612 13524 24622
rect 13356 24388 13412 24398
rect 12908 23716 12964 23726
rect 12908 23378 12964 23660
rect 12908 23326 12910 23378
rect 12962 23326 12964 23378
rect 12908 23314 12964 23326
rect 13020 23154 13076 23166
rect 13020 23102 13022 23154
rect 13074 23102 13076 23154
rect 12796 22764 12964 22820
rect 12460 22278 12516 22316
rect 12796 22596 12852 22606
rect 12684 21474 12740 21486
rect 12684 21422 12686 21474
rect 12738 21422 12740 21474
rect 12684 20804 12740 21422
rect 12684 20738 12740 20748
rect 12796 20356 12852 22540
rect 12908 22484 12964 22764
rect 12908 22390 12964 22428
rect 13020 21812 13076 23102
rect 13132 23156 13188 23166
rect 13356 23156 13412 24332
rect 13132 23154 13412 23156
rect 13132 23102 13134 23154
rect 13186 23102 13412 23154
rect 13132 23100 13412 23102
rect 13132 23090 13188 23100
rect 13020 21746 13076 21756
rect 13132 22820 13188 22830
rect 13132 21586 13188 22764
rect 13132 21534 13134 21586
rect 13186 21534 13188 21586
rect 13132 21522 13188 21534
rect 13356 21028 13412 23100
rect 13468 23156 13524 24556
rect 13580 24052 13636 24062
rect 13580 23958 13636 23996
rect 13804 23716 13860 23726
rect 13692 23714 13860 23716
rect 13692 23662 13806 23714
rect 13858 23662 13860 23714
rect 13692 23660 13860 23662
rect 13468 22484 13524 23100
rect 13580 23156 13636 23166
rect 13692 23156 13748 23660
rect 13804 23650 13860 23660
rect 13580 23154 13748 23156
rect 13580 23102 13582 23154
rect 13634 23102 13748 23154
rect 13580 23100 13748 23102
rect 13916 23154 13972 25564
rect 14028 23826 14084 25676
rect 14252 24948 14308 24958
rect 14252 24854 14308 24892
rect 14364 24500 14420 26236
rect 14476 26198 14532 26236
rect 14364 24434 14420 24444
rect 14476 25956 14532 25966
rect 14476 24276 14532 25900
rect 14252 24220 14532 24276
rect 14140 24052 14196 24062
rect 14140 23938 14196 23996
rect 14140 23886 14142 23938
rect 14194 23886 14196 23938
rect 14140 23874 14196 23886
rect 14028 23774 14030 23826
rect 14082 23774 14084 23826
rect 14028 23762 14084 23774
rect 13916 23102 13918 23154
rect 13970 23102 13972 23154
rect 13580 23090 13636 23100
rect 13916 22820 13972 23102
rect 13916 22754 13972 22764
rect 13580 22484 13636 22494
rect 13468 22482 13636 22484
rect 13468 22430 13582 22482
rect 13634 22430 13636 22482
rect 13468 22428 13636 22430
rect 13580 22418 13636 22428
rect 14028 22260 14084 22270
rect 14028 22146 14084 22204
rect 14028 22094 14030 22146
rect 14082 22094 14084 22146
rect 13580 21812 13636 21822
rect 13580 21586 13636 21756
rect 14028 21700 14084 22094
rect 13580 21534 13582 21586
rect 13634 21534 13636 21586
rect 13580 21522 13636 21534
rect 13916 21644 14028 21700
rect 13580 21140 13636 21150
rect 13580 21028 13636 21084
rect 13356 21026 13636 21028
rect 13356 20974 13582 21026
rect 13634 20974 13636 21026
rect 13356 20972 13636 20974
rect 13580 20962 13636 20972
rect 13804 20804 13860 20814
rect 12124 18732 12404 18788
rect 12684 20300 12852 20356
rect 13692 20748 13804 20804
rect 12124 18452 12180 18732
rect 12124 18386 12180 18396
rect 12348 18452 12404 18462
rect 12348 18358 12404 18396
rect 12460 18450 12516 18462
rect 12460 18398 12462 18450
rect 12514 18398 12516 18450
rect 12236 18338 12292 18350
rect 12236 18286 12238 18338
rect 12290 18286 12292 18338
rect 12012 18226 12068 18238
rect 12012 18174 12014 18226
rect 12066 18174 12068 18226
rect 12012 18116 12068 18174
rect 12012 18050 12068 18060
rect 12124 17780 12180 17790
rect 12236 17780 12292 18286
rect 12124 17778 12292 17780
rect 12124 17726 12126 17778
rect 12178 17726 12292 17778
rect 12124 17724 12292 17726
rect 12460 17780 12516 18398
rect 12124 17714 12180 17724
rect 12460 17714 12516 17724
rect 11340 17054 11342 17106
rect 11394 17054 11396 17106
rect 11340 17042 11396 17054
rect 11564 17388 11956 17444
rect 12012 17666 12068 17678
rect 12012 17614 12014 17666
rect 12066 17614 12068 17666
rect 11564 16658 11620 17388
rect 12012 17220 12068 17614
rect 12012 17154 12068 17164
rect 12236 17554 12292 17566
rect 12236 17502 12238 17554
rect 12290 17502 12292 17554
rect 11900 16996 11956 17006
rect 11900 16902 11956 16940
rect 11564 16606 11566 16658
rect 11618 16606 11620 16658
rect 11564 16210 11620 16606
rect 12124 16660 12180 16670
rect 12124 16566 12180 16604
rect 11564 16158 11566 16210
rect 11618 16158 11620 16210
rect 11564 15876 11620 16158
rect 11564 15810 11620 15820
rect 11676 15316 11732 15326
rect 11676 15222 11732 15260
rect 11564 15092 11620 15102
rect 11564 14642 11620 15036
rect 11564 14590 11566 14642
rect 11618 14590 11620 14642
rect 11564 14578 11620 14590
rect 12236 14644 12292 17502
rect 12460 17556 12516 17566
rect 12460 17106 12516 17500
rect 12460 17054 12462 17106
rect 12514 17054 12516 17106
rect 12460 17042 12516 17054
rect 12684 16996 12740 20300
rect 12796 20132 12852 20142
rect 12796 19236 12852 20076
rect 13356 20132 13412 20142
rect 13356 20018 13412 20076
rect 13356 19966 13358 20018
rect 13410 19966 13412 20018
rect 13356 19954 13412 19966
rect 12796 19234 12964 19236
rect 12796 19182 12798 19234
rect 12850 19182 12964 19234
rect 12796 19180 12964 19182
rect 12796 19170 12852 19180
rect 12908 17778 12964 19180
rect 13692 19234 13748 20748
rect 13804 20710 13860 20748
rect 13916 20130 13972 21644
rect 14028 21634 14084 21644
rect 14252 21026 14308 24220
rect 14476 23940 14532 23950
rect 14588 23940 14644 27132
rect 14812 26908 14868 27918
rect 14924 27188 14980 28588
rect 15036 27858 15092 28924
rect 15036 27806 15038 27858
rect 15090 27806 15092 27858
rect 15036 27794 15092 27806
rect 14924 27122 14980 27132
rect 15036 27524 15092 27534
rect 15036 27076 15092 27468
rect 15036 27010 15092 27020
rect 14812 26852 14980 26908
rect 14924 26516 14980 26852
rect 14812 26460 14980 26516
rect 14812 26066 14868 26460
rect 14924 26292 14980 26302
rect 14924 26198 14980 26236
rect 15148 26292 15204 26302
rect 15260 26292 15316 29148
rect 15148 26290 15316 26292
rect 15148 26238 15150 26290
rect 15202 26238 15316 26290
rect 15148 26236 15316 26238
rect 15372 26964 15428 26974
rect 15148 26226 15204 26236
rect 14812 26014 14814 26066
rect 14866 26014 14868 26066
rect 14812 25284 14868 26014
rect 14812 25218 14868 25228
rect 14924 25956 14980 25966
rect 14924 24836 14980 25900
rect 15372 25844 15428 26908
rect 15932 26908 15988 32396
rect 16380 31892 16436 33516
rect 16492 33236 16548 33246
rect 16492 33142 16548 33180
rect 16044 31836 16380 31892
rect 16044 30098 16100 31836
rect 16380 31826 16436 31836
rect 16604 31108 16660 34412
rect 16828 34132 16884 34638
rect 16716 34076 16828 34132
rect 16716 33346 16772 34076
rect 16828 34038 16884 34076
rect 16716 33294 16718 33346
rect 16770 33294 16772 33346
rect 16716 33282 16772 33294
rect 16604 31042 16660 31052
rect 16044 30046 16046 30098
rect 16098 30046 16100 30098
rect 16044 30034 16100 30046
rect 16380 29986 16436 29998
rect 16380 29934 16382 29986
rect 16434 29934 16436 29986
rect 16380 29652 16436 29934
rect 16380 29586 16436 29596
rect 17052 29428 17108 38612
rect 17724 38276 17780 38286
rect 17612 38164 17668 38174
rect 17164 38162 17668 38164
rect 17164 38110 17614 38162
rect 17666 38110 17668 38162
rect 17164 38108 17668 38110
rect 17164 38050 17220 38108
rect 17612 38098 17668 38108
rect 17164 37998 17166 38050
rect 17218 37998 17220 38050
rect 17164 37986 17220 37998
rect 17500 37938 17556 37950
rect 17500 37886 17502 37938
rect 17554 37886 17556 37938
rect 17500 37044 17556 37886
rect 17724 37940 17780 38220
rect 17724 37846 17780 37884
rect 17500 36978 17556 36988
rect 17612 37828 17668 37838
rect 17388 34356 17444 34366
rect 17388 34262 17444 34300
rect 17276 34020 17332 34030
rect 17164 33570 17220 33582
rect 17164 33518 17166 33570
rect 17218 33518 17220 33570
rect 17164 33458 17220 33518
rect 17164 33406 17166 33458
rect 17218 33406 17220 33458
rect 17164 33394 17220 33406
rect 17276 33236 17332 33964
rect 16156 29314 16212 29326
rect 16156 29262 16158 29314
rect 16210 29262 16212 29314
rect 16156 28532 16212 29262
rect 16156 28084 16212 28476
rect 16604 29204 16660 29214
rect 16604 28866 16660 29148
rect 16604 28814 16606 28866
rect 16658 28814 16660 28866
rect 16492 28084 16548 28094
rect 16156 28082 16548 28084
rect 16156 28030 16494 28082
rect 16546 28030 16548 28082
rect 16156 28028 16548 28030
rect 16492 28018 16548 28028
rect 16604 27186 16660 28814
rect 17052 28756 17108 29372
rect 17052 28690 17108 28700
rect 17164 33180 17332 33236
rect 16940 28644 16996 28682
rect 16940 28578 16996 28588
rect 17164 28532 17220 33180
rect 17388 32452 17444 32462
rect 17276 32450 17444 32452
rect 17276 32398 17390 32450
rect 17442 32398 17444 32450
rect 17276 32396 17444 32398
rect 17276 29540 17332 32396
rect 17388 32386 17444 32396
rect 17500 31220 17556 31230
rect 17500 31126 17556 31164
rect 17388 31108 17444 31118
rect 17388 31014 17444 31052
rect 17276 29474 17332 29484
rect 17388 28756 17444 28766
rect 17388 28662 17444 28700
rect 17052 28476 17220 28532
rect 16716 28418 16772 28430
rect 16716 28366 16718 28418
rect 16770 28366 16772 28418
rect 16716 27636 16772 28366
rect 16940 28420 16996 28430
rect 16828 27970 16884 27982
rect 16828 27918 16830 27970
rect 16882 27918 16884 27970
rect 16828 27860 16884 27918
rect 16828 27794 16884 27804
rect 16716 27570 16772 27580
rect 16604 27134 16606 27186
rect 16658 27134 16660 27186
rect 16604 27122 16660 27134
rect 16940 26962 16996 28364
rect 16940 26910 16942 26962
rect 16994 26910 16996 26962
rect 16940 26908 16996 26910
rect 15932 26852 16100 26908
rect 15372 25778 15428 25788
rect 14812 24780 14980 24836
rect 14700 24724 14756 24762
rect 14700 24658 14756 24668
rect 14476 23938 14644 23940
rect 14476 23886 14478 23938
rect 14530 23886 14644 23938
rect 14476 23884 14644 23886
rect 14700 24500 14756 24510
rect 14700 23938 14756 24444
rect 14700 23886 14702 23938
rect 14754 23886 14756 23938
rect 14476 23716 14532 23884
rect 14476 23650 14532 23660
rect 14588 23714 14644 23726
rect 14588 23662 14590 23714
rect 14642 23662 14644 23714
rect 14476 23156 14532 23166
rect 14588 23156 14644 23662
rect 14700 23716 14756 23886
rect 14700 23650 14756 23660
rect 14476 23154 14644 23156
rect 14476 23102 14478 23154
rect 14530 23102 14644 23154
rect 14476 23100 14644 23102
rect 14476 23090 14532 23100
rect 14252 20974 14254 21026
rect 14306 20974 14308 21026
rect 14252 20962 14308 20974
rect 14364 21812 14420 21822
rect 14364 21026 14420 21756
rect 14812 21364 14868 24780
rect 15148 24612 15204 24622
rect 15036 24610 15204 24612
rect 15036 24558 15150 24610
rect 15202 24558 15204 24610
rect 15036 24556 15204 24558
rect 15036 24052 15092 24556
rect 15148 24546 15204 24556
rect 15484 24164 15540 24174
rect 15036 23716 15092 23996
rect 15148 24162 15540 24164
rect 15148 24110 15486 24162
rect 15538 24110 15540 24162
rect 15148 24108 15540 24110
rect 15148 23938 15204 24108
rect 15484 24098 15540 24108
rect 15148 23886 15150 23938
rect 15202 23886 15204 23938
rect 15148 23874 15204 23886
rect 16044 23938 16100 26852
rect 16604 26852 16996 26908
rect 16604 26178 16660 26852
rect 16604 26126 16606 26178
rect 16658 26126 16660 26178
rect 16044 23886 16046 23938
rect 16098 23886 16100 23938
rect 16044 23874 16100 23886
rect 16156 25284 16212 25294
rect 15372 23828 15428 23838
rect 15260 23826 15428 23828
rect 15260 23774 15374 23826
rect 15426 23774 15428 23826
rect 15260 23772 15428 23774
rect 15260 23716 15316 23772
rect 15372 23762 15428 23772
rect 15484 23828 15540 23838
rect 15484 23734 15540 23772
rect 15036 23660 15316 23716
rect 14588 21308 14812 21364
rect 14364 20974 14366 21026
rect 14418 20974 14420 21026
rect 14364 20962 14420 20974
rect 14476 21252 14532 21262
rect 14140 20692 14196 20702
rect 14140 20598 14196 20636
rect 13916 20078 13918 20130
rect 13970 20078 13972 20130
rect 13916 20066 13972 20078
rect 14364 20244 14420 20254
rect 14476 20244 14532 21196
rect 14420 20188 14532 20244
rect 14364 20130 14420 20188
rect 14364 20078 14366 20130
rect 14418 20078 14420 20130
rect 14364 20066 14420 20078
rect 13692 19182 13694 19234
rect 13746 19182 13748 19234
rect 13468 19012 13524 19022
rect 13468 18918 13524 18956
rect 13692 18788 13748 19182
rect 14364 19234 14420 19246
rect 14364 19182 14366 19234
rect 14418 19182 14420 19234
rect 14364 19124 14420 19182
rect 13356 18732 13748 18788
rect 13916 19012 13972 19022
rect 13132 18340 13188 18350
rect 13356 18340 13412 18732
rect 13132 18338 13412 18340
rect 13132 18286 13134 18338
rect 13186 18286 13412 18338
rect 13132 18284 13412 18286
rect 13804 18340 13860 18350
rect 12908 17726 12910 17778
rect 12962 17726 12964 17778
rect 12908 17714 12964 17726
rect 13020 18116 13076 18126
rect 13020 17106 13076 18060
rect 13020 17054 13022 17106
rect 13074 17054 13076 17106
rect 13020 17042 13076 17054
rect 12684 16212 12740 16940
rect 12796 16212 12852 16222
rect 12684 16210 12852 16212
rect 12684 16158 12798 16210
rect 12850 16158 12852 16210
rect 12684 16156 12852 16158
rect 12796 16146 12852 16156
rect 12796 15428 12852 15438
rect 12348 15202 12404 15214
rect 12348 15150 12350 15202
rect 12402 15150 12404 15202
rect 12348 15148 12404 15150
rect 12348 15092 12628 15148
rect 12572 14754 12628 15092
rect 12572 14702 12574 14754
rect 12626 14702 12628 14754
rect 12572 14690 12628 14702
rect 12236 14578 12292 14588
rect 8764 11666 8820 11676
rect 8876 12740 8932 12750
rect 8092 10834 8260 10836
rect 8092 10782 8206 10834
rect 8258 10782 8260 10834
rect 8092 10780 8260 10782
rect 7980 9998 7982 10050
rect 8034 9998 8036 10050
rect 7980 9986 8036 9998
rect 7644 9716 7700 9726
rect 8204 9716 8260 10780
rect 8428 10780 8708 10836
rect 7644 9622 7700 9660
rect 7756 9660 8204 9716
rect 7756 9042 7812 9660
rect 8204 9650 8260 9660
rect 8316 9714 8372 9726
rect 8316 9662 8318 9714
rect 8370 9662 8372 9714
rect 8316 9044 8372 9662
rect 7756 8990 7758 9042
rect 7810 8990 7812 9042
rect 7756 8978 7812 8990
rect 7868 8988 8316 9044
rect 7532 7634 7588 7644
rect 7756 7700 7812 7710
rect 7868 7700 7924 8988
rect 8316 8950 8372 8988
rect 8428 9154 8484 10780
rect 8652 10612 8708 10622
rect 8652 10518 8708 10556
rect 8540 9716 8596 9726
rect 8540 9622 8596 9660
rect 8428 9102 8430 9154
rect 8482 9102 8484 9154
rect 8428 8372 8484 9102
rect 8652 8372 8708 8382
rect 8428 8370 8708 8372
rect 8428 8318 8654 8370
rect 8706 8318 8708 8370
rect 8428 8316 8708 8318
rect 8204 7700 8260 7710
rect 7756 7698 8148 7700
rect 7756 7646 7758 7698
rect 7810 7646 8148 7698
rect 7756 7644 8148 7646
rect 7756 7634 7812 7644
rect 7868 7250 7924 7262
rect 7868 7198 7870 7250
rect 7922 7198 7924 7250
rect 7868 6914 7924 7198
rect 7868 6862 7870 6914
rect 7922 6862 7924 6914
rect 7868 6850 7924 6862
rect 7532 6580 7588 6590
rect 7532 6486 7588 6524
rect 8092 6578 8148 7644
rect 8204 6804 8260 7644
rect 8428 7250 8484 8316
rect 8652 8306 8708 8316
rect 8540 7364 8596 7374
rect 8540 7270 8596 7308
rect 8428 7198 8430 7250
rect 8482 7198 8484 7250
rect 8428 7186 8484 7198
rect 8876 7028 8932 12684
rect 11228 12292 11284 12796
rect 11004 12236 11284 12292
rect 11340 14308 11396 14318
rect 11340 13746 11396 14252
rect 12684 14306 12740 14318
rect 12684 14254 12686 14306
rect 12738 14254 12740 14306
rect 12012 13972 12068 13982
rect 12012 13858 12068 13916
rect 12012 13806 12014 13858
rect 12066 13806 12068 13858
rect 12012 13794 12068 13806
rect 11340 13694 11342 13746
rect 11394 13694 11396 13746
rect 11004 11506 11060 12236
rect 11004 11454 11006 11506
rect 11058 11454 11060 11506
rect 11004 11442 11060 11454
rect 11340 11508 11396 13694
rect 12124 12740 12180 12750
rect 12348 12740 12404 12750
rect 12180 12738 12404 12740
rect 12180 12686 12350 12738
rect 12402 12686 12404 12738
rect 12180 12684 12404 12686
rect 12124 12646 12180 12684
rect 12348 12180 12404 12684
rect 12348 12114 12404 12124
rect 11452 11508 11508 11518
rect 11340 11506 11508 11508
rect 11340 11454 11454 11506
rect 11506 11454 11508 11506
rect 11340 11452 11508 11454
rect 9324 10948 9380 10958
rect 8988 8258 9044 8270
rect 8988 8206 8990 8258
rect 9042 8206 9044 8258
rect 8988 7364 9044 8206
rect 9324 7700 9380 10892
rect 9660 10612 9716 10622
rect 9660 10518 9716 10556
rect 11452 10612 11508 11452
rect 10332 10500 10388 10510
rect 10332 10498 10612 10500
rect 10332 10446 10334 10498
rect 10386 10446 10612 10498
rect 10332 10444 10612 10446
rect 10332 10434 10388 10444
rect 10556 9714 10612 10444
rect 10892 10388 10948 10398
rect 10892 9826 10948 10332
rect 11452 9940 11508 10556
rect 12348 11282 12404 11294
rect 12348 11230 12350 11282
rect 12402 11230 12404 11282
rect 12348 10050 12404 11230
rect 12348 9998 12350 10050
rect 12402 9998 12404 10050
rect 12348 9986 12404 9998
rect 12460 10500 12516 10510
rect 10892 9774 10894 9826
rect 10946 9774 10948 9826
rect 10892 9762 10948 9774
rect 11340 9884 11452 9940
rect 10556 9662 10558 9714
rect 10610 9662 10612 9714
rect 10556 9650 10612 9662
rect 9436 9602 9492 9614
rect 9436 9550 9438 9602
rect 9490 9550 9492 9602
rect 9436 9044 9492 9550
rect 11004 9604 11060 9614
rect 11004 9266 11060 9548
rect 11004 9214 11006 9266
rect 11058 9214 11060 9266
rect 11004 9202 11060 9214
rect 11340 9266 11396 9884
rect 11452 9874 11508 9884
rect 11900 9604 11956 9614
rect 11340 9214 11342 9266
rect 11394 9214 11396 9266
rect 11340 9202 11396 9214
rect 11788 9602 11956 9604
rect 11788 9550 11902 9602
rect 11954 9550 11956 9602
rect 11788 9548 11956 9550
rect 9436 8932 9492 8988
rect 9660 8932 9716 8942
rect 9436 8930 9716 8932
rect 9436 8878 9662 8930
rect 9714 8878 9716 8930
rect 9436 8876 9716 8878
rect 9660 8708 9716 8876
rect 9660 8642 9716 8652
rect 9772 8148 9828 8158
rect 10780 8148 10836 8158
rect 9772 8146 10164 8148
rect 9772 8094 9774 8146
rect 9826 8094 10164 8146
rect 9772 8092 10164 8094
rect 9772 8082 9828 8092
rect 9324 7634 9380 7644
rect 10108 7698 10164 8092
rect 10108 7646 10110 7698
rect 10162 7646 10164 7698
rect 10108 7634 10164 7646
rect 10444 7476 10500 7486
rect 10444 7382 10500 7420
rect 8988 7298 9044 7308
rect 9100 7362 9156 7374
rect 9100 7310 9102 7362
rect 9154 7310 9156 7362
rect 8204 6738 8260 6748
rect 8428 6972 8932 7028
rect 8988 7028 9044 7038
rect 8092 6526 8094 6578
rect 8146 6526 8148 6578
rect 8092 6514 8148 6526
rect 7532 5124 7588 5134
rect 7532 5030 7588 5068
rect 8204 5124 8260 5134
rect 8204 5122 8372 5124
rect 8204 5070 8206 5122
rect 8258 5070 8372 5122
rect 8204 5068 8372 5070
rect 8204 5058 8260 5068
rect 7420 4946 7476 4956
rect 6748 4898 6804 4910
rect 6748 4846 6750 4898
rect 6802 4846 6804 4898
rect 6748 4452 6804 4846
rect 7644 4900 7700 4910
rect 6860 4452 6916 4462
rect 6748 4450 6916 4452
rect 6748 4398 6862 4450
rect 6914 4398 6916 4450
rect 6748 4396 6916 4398
rect 6860 4386 6916 4396
rect 7196 4004 7252 4014
rect 6972 3780 7028 3790
rect 6972 3554 7028 3724
rect 6972 3502 6974 3554
rect 7026 3502 7028 3554
rect 6972 3490 7028 3502
rect 7196 3442 7252 3948
rect 7644 3554 7700 4844
rect 7644 3502 7646 3554
rect 7698 3502 7700 3554
rect 7644 3490 7700 3502
rect 7756 4898 7812 4910
rect 7756 4846 7758 4898
rect 7810 4846 7812 4898
rect 7196 3390 7198 3442
rect 7250 3390 7252 3442
rect 7196 3378 7252 3390
rect 7756 2996 7812 4846
rect 8204 4340 8260 4350
rect 8204 3666 8260 4284
rect 8204 3614 8206 3666
rect 8258 3614 8260 3666
rect 8204 3602 8260 3614
rect 8316 3668 8372 5068
rect 8428 5010 8484 6972
rect 8540 6804 8596 6814
rect 8540 6580 8596 6748
rect 8540 6578 8708 6580
rect 8540 6526 8542 6578
rect 8594 6526 8708 6578
rect 8540 6524 8708 6526
rect 8540 6514 8596 6524
rect 8652 6130 8708 6524
rect 8988 6356 9044 6972
rect 9100 6692 9156 7310
rect 9772 7364 9828 7374
rect 9100 6636 9604 6692
rect 9212 6466 9268 6478
rect 9212 6414 9214 6466
rect 9266 6414 9268 6466
rect 8988 6300 9156 6356
rect 8652 6078 8654 6130
rect 8706 6078 8708 6130
rect 8652 6066 8708 6078
rect 8764 6244 8820 6254
rect 8428 4958 8430 5010
rect 8482 4958 8484 5010
rect 8428 4946 8484 4958
rect 8316 3602 8372 3612
rect 8764 3554 8820 6188
rect 8988 6132 9044 6142
rect 8876 5908 8932 5918
rect 8876 5122 8932 5852
rect 8876 5070 8878 5122
rect 8930 5070 8932 5122
rect 8876 5058 8932 5070
rect 8988 4226 9044 6076
rect 9100 5460 9156 6300
rect 9212 6244 9268 6414
rect 9212 6178 9268 6188
rect 9548 6466 9604 6636
rect 9548 6414 9550 6466
rect 9602 6414 9604 6466
rect 9548 5572 9604 6414
rect 9660 6580 9716 6590
rect 9660 5794 9716 6524
rect 9772 6468 9828 7308
rect 10220 6916 10276 6926
rect 9884 6692 9940 6702
rect 9884 6598 9940 6636
rect 10220 6578 10276 6860
rect 10668 6692 10724 6702
rect 10668 6598 10724 6636
rect 10220 6526 10222 6578
rect 10274 6526 10276 6578
rect 10220 6514 10276 6526
rect 9772 6412 9940 6468
rect 9660 5742 9662 5794
rect 9714 5742 9716 5794
rect 9660 5730 9716 5742
rect 9772 6018 9828 6030
rect 9772 5966 9774 6018
rect 9826 5966 9828 6018
rect 9772 5572 9828 5966
rect 9884 5908 9940 6412
rect 9996 6356 10052 6366
rect 9996 6018 10052 6300
rect 9996 5966 9998 6018
rect 10050 5966 10052 6018
rect 9996 5954 10052 5966
rect 10668 6018 10724 6030
rect 10668 5966 10670 6018
rect 10722 5966 10724 6018
rect 9884 5842 9940 5852
rect 10444 5906 10500 5918
rect 10444 5854 10446 5906
rect 10498 5854 10500 5906
rect 9548 5516 9716 5572
rect 9100 5404 9604 5460
rect 9548 5234 9604 5404
rect 9548 5182 9550 5234
rect 9602 5182 9604 5234
rect 9548 5170 9604 5182
rect 8988 4174 8990 4226
rect 9042 4174 9044 4226
rect 8988 4162 9044 4174
rect 9324 3668 9380 3678
rect 9324 3574 9380 3612
rect 8764 3502 8766 3554
rect 8818 3502 8820 3554
rect 8764 3490 8820 3502
rect 7868 3444 7924 3482
rect 7868 3378 7924 3388
rect 9660 3388 9716 5516
rect 9772 5506 9828 5516
rect 10444 5348 10500 5854
rect 10668 5460 10724 5966
rect 10668 5394 10724 5404
rect 10444 5282 10500 5292
rect 10444 5124 10500 5134
rect 10220 4340 10276 4350
rect 10220 4246 10276 4284
rect 10444 3388 10500 5068
rect 10556 4452 10612 4462
rect 10556 4358 10612 4396
rect 10668 4228 10724 4238
rect 10780 4228 10836 8092
rect 11788 7700 11844 9548
rect 11900 9538 11956 9548
rect 12348 9604 12404 9614
rect 12348 9510 12404 9548
rect 11900 8930 11956 8942
rect 11900 8878 11902 8930
rect 11954 8878 11956 8930
rect 11900 8596 11956 8878
rect 12124 8932 12180 8942
rect 12124 8930 12292 8932
rect 12124 8878 12126 8930
rect 12178 8878 12292 8930
rect 12124 8876 12292 8878
rect 12124 8866 12180 8876
rect 11900 8530 11956 8540
rect 11900 8372 11956 8382
rect 11900 8370 12180 8372
rect 11900 8318 11902 8370
rect 11954 8318 12180 8370
rect 11900 8316 12180 8318
rect 11900 8306 11956 8316
rect 11788 7644 11956 7700
rect 11228 7586 11284 7598
rect 11228 7534 11230 7586
rect 11282 7534 11284 7586
rect 11004 7476 11060 7486
rect 11004 7474 11172 7476
rect 11004 7422 11006 7474
rect 11058 7422 11172 7474
rect 11004 7420 11172 7422
rect 11004 7410 11060 7420
rect 11004 6690 11060 6702
rect 11004 6638 11006 6690
rect 11058 6638 11060 6690
rect 11004 6132 11060 6638
rect 11004 6066 11060 6076
rect 11004 5908 11060 5918
rect 11004 5814 11060 5852
rect 11116 4338 11172 7420
rect 11228 7364 11284 7534
rect 11340 7588 11396 7598
rect 11340 7586 11732 7588
rect 11340 7534 11342 7586
rect 11394 7534 11732 7586
rect 11340 7532 11732 7534
rect 11340 7522 11396 7532
rect 11228 7308 11396 7364
rect 11340 6692 11396 7308
rect 11116 4286 11118 4338
rect 11170 4286 11172 4338
rect 11116 4274 11172 4286
rect 11228 6580 11284 6590
rect 11340 6580 11396 6636
rect 11228 6578 11396 6580
rect 11228 6526 11230 6578
rect 11282 6526 11396 6578
rect 11228 6524 11396 6526
rect 11564 7252 11620 7262
rect 11564 6578 11620 7196
rect 11564 6526 11566 6578
rect 11618 6526 11620 6578
rect 11228 4340 11284 6524
rect 11564 6514 11620 6526
rect 11676 5234 11732 7532
rect 11788 7476 11844 7486
rect 11788 7382 11844 7420
rect 11788 6804 11844 6814
rect 11788 6018 11844 6748
rect 11788 5966 11790 6018
rect 11842 5966 11844 6018
rect 11788 5954 11844 5966
rect 11676 5182 11678 5234
rect 11730 5182 11732 5234
rect 11676 5170 11732 5182
rect 11788 5684 11844 5694
rect 11788 4564 11844 5628
rect 11788 4498 11844 4508
rect 11900 5012 11956 7644
rect 12124 7474 12180 8316
rect 12236 8148 12292 8876
rect 12460 8930 12516 10444
rect 12684 10164 12740 14254
rect 12796 13076 12852 15372
rect 13132 15092 13188 18284
rect 13804 18246 13860 18284
rect 13804 18004 13860 18014
rect 13692 17948 13804 18004
rect 13580 17780 13636 17790
rect 13580 17686 13636 17724
rect 13692 17554 13748 17948
rect 13804 17938 13860 17948
rect 13692 17502 13694 17554
rect 13746 17502 13748 17554
rect 13692 17490 13748 17502
rect 13804 17556 13860 17566
rect 13804 17462 13860 17500
rect 13916 17554 13972 18956
rect 14252 18452 14308 18462
rect 14252 18358 14308 18396
rect 14028 18228 14084 18238
rect 14028 18134 14084 18172
rect 13916 17502 13918 17554
rect 13970 17502 13972 17554
rect 13916 17490 13972 17502
rect 14252 17780 14308 17790
rect 13468 17444 13524 17454
rect 13468 17350 13524 17388
rect 13468 17220 13524 17230
rect 13468 17106 13524 17164
rect 13468 17054 13470 17106
rect 13522 17054 13524 17106
rect 13468 17042 13524 17054
rect 14028 17108 14084 17118
rect 14252 17108 14308 17724
rect 14028 17106 14308 17108
rect 14028 17054 14030 17106
rect 14082 17054 14254 17106
rect 14306 17054 14308 17106
rect 14028 17052 14308 17054
rect 14028 17042 14084 17052
rect 14252 15148 14308 17052
rect 14364 15316 14420 19068
rect 14588 17220 14644 21308
rect 14812 21298 14868 21308
rect 14924 22484 14980 22494
rect 14924 21924 14980 22428
rect 14812 20804 14868 20814
rect 14812 20710 14868 20748
rect 14700 20020 14756 20030
rect 14700 19926 14756 19964
rect 14924 19236 14980 21868
rect 16044 21476 16100 21486
rect 15260 21474 16100 21476
rect 15260 21422 16046 21474
rect 16098 21422 16100 21474
rect 15260 21420 16100 21422
rect 15148 21140 15204 21150
rect 15148 21026 15204 21084
rect 15148 20974 15150 21026
rect 15202 20974 15204 21026
rect 15148 20962 15204 20974
rect 15260 20914 15316 21420
rect 16044 21410 16100 21420
rect 15260 20862 15262 20914
rect 15314 20862 15316 20914
rect 15260 20850 15316 20862
rect 15148 20132 15204 20142
rect 15148 20038 15204 20076
rect 14812 19180 14980 19236
rect 15820 19684 15876 19694
rect 14700 18452 14756 18462
rect 14700 18358 14756 18396
rect 14812 18228 14868 19180
rect 15148 19124 15204 19134
rect 14924 19122 15204 19124
rect 14924 19070 15150 19122
rect 15202 19070 15204 19122
rect 14924 19068 15204 19070
rect 14924 18674 14980 19068
rect 15148 19058 15204 19068
rect 14924 18622 14926 18674
rect 14978 18622 14980 18674
rect 14924 18610 14980 18622
rect 14700 18172 14868 18228
rect 15260 18450 15316 18462
rect 15260 18398 15262 18450
rect 15314 18398 15316 18450
rect 14700 18004 14756 18172
rect 14700 17778 14756 17948
rect 14700 17726 14702 17778
rect 14754 17726 14756 17778
rect 14700 17714 14756 17726
rect 14588 17154 14644 17164
rect 14812 17668 14868 17678
rect 14588 16996 14644 17006
rect 14476 16940 14588 16996
rect 14476 15652 14532 16940
rect 14588 16902 14644 16940
rect 14700 16100 14756 16110
rect 14812 16100 14868 17612
rect 15260 16436 15316 18398
rect 15708 18452 15764 18462
rect 15708 18358 15764 18396
rect 15820 17892 15876 19628
rect 16156 18116 16212 25228
rect 16380 24164 16436 24174
rect 16380 23938 16436 24108
rect 16380 23886 16382 23938
rect 16434 23886 16436 23938
rect 16380 23874 16436 23886
rect 16268 23714 16324 23726
rect 16604 23716 16660 26126
rect 17052 24052 17108 28476
rect 17388 27860 17444 27870
rect 17276 27858 17444 27860
rect 17276 27806 17390 27858
rect 17442 27806 17444 27858
rect 17276 27804 17444 27806
rect 17164 26964 17220 27002
rect 17164 26898 17220 26908
rect 17276 24164 17332 27804
rect 17388 27794 17444 27804
rect 17500 27746 17556 27758
rect 17500 27694 17502 27746
rect 17554 27694 17556 27746
rect 17500 27298 17556 27694
rect 17612 27412 17668 37772
rect 17836 37044 17892 38612
rect 17724 34244 17780 34254
rect 17836 34244 17892 36988
rect 17948 35028 18004 39004
rect 18060 38836 18116 38846
rect 18060 38742 18116 38780
rect 18172 37492 18228 42700
rect 18396 42662 18452 42700
rect 18284 42084 18340 42094
rect 18284 40402 18340 42028
rect 18284 40350 18286 40402
rect 18338 40350 18340 40402
rect 18284 40338 18340 40350
rect 18396 41972 18452 41982
rect 18620 41972 18676 47292
rect 19292 47348 19348 47966
rect 19852 48020 19908 48302
rect 20076 48356 20132 48366
rect 20076 48242 20132 48300
rect 20076 48190 20078 48242
rect 20130 48190 20132 48242
rect 20076 48178 20132 48190
rect 19852 47954 19908 47964
rect 20748 48020 20804 48750
rect 20748 47954 20804 47964
rect 20972 48020 21028 48030
rect 21308 48020 21364 48030
rect 20972 48018 21140 48020
rect 20972 47966 20974 48018
rect 21026 47966 21140 48018
rect 20972 47964 21140 47966
rect 20972 47954 21028 47964
rect 21084 47460 21140 47964
rect 21308 47926 21364 47964
rect 21308 47460 21364 47470
rect 21084 47458 21364 47460
rect 21084 47406 21310 47458
rect 21362 47406 21364 47458
rect 21084 47404 21364 47406
rect 21308 47394 21364 47404
rect 19292 47282 19348 47292
rect 21420 47236 21476 48974
rect 21644 49026 21924 49028
rect 21644 48974 21870 49026
rect 21922 48974 21924 49026
rect 21644 48972 21924 48974
rect 21532 48356 21588 48366
rect 21532 48262 21588 48300
rect 21644 47346 21700 48972
rect 21868 48962 21924 48972
rect 24332 48802 24388 48814
rect 24332 48750 24334 48802
rect 24386 48750 24388 48802
rect 21980 48356 22036 48366
rect 21980 48262 22036 48300
rect 22652 48356 22708 48366
rect 24108 48356 24164 48366
rect 21644 47294 21646 47346
rect 21698 47294 21700 47346
rect 21644 47282 21700 47294
rect 21980 48020 22036 48030
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 18732 46116 18788 46126
rect 18732 43652 18788 46060
rect 19628 46116 19684 46126
rect 19628 46002 19684 46060
rect 19628 45950 19630 46002
rect 19682 45950 19684 46002
rect 19628 45938 19684 45950
rect 21196 46116 21252 46126
rect 21420 46116 21476 47180
rect 21252 46060 21476 46116
rect 20524 45892 20580 45902
rect 20748 45892 20804 45902
rect 21196 45892 21252 46060
rect 20524 45890 20692 45892
rect 20524 45838 20526 45890
rect 20578 45838 20692 45890
rect 20524 45836 20692 45838
rect 20524 45826 20580 45836
rect 19180 45668 19236 45678
rect 19180 45666 19348 45668
rect 19180 45614 19182 45666
rect 19234 45614 19348 45666
rect 19180 45612 19348 45614
rect 19180 45602 19236 45612
rect 19292 45444 19348 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19180 44884 19236 44894
rect 18732 43650 19012 43652
rect 18732 43598 18734 43650
rect 18786 43598 19012 43650
rect 18732 43596 19012 43598
rect 18732 43586 18788 43596
rect 18844 42868 18900 43596
rect 18956 43538 19012 43596
rect 18956 43486 18958 43538
rect 19010 43486 19012 43538
rect 18956 43474 19012 43486
rect 18844 42866 19012 42868
rect 18844 42814 18846 42866
rect 18898 42814 19012 42866
rect 18844 42812 19012 42814
rect 18844 42802 18900 42812
rect 18956 42196 19012 42812
rect 19180 42308 19236 44828
rect 19292 43652 19348 45388
rect 20636 44884 20692 45836
rect 20748 45778 20804 45836
rect 20748 45726 20750 45778
rect 20802 45726 20804 45778
rect 20748 45714 20804 45726
rect 20972 45890 21252 45892
rect 20972 45838 21198 45890
rect 21250 45838 21252 45890
rect 20972 45836 21252 45838
rect 20972 45330 21028 45836
rect 21196 45826 21252 45836
rect 21868 45892 21924 45902
rect 21868 45798 21924 45836
rect 21980 45668 22036 47964
rect 20972 45278 20974 45330
rect 21026 45278 21028 45330
rect 20748 44884 20804 44894
rect 20636 44882 20804 44884
rect 20636 44830 20750 44882
rect 20802 44830 20804 44882
rect 20636 44828 20804 44830
rect 20748 44818 20804 44828
rect 20972 44324 21028 45278
rect 21868 45612 22036 45668
rect 21084 44884 21140 44894
rect 21084 44882 21700 44884
rect 21084 44830 21086 44882
rect 21138 44830 21700 44882
rect 21084 44828 21700 44830
rect 21084 44818 21140 44828
rect 21644 44546 21700 44828
rect 21644 44494 21646 44546
rect 21698 44494 21700 44546
rect 21644 44482 21700 44494
rect 20972 44258 21028 44268
rect 20188 44210 20244 44222
rect 20188 44158 20190 44210
rect 20242 44158 20244 44210
rect 19852 44100 19908 44110
rect 19628 44098 19908 44100
rect 19628 44046 19854 44098
rect 19906 44046 19908 44098
rect 19628 44044 19908 44046
rect 19404 43652 19460 43662
rect 19292 43596 19404 43652
rect 19404 43586 19460 43596
rect 19628 43538 19684 44044
rect 19852 44034 19908 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19628 43486 19630 43538
rect 19682 43486 19684 43538
rect 19628 43474 19684 43486
rect 20188 42980 20244 44158
rect 20188 42914 20244 42924
rect 20412 43652 20468 43662
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19180 42252 19348 42308
rect 19836 42298 20100 42308
rect 18956 42194 19236 42196
rect 18956 42142 18958 42194
rect 19010 42142 19236 42194
rect 18956 42140 19236 42142
rect 18956 42130 19012 42140
rect 19180 41972 19236 42140
rect 18620 41916 19012 41972
rect 18396 38668 18452 41916
rect 18620 40180 18676 40190
rect 18620 40178 18788 40180
rect 18620 40126 18622 40178
rect 18674 40126 18788 40178
rect 18620 40124 18788 40126
rect 18620 40114 18676 40124
rect 18508 39060 18564 39070
rect 18508 38946 18564 39004
rect 18508 38894 18510 38946
rect 18562 38894 18564 38946
rect 18508 38882 18564 38894
rect 18620 38946 18676 38958
rect 18620 38894 18622 38946
rect 18674 38894 18676 38946
rect 18172 37156 18228 37436
rect 18284 38612 18452 38668
rect 18620 38724 18676 38894
rect 18620 38658 18676 38668
rect 18732 38668 18788 40124
rect 18844 38836 18900 38846
rect 18844 38742 18900 38780
rect 18732 38612 18900 38668
rect 18284 37378 18340 38612
rect 18284 37326 18286 37378
rect 18338 37326 18340 37378
rect 18284 37314 18340 37326
rect 18732 37826 18788 37838
rect 18732 37774 18734 37826
rect 18786 37774 18788 37826
rect 18732 37156 18788 37774
rect 18172 37100 18452 37156
rect 18284 36260 18340 36270
rect 17948 34356 18004 34972
rect 18172 35588 18228 35598
rect 18060 34916 18116 34926
rect 18060 34822 18116 34860
rect 18060 34356 18116 34366
rect 17948 34354 18116 34356
rect 17948 34302 18062 34354
rect 18114 34302 18116 34354
rect 17948 34300 18116 34302
rect 18060 34290 18116 34300
rect 17724 34242 17892 34244
rect 17724 34190 17726 34242
rect 17778 34190 17892 34242
rect 17724 34188 17892 34190
rect 17724 33458 17780 34188
rect 17724 33406 17726 33458
rect 17778 33406 17780 33458
rect 17724 32676 17780 33406
rect 18060 33572 18116 33582
rect 18172 33572 18228 35532
rect 18284 34914 18340 36204
rect 18396 35476 18452 37100
rect 18508 36372 18564 36382
rect 18508 36278 18564 36316
rect 18732 35924 18788 37100
rect 18844 36820 18900 38612
rect 18956 38050 19012 41916
rect 19180 41878 19236 41916
rect 19180 41300 19236 41310
rect 19292 41300 19348 42252
rect 19236 41244 19348 41300
rect 19628 41972 19684 41982
rect 19628 41298 19684 41916
rect 19964 41972 20020 41982
rect 19964 41970 20244 41972
rect 19964 41918 19966 41970
rect 20018 41918 20244 41970
rect 19964 41916 20244 41918
rect 19964 41906 20020 41916
rect 19628 41246 19630 41298
rect 19682 41246 19684 41298
rect 19180 41206 19236 41244
rect 19628 41234 19684 41246
rect 20188 41074 20244 41916
rect 20188 41022 20190 41074
rect 20242 41022 20244 41074
rect 20188 41010 20244 41022
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19180 40404 19236 40414
rect 19180 40310 19236 40348
rect 20188 40404 20244 40414
rect 19740 40290 19796 40302
rect 19740 40238 19742 40290
rect 19794 40238 19796 40290
rect 19180 40178 19236 40190
rect 19180 40126 19182 40178
rect 19234 40126 19236 40178
rect 19068 38612 19124 38622
rect 19068 38276 19124 38556
rect 19068 38210 19124 38220
rect 18956 37998 18958 38050
rect 19010 37998 19012 38050
rect 18956 37986 19012 37998
rect 19180 38052 19236 40126
rect 19740 40178 19796 40238
rect 19740 40126 19742 40178
rect 19794 40126 19796 40178
rect 19740 40114 19796 40126
rect 20188 39620 20244 40348
rect 19852 39396 19908 39406
rect 19628 39394 19908 39396
rect 19628 39342 19854 39394
rect 19906 39342 19908 39394
rect 19628 39340 19908 39342
rect 19628 38946 19684 39340
rect 19852 39330 19908 39340
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19628 38894 19630 38946
rect 19682 38894 19684 38946
rect 19628 38882 19684 38894
rect 19516 38836 19572 38846
rect 19516 38742 19572 38780
rect 20188 38834 20244 39564
rect 20188 38782 20190 38834
rect 20242 38782 20244 38834
rect 19292 38722 19348 38734
rect 19292 38670 19294 38722
rect 19346 38670 19348 38722
rect 19292 38612 19348 38670
rect 19292 38546 19348 38556
rect 20076 38612 20132 38622
rect 19740 38052 19796 38062
rect 19180 37958 19236 37996
rect 19628 38050 19796 38052
rect 19628 37998 19742 38050
rect 19794 37998 19796 38050
rect 19628 37996 19796 37998
rect 19628 37940 19684 37996
rect 19740 37986 19796 37996
rect 20076 38050 20132 38556
rect 20076 37998 20078 38050
rect 20130 37998 20132 38050
rect 19628 37874 19684 37884
rect 19404 37828 19460 37838
rect 19404 37734 19460 37772
rect 19516 37826 19572 37838
rect 19516 37774 19518 37826
rect 19570 37774 19572 37826
rect 19404 36932 19460 36942
rect 18844 36754 18900 36764
rect 19292 36820 19348 36830
rect 19068 36708 19124 36718
rect 18956 36372 19012 36382
rect 18956 36278 19012 36316
rect 18844 36260 18900 36270
rect 18844 36166 18900 36204
rect 18396 35410 18452 35420
rect 18620 35700 18676 35710
rect 18284 34862 18286 34914
rect 18338 34862 18340 34914
rect 18284 34850 18340 34862
rect 18620 34916 18676 35644
rect 18732 35698 18788 35868
rect 18732 35646 18734 35698
rect 18786 35646 18788 35698
rect 18732 35634 18788 35646
rect 18956 36148 19012 36158
rect 18844 35252 18900 35262
rect 18844 35138 18900 35196
rect 18844 35086 18846 35138
rect 18898 35086 18900 35138
rect 18844 35074 18900 35086
rect 18620 34356 18676 34860
rect 18956 34916 19012 36092
rect 19068 34916 19124 36652
rect 19292 34916 19348 36764
rect 19404 36482 19460 36876
rect 19404 36430 19406 36482
rect 19458 36430 19460 36482
rect 19404 36418 19460 36430
rect 19516 36484 19572 37774
rect 19852 37828 19908 37838
rect 19852 37734 19908 37772
rect 20076 37828 20132 37998
rect 20076 37762 20132 37772
rect 19628 37716 19684 37726
rect 19628 37156 19684 37660
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20076 37266 20132 37278
rect 20076 37214 20078 37266
rect 20130 37214 20132 37266
rect 20076 37156 20132 37214
rect 19628 37100 19908 37156
rect 19852 36706 19908 37100
rect 20076 37090 20132 37100
rect 19852 36654 19854 36706
rect 19906 36654 19908 36706
rect 19852 36642 19908 36654
rect 19516 36418 19572 36428
rect 19628 36596 19684 36606
rect 19628 36370 19684 36540
rect 19628 36318 19630 36370
rect 19682 36318 19684 36370
rect 19516 36258 19572 36270
rect 19516 36206 19518 36258
rect 19570 36206 19572 36258
rect 19516 35140 19572 36206
rect 19628 35700 19684 36318
rect 19964 36482 20020 36494
rect 19964 36430 19966 36482
rect 20018 36430 20020 36482
rect 19964 36260 20020 36430
rect 19964 36194 20020 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19628 35634 19684 35644
rect 20188 35588 20244 38782
rect 20412 38668 20468 43596
rect 21420 42980 21476 42990
rect 21420 42886 21476 42924
rect 21756 42754 21812 42766
rect 21756 42702 21758 42754
rect 21810 42702 21812 42754
rect 21756 41860 21812 42702
rect 21756 41794 21812 41804
rect 21756 41186 21812 41198
rect 21756 41134 21758 41186
rect 21810 41134 21812 41186
rect 20524 41076 20580 41086
rect 21420 41076 21476 41086
rect 20524 41074 21476 41076
rect 20524 41022 20526 41074
rect 20578 41022 21422 41074
rect 21474 41022 21476 41074
rect 20524 41020 21476 41022
rect 20524 41010 20580 41020
rect 21420 41010 21476 41020
rect 21756 40964 21812 41134
rect 21756 40898 21812 40908
rect 20972 40290 21028 40302
rect 21756 40292 21812 40302
rect 20972 40238 20974 40290
rect 21026 40238 21028 40290
rect 20524 39618 20580 39630
rect 20524 39566 20526 39618
rect 20578 39566 20580 39618
rect 20524 39508 20580 39566
rect 20636 39508 20692 39518
rect 20524 39452 20636 39508
rect 20636 39442 20692 39452
rect 20748 39394 20804 39406
rect 20748 39342 20750 39394
rect 20802 39342 20804 39394
rect 20748 38834 20804 39342
rect 20748 38782 20750 38834
rect 20802 38782 20804 38834
rect 20748 38770 20804 38782
rect 20412 38612 20580 38668
rect 20412 37940 20468 37950
rect 20412 37846 20468 37884
rect 20524 37938 20580 38612
rect 20524 37886 20526 37938
rect 20578 37886 20580 37938
rect 20524 37874 20580 37886
rect 20972 38612 21028 40238
rect 20972 37940 21028 38556
rect 20748 37826 20804 37838
rect 20748 37774 20750 37826
rect 20802 37774 20804 37826
rect 20188 35494 20244 35532
rect 20300 37716 20356 37726
rect 19516 35074 19572 35084
rect 20188 35140 20244 35150
rect 20188 35046 20244 35084
rect 19740 34916 19796 34926
rect 19068 34860 19236 34916
rect 19292 34914 19796 34916
rect 19292 34862 19742 34914
rect 19794 34862 19796 34914
rect 19292 34860 19796 34862
rect 18956 34822 19012 34860
rect 18620 34290 18676 34300
rect 19068 34690 19124 34702
rect 19068 34638 19070 34690
rect 19122 34638 19124 34690
rect 18396 34130 18452 34142
rect 18396 34078 18398 34130
rect 18450 34078 18452 34130
rect 18060 33570 18228 33572
rect 18060 33518 18062 33570
rect 18114 33518 18228 33570
rect 18060 33516 18228 33518
rect 18284 33570 18340 33582
rect 18284 33518 18286 33570
rect 18338 33518 18340 33570
rect 17724 32610 17780 32620
rect 17836 33124 17892 33134
rect 17724 31668 17780 31678
rect 17724 31106 17780 31612
rect 17724 31054 17726 31106
rect 17778 31054 17780 31106
rect 17724 31042 17780 31054
rect 17836 30884 17892 33068
rect 17948 32562 18004 32574
rect 17948 32510 17950 32562
rect 18002 32510 18004 32562
rect 17948 32452 18004 32510
rect 17948 32386 18004 32396
rect 18060 32340 18116 33516
rect 18172 33124 18228 33134
rect 18284 33124 18340 33518
rect 18172 33122 18340 33124
rect 18172 33070 18174 33122
rect 18226 33070 18340 33122
rect 18172 33068 18340 33070
rect 18396 33124 18452 34078
rect 18732 34130 18788 34142
rect 18732 34078 18734 34130
rect 18786 34078 18788 34130
rect 18732 33570 18788 34078
rect 18956 34132 19012 34142
rect 19068 34132 19124 34638
rect 19180 34356 19236 34860
rect 19740 34850 19796 34860
rect 20076 34916 20132 34926
rect 20076 34914 20244 34916
rect 20076 34862 20078 34914
rect 20130 34862 20244 34914
rect 20076 34860 20244 34862
rect 20076 34850 20132 34860
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19180 34300 19348 34356
rect 19180 34132 19236 34142
rect 19068 34130 19236 34132
rect 19068 34078 19182 34130
rect 19234 34078 19236 34130
rect 19068 34076 19236 34078
rect 18956 34038 19012 34076
rect 19180 34066 19236 34076
rect 18732 33518 18734 33570
rect 18786 33518 18788 33570
rect 18732 33506 18788 33518
rect 19292 33348 19348 34300
rect 19516 34354 19572 34366
rect 19516 34302 19518 34354
rect 19570 34302 19572 34354
rect 19404 34130 19460 34142
rect 19404 34078 19406 34130
rect 19458 34078 19460 34130
rect 19404 33458 19460 34078
rect 19516 33572 19572 34302
rect 19964 34020 20020 34030
rect 20188 34020 20244 34860
rect 20020 33964 20244 34020
rect 19964 33926 20020 33964
rect 19516 33506 19572 33516
rect 19404 33406 19406 33458
rect 19458 33406 19460 33458
rect 19404 33394 19460 33406
rect 19180 33292 19348 33348
rect 19516 33348 19572 33358
rect 18620 33124 18676 33134
rect 18396 33122 18676 33124
rect 18396 33070 18622 33122
rect 18674 33070 18676 33122
rect 18396 33068 18676 33070
rect 18172 33058 18228 33068
rect 18172 32340 18228 32350
rect 18060 32338 18228 32340
rect 18060 32286 18174 32338
rect 18226 32286 18228 32338
rect 18060 32284 18228 32286
rect 18060 31780 18116 32284
rect 18172 32274 18228 32284
rect 18284 32116 18340 33068
rect 18396 32450 18452 32462
rect 18396 32398 18398 32450
rect 18450 32398 18452 32450
rect 18396 32338 18452 32398
rect 18396 32286 18398 32338
rect 18450 32286 18452 32338
rect 18396 32274 18452 32286
rect 18284 32060 18452 32116
rect 17948 31556 18004 31566
rect 17948 31106 18004 31500
rect 17948 31054 17950 31106
rect 18002 31054 18004 31106
rect 17948 31042 18004 31054
rect 17724 30828 17892 30884
rect 18060 30884 18116 31724
rect 18284 31780 18340 31790
rect 18172 31556 18228 31566
rect 18284 31556 18340 31724
rect 18396 31668 18452 32060
rect 18508 31892 18564 31902
rect 18508 31798 18564 31836
rect 18396 31612 18564 31668
rect 18172 31554 18340 31556
rect 18172 31502 18174 31554
rect 18226 31502 18340 31554
rect 18172 31500 18340 31502
rect 18172 31490 18228 31500
rect 17724 30548 17780 30828
rect 18060 30818 18116 30828
rect 17724 30098 17780 30492
rect 17724 30046 17726 30098
rect 17778 30046 17780 30098
rect 17724 30034 17780 30046
rect 18060 29988 18116 29998
rect 18060 29986 18228 29988
rect 18060 29934 18062 29986
rect 18114 29934 18228 29986
rect 18060 29932 18228 29934
rect 18060 29922 18116 29932
rect 18172 29540 18228 29932
rect 18172 29426 18228 29484
rect 18172 29374 18174 29426
rect 18226 29374 18228 29426
rect 17836 29316 17892 29326
rect 17836 28868 17892 29260
rect 17836 28812 18116 28868
rect 17724 28084 17780 28094
rect 17724 27858 17780 28028
rect 17724 27806 17726 27858
rect 17778 27806 17780 27858
rect 17724 27794 17780 27806
rect 17836 27746 17892 27758
rect 17836 27694 17838 27746
rect 17890 27694 17892 27746
rect 17724 27636 17780 27646
rect 17836 27636 17892 27694
rect 17780 27580 17892 27636
rect 17724 27570 17780 27580
rect 17612 27356 18004 27412
rect 17500 27246 17502 27298
rect 17554 27246 17556 27298
rect 17500 27234 17556 27246
rect 17612 27188 17668 27198
rect 17500 26964 17556 26974
rect 17388 26180 17444 26190
rect 17388 25284 17444 26124
rect 17388 25218 17444 25228
rect 17500 24948 17556 26908
rect 17612 26290 17668 27132
rect 17724 27076 17780 27114
rect 17724 27010 17780 27020
rect 17724 26852 17780 26862
rect 17724 26850 17892 26852
rect 17724 26798 17726 26850
rect 17778 26798 17892 26850
rect 17724 26796 17892 26798
rect 17724 26786 17780 26796
rect 17612 26238 17614 26290
rect 17666 26238 17668 26290
rect 17612 26226 17668 26238
rect 17836 26290 17892 26796
rect 17836 26238 17838 26290
rect 17890 26238 17892 26290
rect 17836 26226 17892 26238
rect 17948 25732 18004 27356
rect 17724 25676 18004 25732
rect 17724 25060 17780 25676
rect 18060 25620 18116 28812
rect 18172 28530 18228 29374
rect 18172 28478 18174 28530
rect 18226 28478 18228 28530
rect 18172 27858 18228 28478
rect 18172 27806 18174 27858
rect 18226 27806 18228 27858
rect 18172 27794 18228 27806
rect 18284 27636 18340 31500
rect 18508 30996 18564 31612
rect 18620 31220 18676 33068
rect 19180 32900 19236 33292
rect 19516 33254 19572 33292
rect 19964 33346 20020 33358
rect 19964 33294 19966 33346
rect 20018 33294 20020 33346
rect 19292 33124 19348 33134
rect 19964 33124 20020 33294
rect 20300 33348 20356 37660
rect 20636 37154 20692 37166
rect 20636 37102 20638 37154
rect 20690 37102 20692 37154
rect 20636 36596 20692 37102
rect 20636 36530 20692 36540
rect 20748 36484 20804 37774
rect 20972 37044 21028 37884
rect 21420 40290 21812 40292
rect 21420 40238 21758 40290
rect 21810 40238 21812 40290
rect 21420 40236 21812 40238
rect 21420 37828 21476 40236
rect 21756 40226 21812 40236
rect 21756 39508 21812 39518
rect 21756 39414 21812 39452
rect 21644 39284 21700 39294
rect 21868 39284 21924 45612
rect 21980 44322 22036 44334
rect 21980 44270 21982 44322
rect 22034 44270 22036 44322
rect 21980 43428 22036 44270
rect 22428 44322 22484 44334
rect 22428 44270 22430 44322
rect 22482 44270 22484 44322
rect 22092 43428 22148 43438
rect 21980 43372 22092 43428
rect 22092 43334 22148 43372
rect 22204 42756 22260 42766
rect 22428 42756 22484 44270
rect 22204 42754 22484 42756
rect 22204 42702 22206 42754
rect 22258 42702 22484 42754
rect 22204 42700 22484 42702
rect 22540 43428 22596 43438
rect 22204 41188 22260 42700
rect 22540 42642 22596 43372
rect 22540 42590 22542 42642
rect 22594 42590 22596 42642
rect 22316 41860 22372 41870
rect 22372 41804 22484 41860
rect 22316 41766 22372 41804
rect 22204 41186 22372 41188
rect 22204 41134 22206 41186
rect 22258 41134 22372 41186
rect 22204 41132 22372 41134
rect 22204 41122 22260 41132
rect 22092 39620 22148 39630
rect 22092 39526 22148 39564
rect 22316 39508 22372 41132
rect 22428 41074 22484 41804
rect 22428 41022 22430 41074
rect 22482 41022 22484 41074
rect 22428 40852 22484 41022
rect 22428 40786 22484 40796
rect 22316 39506 22484 39508
rect 22316 39454 22318 39506
rect 22370 39454 22484 39506
rect 22316 39452 22484 39454
rect 22316 39442 22372 39452
rect 21868 39228 22372 39284
rect 21644 38164 21700 39228
rect 21644 38070 21700 38108
rect 21868 39060 21924 39070
rect 21756 37828 21812 37838
rect 21420 37772 21756 37828
rect 21308 37156 21364 37166
rect 21308 37062 21364 37100
rect 20972 36978 21028 36988
rect 20748 36418 20804 36428
rect 21532 36482 21588 36494
rect 21532 36430 21534 36482
rect 21586 36430 21588 36482
rect 21420 36372 21476 36382
rect 21420 36278 21476 36316
rect 20860 36260 20916 36270
rect 20748 36204 20860 36260
rect 20524 34916 20580 34926
rect 20524 34914 20692 34916
rect 20524 34862 20526 34914
rect 20578 34862 20692 34914
rect 20524 34860 20692 34862
rect 20524 34850 20580 34860
rect 20524 34690 20580 34702
rect 20524 34638 20526 34690
rect 20578 34638 20580 34690
rect 20524 33460 20580 34638
rect 20636 34468 20692 34860
rect 20636 34354 20692 34412
rect 20636 34302 20638 34354
rect 20690 34302 20692 34354
rect 20636 34290 20692 34302
rect 20524 33394 20580 33404
rect 20300 33282 20356 33292
rect 20412 33124 20468 33134
rect 19964 33122 20468 33124
rect 19964 33070 20414 33122
rect 20466 33070 20468 33122
rect 19964 33068 20468 33070
rect 19292 33030 19348 33068
rect 19836 32956 20100 32966
rect 19180 32834 19236 32844
rect 19628 32900 19684 32910
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32900 20244 32910
rect 18844 32452 18900 32462
rect 18844 32358 18900 32396
rect 19516 32340 19572 32350
rect 19404 32338 19572 32340
rect 19404 32286 19518 32338
rect 19570 32286 19572 32338
rect 19404 32284 19572 32286
rect 18844 31890 18900 31902
rect 18844 31838 18846 31890
rect 18898 31838 18900 31890
rect 18732 31780 18788 31790
rect 18732 31666 18788 31724
rect 18732 31614 18734 31666
rect 18786 31614 18788 31666
rect 18732 31332 18788 31614
rect 18844 31556 18900 31838
rect 18844 31490 18900 31500
rect 19404 31556 19460 32284
rect 19516 32274 19572 32284
rect 19628 31778 19684 32844
rect 20412 32900 20468 33068
rect 20412 32844 20692 32900
rect 20188 32788 20244 32844
rect 20076 32732 20244 32788
rect 19740 32450 19796 32462
rect 19740 32398 19742 32450
rect 19794 32398 19796 32450
rect 19740 32338 19796 32398
rect 19740 32286 19742 32338
rect 19794 32286 19796 32338
rect 19740 32274 19796 32286
rect 20076 32338 20132 32732
rect 20524 32676 20580 32686
rect 20412 32674 20580 32676
rect 20412 32622 20526 32674
rect 20578 32622 20580 32674
rect 20412 32620 20580 32622
rect 20300 32452 20356 32462
rect 20076 32286 20078 32338
rect 20130 32286 20132 32338
rect 20076 32274 20132 32286
rect 20188 32450 20356 32452
rect 20188 32398 20302 32450
rect 20354 32398 20356 32450
rect 20188 32396 20356 32398
rect 20188 32116 20244 32396
rect 20300 32386 20356 32396
rect 19628 31726 19630 31778
rect 19682 31726 19684 31778
rect 19628 31668 19684 31726
rect 19964 32060 20244 32116
rect 19964 31780 20020 32060
rect 20412 31892 20468 32620
rect 20524 32610 20580 32620
rect 20636 32228 20692 32844
rect 20636 32162 20692 32172
rect 19964 31686 20020 31724
rect 20300 31836 20468 31892
rect 19628 31602 19684 31612
rect 19404 31462 19460 31500
rect 19516 31554 19572 31566
rect 19516 31502 19518 31554
rect 19570 31502 19572 31554
rect 18732 31276 18900 31332
rect 18620 31164 18788 31220
rect 18620 30996 18676 31006
rect 18508 30994 18676 30996
rect 18508 30942 18622 30994
rect 18674 30942 18676 30994
rect 18508 30940 18676 30942
rect 18732 30996 18788 31164
rect 18844 31108 18900 31276
rect 19068 31218 19124 31230
rect 19516 31220 19572 31502
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19068 31166 19070 31218
rect 19122 31166 19124 31218
rect 18844 31052 19012 31108
rect 18732 30940 18900 30996
rect 18508 29988 18564 29998
rect 18620 29988 18676 30940
rect 18844 30772 18900 30940
rect 18956 30994 19012 31052
rect 18956 30942 18958 30994
rect 19010 30942 19012 30994
rect 18956 30930 19012 30942
rect 18508 29986 18676 29988
rect 18508 29934 18510 29986
rect 18562 29934 18676 29986
rect 18508 29932 18676 29934
rect 18732 30716 18900 30772
rect 18396 29092 18452 29102
rect 18396 28642 18452 29036
rect 18396 28590 18398 28642
rect 18450 28590 18452 28642
rect 18396 28578 18452 28590
rect 18508 28420 18564 29932
rect 18620 29540 18676 29550
rect 18620 29446 18676 29484
rect 18508 28354 18564 28364
rect 18620 28084 18676 28094
rect 18620 27990 18676 28028
rect 18060 25284 18116 25564
rect 18172 27580 18340 27636
rect 18508 27748 18564 27758
rect 18172 25396 18228 27580
rect 18508 26514 18564 27692
rect 18508 26462 18510 26514
rect 18562 26462 18564 26514
rect 18508 26450 18564 26462
rect 18284 26066 18340 26078
rect 18284 26014 18286 26066
rect 18338 26014 18340 26066
rect 18284 25956 18340 26014
rect 18284 25890 18340 25900
rect 18284 25732 18340 25742
rect 18284 25730 18676 25732
rect 18284 25678 18286 25730
rect 18338 25678 18676 25730
rect 18284 25676 18676 25678
rect 18284 25666 18340 25676
rect 18396 25508 18452 25518
rect 18396 25414 18452 25452
rect 18620 25506 18676 25676
rect 18732 25620 18788 30716
rect 19068 30660 19124 31166
rect 19404 31164 19572 31220
rect 19404 30994 19460 31164
rect 19404 30942 19406 30994
rect 19458 30942 19460 30994
rect 19404 30930 19460 30942
rect 19740 30994 19796 31006
rect 19740 30942 19742 30994
rect 19794 30942 19796 30994
rect 19740 30884 19796 30942
rect 20300 30994 20356 31836
rect 20412 31668 20468 31678
rect 20412 31574 20468 31612
rect 20636 31668 20692 31678
rect 20300 30942 20302 30994
rect 20354 30942 20356 30994
rect 20300 30930 20356 30942
rect 20524 31554 20580 31566
rect 20524 31502 20526 31554
rect 20578 31502 20580 31554
rect 19180 30772 19236 30782
rect 19180 30770 19572 30772
rect 19180 30718 19182 30770
rect 19234 30718 19572 30770
rect 19180 30716 19572 30718
rect 19180 30706 19236 30716
rect 19068 30594 19124 30604
rect 19516 30324 19572 30716
rect 19628 30324 19684 30334
rect 19516 30322 19684 30324
rect 19516 30270 19630 30322
rect 19682 30270 19684 30322
rect 19516 30268 19684 30270
rect 19628 30258 19684 30268
rect 19740 30324 19796 30828
rect 20524 30772 20580 31502
rect 20076 30716 20580 30772
rect 20076 30434 20132 30716
rect 20076 30382 20078 30434
rect 20130 30382 20132 30434
rect 20076 30370 20132 30382
rect 19740 30258 19796 30268
rect 19404 30212 19460 30222
rect 18844 29988 18900 29998
rect 18844 28084 18900 29932
rect 19180 29540 19236 29550
rect 19180 29446 19236 29484
rect 18844 28018 18900 28028
rect 18956 28868 19012 28878
rect 18732 25554 18788 25564
rect 18844 26402 18900 26414
rect 18844 26350 18846 26402
rect 18898 26350 18900 26402
rect 18620 25454 18622 25506
rect 18674 25454 18676 25506
rect 18620 25442 18676 25454
rect 18284 25396 18340 25406
rect 18172 25394 18340 25396
rect 18172 25342 18286 25394
rect 18338 25342 18340 25394
rect 18172 25340 18340 25342
rect 18284 25330 18340 25340
rect 18844 25396 18900 26350
rect 18844 25330 18900 25340
rect 18060 25228 18228 25284
rect 18060 25060 18116 25070
rect 17724 25004 18004 25060
rect 17500 24892 17780 24948
rect 17500 24722 17556 24734
rect 17500 24670 17502 24722
rect 17554 24670 17556 24722
rect 17276 24108 17444 24164
rect 17052 23996 17332 24052
rect 16268 23662 16270 23714
rect 16322 23662 16324 23714
rect 16268 22148 16324 23662
rect 16268 22082 16324 22092
rect 16380 23660 16660 23716
rect 16716 23826 16772 23838
rect 17052 23828 17108 23838
rect 16716 23774 16718 23826
rect 16770 23774 16772 23826
rect 16380 20020 16436 23660
rect 16716 23604 16772 23774
rect 16716 23538 16772 23548
rect 16828 23826 17108 23828
rect 16828 23774 17054 23826
rect 17106 23774 17108 23826
rect 16828 23772 17108 23774
rect 16828 23378 16884 23772
rect 17052 23762 17108 23772
rect 17164 23716 17220 23726
rect 17164 23622 17220 23660
rect 16828 23326 16830 23378
rect 16882 23326 16884 23378
rect 16828 23314 16884 23326
rect 16940 23156 16996 23166
rect 16492 22372 16548 22382
rect 16940 22372 16996 23100
rect 16548 22370 16996 22372
rect 16548 22318 16942 22370
rect 16994 22318 16996 22370
rect 16548 22316 16996 22318
rect 16492 21810 16548 22316
rect 16940 22306 16996 22316
rect 16492 21758 16494 21810
rect 16546 21758 16548 21810
rect 16492 21746 16548 21758
rect 16828 21588 16884 21598
rect 16828 21586 17108 21588
rect 16828 21534 16830 21586
rect 16882 21534 17108 21586
rect 16828 21532 17108 21534
rect 16828 21522 16884 21532
rect 17052 20580 17108 21532
rect 17052 20486 17108 20524
rect 16380 19954 16436 19964
rect 16828 20018 16884 20030
rect 16828 19966 16830 20018
rect 16882 19966 16884 20018
rect 16156 18050 16212 18060
rect 16268 19906 16324 19918
rect 16268 19854 16270 19906
rect 16322 19854 16324 19906
rect 15820 17826 15876 17836
rect 16044 17892 16100 17902
rect 16268 17892 16324 19854
rect 16828 19348 16884 19966
rect 17276 19572 17332 23996
rect 17388 23716 17444 24108
rect 17388 23650 17444 23660
rect 17500 23380 17556 24670
rect 17724 23828 17780 24892
rect 17612 23716 17668 23726
rect 17612 23622 17668 23660
rect 17388 23156 17444 23166
rect 17388 23062 17444 23100
rect 17500 22820 17556 23324
rect 17500 22754 17556 22764
rect 17388 22484 17444 22494
rect 17388 22390 17444 22428
rect 17724 22482 17780 23772
rect 17948 23492 18004 25004
rect 18060 24722 18116 25004
rect 18060 24670 18062 24722
rect 18114 24670 18116 24722
rect 18060 24658 18116 24670
rect 18172 24388 18228 25228
rect 18172 24322 18228 24332
rect 17948 23154 18004 23436
rect 17948 23102 17950 23154
rect 18002 23102 18004 23154
rect 17948 23090 18004 23102
rect 18172 23268 18228 23278
rect 17724 22430 17726 22482
rect 17778 22430 17780 22482
rect 17724 22418 17780 22430
rect 18172 22260 18228 23212
rect 18956 23156 19012 28812
rect 19292 28644 19348 28654
rect 19068 28084 19124 28094
rect 19068 27858 19124 28028
rect 19068 27806 19070 27858
rect 19122 27806 19124 27858
rect 19068 27794 19124 27806
rect 19292 26908 19348 28588
rect 19404 28084 19460 30156
rect 19852 30210 19908 30222
rect 19852 30158 19854 30210
rect 19906 30158 19908 30210
rect 19516 30100 19572 30110
rect 19516 30098 19684 30100
rect 19516 30046 19518 30098
rect 19570 30046 19684 30098
rect 19516 30044 19684 30046
rect 19516 30034 19572 30044
rect 19404 28018 19460 28028
rect 19516 28868 19572 28878
rect 19516 28642 19572 28812
rect 19516 28590 19518 28642
rect 19570 28590 19572 28642
rect 19516 27860 19572 28590
rect 19628 28644 19684 30044
rect 19852 29988 19908 30158
rect 20076 30212 20132 30222
rect 20076 30118 20132 30156
rect 19852 29922 19908 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20412 28754 20468 28766
rect 20412 28702 20414 28754
rect 20466 28702 20468 28754
rect 19740 28644 19796 28654
rect 19628 28588 19740 28644
rect 19740 28550 19796 28588
rect 20076 28644 20132 28654
rect 20412 28644 20468 28702
rect 20076 28642 20468 28644
rect 20076 28590 20078 28642
rect 20130 28590 20468 28642
rect 20076 28588 20468 28590
rect 20076 28578 20132 28588
rect 20524 28530 20580 28542
rect 20524 28478 20526 28530
rect 20578 28478 20580 28530
rect 19292 26852 19460 26908
rect 19292 26180 19348 26190
rect 19292 26086 19348 26124
rect 19404 25620 19460 26852
rect 19516 26290 19572 27804
rect 19628 28418 19684 28430
rect 19628 28366 19630 28418
rect 19682 28366 19684 28418
rect 19628 27858 19684 28366
rect 20524 28420 20580 28478
rect 20636 28420 20692 31612
rect 20748 28756 20804 36204
rect 20860 36166 20916 36204
rect 21084 35588 21140 35598
rect 21084 34356 21140 35532
rect 21532 34468 21588 36430
rect 21644 35924 21700 35934
rect 21644 35830 21700 35868
rect 21532 34402 21588 34412
rect 21644 35700 21700 35710
rect 21644 35026 21700 35644
rect 21644 34974 21646 35026
rect 21698 34974 21700 35026
rect 21084 34354 21364 34356
rect 21084 34302 21086 34354
rect 21138 34302 21364 34354
rect 21084 34300 21364 34302
rect 21084 34290 21140 34300
rect 21308 34130 21364 34300
rect 21308 34078 21310 34130
rect 21362 34078 21364 34130
rect 21308 34066 21364 34078
rect 20860 33122 20916 33134
rect 20860 33070 20862 33122
rect 20914 33070 20916 33122
rect 20860 32900 20916 33070
rect 20860 32834 20916 32844
rect 21308 32900 21364 32910
rect 20860 32564 20916 32574
rect 20860 32562 21140 32564
rect 20860 32510 20862 32562
rect 20914 32510 21140 32562
rect 20860 32508 21140 32510
rect 20860 32498 20916 32508
rect 21084 32004 21140 32508
rect 21308 32452 21364 32844
rect 21308 32358 21364 32396
rect 21532 32004 21588 32014
rect 21084 32002 21588 32004
rect 21084 31950 21534 32002
rect 21586 31950 21588 32002
rect 21084 31948 21588 31950
rect 21532 31938 21588 31948
rect 20860 29988 20916 29998
rect 20860 29894 20916 29932
rect 21644 29540 21700 34974
rect 21756 32564 21812 37772
rect 21868 35700 21924 39004
rect 22204 38052 22260 38062
rect 21980 37828 22036 37838
rect 21980 37734 22036 37772
rect 22204 37266 22260 37996
rect 22204 37214 22206 37266
rect 22258 37214 22260 37266
rect 22204 37202 22260 37214
rect 22316 37154 22372 39228
rect 22428 38162 22484 39452
rect 22428 38110 22430 38162
rect 22482 38110 22484 38162
rect 22428 38098 22484 38110
rect 22540 37156 22596 42590
rect 22652 39060 22708 48300
rect 23996 48354 24164 48356
rect 23996 48302 24110 48354
rect 24162 48302 24164 48354
rect 23996 48300 24164 48302
rect 23212 47458 23268 47470
rect 23212 47406 23214 47458
rect 23266 47406 23268 47458
rect 22988 47236 23044 47246
rect 23212 47236 23268 47406
rect 23996 47458 24052 48300
rect 24108 48290 24164 48300
rect 24332 48356 24388 48750
rect 25564 48804 25620 48814
rect 25564 48802 25732 48804
rect 25564 48750 25566 48802
rect 25618 48750 25732 48802
rect 25564 48748 25732 48750
rect 25564 48738 25620 48748
rect 24332 48290 24388 48300
rect 25676 48356 25732 48748
rect 27356 48466 27412 49756
rect 27916 49026 27972 50318
rect 29484 49922 29540 49934
rect 29484 49870 29486 49922
rect 29538 49870 29540 49922
rect 28924 49698 28980 49710
rect 28924 49646 28926 49698
rect 28978 49646 28980 49698
rect 27916 48974 27918 49026
rect 27970 48974 27972 49026
rect 27916 48962 27972 48974
rect 28700 49028 28756 49038
rect 28924 49028 28980 49646
rect 28700 49026 28980 49028
rect 28700 48974 28702 49026
rect 28754 48974 28980 49026
rect 28700 48972 28980 48974
rect 29260 49028 29316 49038
rect 29484 49028 29540 49870
rect 32844 49922 32900 49934
rect 32844 49870 32846 49922
rect 32898 49870 32900 49922
rect 29820 49810 29876 49822
rect 29820 49758 29822 49810
rect 29874 49758 29876 49810
rect 29708 49028 29764 49038
rect 29484 49026 29764 49028
rect 29484 48974 29710 49026
rect 29762 48974 29764 49026
rect 29484 48972 29764 48974
rect 27356 48414 27358 48466
rect 27410 48414 27412 48466
rect 27356 48402 27412 48414
rect 23996 47406 23998 47458
rect 24050 47406 24052 47458
rect 23996 47394 24052 47406
rect 24444 48242 24500 48254
rect 24444 48190 24446 48242
rect 24498 48190 24500 48242
rect 23044 47180 23268 47236
rect 22988 47142 23044 47180
rect 24444 46900 24500 48190
rect 24444 46834 24500 46844
rect 25340 46900 25396 46910
rect 25340 46806 25396 46844
rect 25676 46450 25732 48300
rect 28252 48356 28308 48366
rect 28252 48262 28308 48300
rect 28476 48242 28532 48254
rect 28476 48190 28478 48242
rect 28530 48190 28532 48242
rect 26908 48132 26964 48142
rect 26348 47234 26404 47246
rect 26348 47182 26350 47234
rect 26402 47182 26404 47234
rect 26348 46786 26404 47182
rect 26348 46734 26350 46786
rect 26402 46734 26404 46786
rect 25676 46398 25678 46450
rect 25730 46398 25732 46450
rect 25004 45780 25060 45790
rect 25004 45778 25172 45780
rect 25004 45726 25006 45778
rect 25058 45726 25172 45778
rect 25004 45724 25172 45726
rect 25004 45714 25060 45724
rect 22764 45668 22820 45678
rect 22764 44210 22820 45612
rect 24332 45668 24388 45678
rect 24668 45668 24724 45678
rect 24332 45574 24388 45612
rect 24444 45666 24724 45668
rect 24444 45614 24670 45666
rect 24722 45614 24724 45666
rect 24444 45612 24724 45614
rect 23324 44324 23380 44334
rect 24108 44324 24164 44334
rect 24444 44324 24500 45612
rect 24668 45602 24724 45612
rect 25116 45332 25172 45724
rect 25676 45668 25732 46398
rect 26124 46674 26180 46686
rect 26124 46622 26126 46674
rect 26178 46622 26180 46674
rect 25676 45612 26068 45668
rect 25340 45332 25396 45342
rect 25116 45330 25396 45332
rect 25116 45278 25342 45330
rect 25394 45278 25396 45330
rect 25116 45276 25396 45278
rect 25340 45266 25396 45276
rect 25676 44884 25732 44894
rect 25788 44884 25844 44894
rect 25676 44882 25788 44884
rect 25676 44830 25678 44882
rect 25730 44830 25788 44882
rect 25676 44828 25788 44830
rect 25676 44818 25732 44828
rect 22764 44158 22766 44210
rect 22818 44158 22820 44210
rect 22764 39620 22820 44158
rect 23100 44268 23324 44324
rect 23380 44268 23492 44324
rect 23100 43764 23156 44268
rect 23324 44230 23380 44268
rect 22988 43762 23156 43764
rect 22988 43710 23102 43762
rect 23154 43710 23156 43762
rect 22988 43708 23156 43710
rect 22988 40628 23044 43708
rect 23100 43698 23156 43708
rect 23436 42868 23492 44268
rect 24108 44322 24500 44324
rect 24108 44270 24110 44322
rect 24162 44270 24500 44322
rect 24108 44268 24500 44270
rect 24108 44258 24164 44268
rect 25676 44100 25732 44110
rect 25228 43650 25284 43662
rect 25228 43598 25230 43650
rect 25282 43598 25284 43650
rect 23548 42868 23604 42878
rect 23436 42866 23828 42868
rect 23436 42814 23550 42866
rect 23602 42814 23828 42866
rect 23436 42812 23828 42814
rect 23548 42802 23604 42812
rect 23772 42754 23828 42812
rect 23772 42702 23774 42754
rect 23826 42702 23828 42754
rect 23772 42690 23828 42702
rect 24556 42756 24612 42766
rect 24556 42662 24612 42700
rect 25228 42756 25284 43598
rect 25228 42690 25284 42700
rect 25452 43538 25508 43550
rect 25452 43486 25454 43538
rect 25506 43486 25508 43538
rect 25340 42196 25396 42206
rect 25452 42196 25508 43486
rect 25340 42194 25508 42196
rect 25340 42142 25342 42194
rect 25394 42142 25508 42194
rect 25340 42140 25508 42142
rect 25340 42130 25396 42140
rect 25564 42084 25620 42094
rect 24444 41076 24500 41086
rect 24444 40982 24500 41020
rect 25340 41076 25396 41086
rect 23100 40964 23156 40974
rect 23100 40740 23156 40908
rect 24108 40962 24164 40974
rect 24108 40910 24110 40962
rect 24162 40910 24164 40962
rect 23100 40684 23492 40740
rect 22988 40626 23380 40628
rect 22988 40574 22990 40626
rect 23042 40574 23380 40626
rect 22988 40572 23380 40574
rect 22988 40562 23044 40572
rect 22764 39554 22820 39564
rect 23324 39618 23380 40572
rect 23324 39566 23326 39618
rect 23378 39566 23380 39618
rect 23324 39554 23380 39566
rect 22876 39508 22932 39518
rect 22876 39506 23268 39508
rect 22876 39454 22878 39506
rect 22930 39454 23268 39506
rect 22876 39452 23268 39454
rect 22876 39442 22932 39452
rect 22652 38994 22708 39004
rect 23212 39058 23268 39452
rect 23212 39006 23214 39058
rect 23266 39006 23268 39058
rect 22988 38164 23044 38174
rect 22988 38070 23044 38108
rect 23212 38050 23268 39006
rect 23324 38724 23380 38734
rect 23324 38164 23380 38668
rect 23324 38098 23380 38108
rect 23212 37998 23214 38050
rect 23266 37998 23268 38050
rect 22316 37102 22318 37154
rect 22370 37102 22372 37154
rect 22316 37090 22372 37102
rect 22428 37100 22596 37156
rect 22764 37266 22820 37278
rect 22764 37214 22766 37266
rect 22818 37214 22820 37266
rect 22092 37042 22148 37054
rect 22092 36990 22094 37042
rect 22146 36990 22148 37042
rect 22092 36482 22148 36990
rect 22204 37044 22260 37054
rect 22204 36932 22260 36988
rect 22204 36876 22372 36932
rect 22092 36430 22094 36482
rect 22146 36430 22148 36482
rect 22092 36418 22148 36430
rect 22204 35812 22260 35822
rect 22204 35718 22260 35756
rect 21980 35700 22036 35710
rect 21868 35698 22036 35700
rect 21868 35646 21982 35698
rect 22034 35646 22036 35698
rect 21868 35644 22036 35646
rect 21980 35028 22036 35644
rect 22316 35588 22372 36876
rect 22428 35812 22484 37100
rect 22540 36484 22596 36494
rect 22540 36390 22596 36428
rect 22652 36258 22708 36270
rect 22652 36206 22654 36258
rect 22706 36206 22708 36258
rect 22540 35812 22596 35822
rect 22428 35810 22596 35812
rect 22428 35758 22542 35810
rect 22594 35758 22596 35810
rect 22428 35756 22596 35758
rect 22540 35746 22596 35756
rect 21980 34962 22036 34972
rect 22204 35532 22372 35588
rect 21980 34690 22036 34702
rect 21980 34638 21982 34690
rect 22034 34638 22036 34690
rect 21980 34130 22036 34638
rect 21980 34078 21982 34130
rect 22034 34078 22036 34130
rect 21980 34066 22036 34078
rect 21756 32498 21812 32508
rect 22092 32676 22148 32686
rect 21532 29484 21644 29540
rect 20748 28700 21028 28756
rect 20748 28532 20804 28542
rect 20748 28438 20804 28476
rect 20524 28364 20636 28420
rect 20636 28354 20692 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 27806 19630 27858
rect 19682 27806 19684 27858
rect 19628 27794 19684 27806
rect 19628 27188 19684 27198
rect 20636 27188 20692 27198
rect 20860 27188 20916 27198
rect 19628 27074 19684 27132
rect 20300 27186 20860 27188
rect 20300 27134 20638 27186
rect 20690 27134 20860 27186
rect 20300 27132 20860 27134
rect 19628 27022 19630 27074
rect 19682 27022 19684 27074
rect 19628 27010 19684 27022
rect 19740 27076 19796 27086
rect 19740 26982 19796 27020
rect 20300 27074 20356 27132
rect 20636 27122 20692 27132
rect 20860 27122 20916 27132
rect 20300 27022 20302 27074
rect 20354 27022 20356 27074
rect 20300 27010 20356 27022
rect 19852 26852 19908 26862
rect 19516 26238 19518 26290
rect 19570 26238 19572 26290
rect 19516 26226 19572 26238
rect 19628 26850 19908 26852
rect 19628 26798 19854 26850
rect 19906 26798 19908 26850
rect 19628 26796 19908 26798
rect 19628 26292 19684 26796
rect 19852 26786 19908 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20188 26628 20244 26638
rect 19852 26516 19908 26526
rect 19852 26514 20132 26516
rect 19852 26462 19854 26514
rect 19906 26462 20132 26514
rect 19852 26460 20132 26462
rect 19852 26450 19908 26460
rect 19852 26292 19908 26302
rect 19628 26290 19908 26292
rect 19628 26238 19854 26290
rect 19906 26238 19908 26290
rect 19628 26236 19908 26238
rect 19068 25564 19460 25620
rect 19740 25620 19796 25630
rect 19068 25282 19124 25564
rect 19740 25506 19796 25564
rect 19740 25454 19742 25506
rect 19794 25454 19796 25506
rect 19740 25442 19796 25454
rect 19292 25396 19348 25406
rect 19292 25302 19348 25340
rect 19068 25230 19070 25282
rect 19122 25230 19124 25282
rect 19068 24948 19124 25230
rect 19180 25284 19236 25294
rect 19180 25190 19236 25228
rect 19852 25284 19908 26236
rect 19964 25508 20020 25518
rect 19964 25394 20020 25452
rect 19964 25342 19966 25394
rect 20018 25342 20020 25394
rect 19964 25330 20020 25342
rect 20076 25284 20132 26460
rect 20188 26402 20244 26572
rect 20748 26628 20804 26638
rect 20748 26514 20804 26572
rect 20748 26462 20750 26514
rect 20802 26462 20804 26514
rect 20748 26450 20804 26462
rect 20188 26350 20190 26402
rect 20242 26350 20244 26402
rect 20188 26338 20244 26350
rect 20300 25620 20356 25630
rect 20300 25284 20356 25564
rect 20412 25284 20468 25294
rect 20076 25228 20244 25284
rect 19852 25218 19908 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19068 24882 19124 24892
rect 20188 24276 20244 25228
rect 20300 25282 20468 25284
rect 20300 25230 20414 25282
rect 20466 25230 20468 25282
rect 20300 25228 20468 25230
rect 20300 24500 20356 25228
rect 20412 25218 20468 25228
rect 20748 24948 20804 24958
rect 20748 24854 20804 24892
rect 20412 24724 20468 24734
rect 20860 24724 20916 24734
rect 20412 24722 20916 24724
rect 20412 24670 20414 24722
rect 20466 24670 20862 24722
rect 20914 24670 20916 24722
rect 20412 24668 20916 24670
rect 20412 24658 20468 24668
rect 20860 24658 20916 24668
rect 20972 24500 21028 28700
rect 21308 27074 21364 27086
rect 21308 27022 21310 27074
rect 21362 27022 21364 27074
rect 21308 26964 21364 27022
rect 21532 27076 21588 29484
rect 21644 29474 21700 29484
rect 21756 31780 21812 31790
rect 21756 29876 21812 31724
rect 21868 31778 21924 31790
rect 21868 31726 21870 31778
rect 21922 31726 21924 31778
rect 21868 31668 21924 31726
rect 21868 31602 21924 31612
rect 22092 30434 22148 32620
rect 22092 30382 22094 30434
rect 22146 30382 22148 30434
rect 22092 30370 22148 30382
rect 21756 29426 21812 29820
rect 21756 29374 21758 29426
rect 21810 29374 21812 29426
rect 21644 28532 21700 28542
rect 21644 27298 21700 28476
rect 21644 27246 21646 27298
rect 21698 27246 21700 27298
rect 21644 27234 21700 27246
rect 21756 27188 21812 29374
rect 22092 29314 22148 29326
rect 22092 29262 22094 29314
rect 22146 29262 22148 29314
rect 21980 28420 22036 28430
rect 21980 28082 22036 28364
rect 21980 28030 21982 28082
rect 22034 28030 22036 28082
rect 21980 28018 22036 28030
rect 22092 27300 22148 29262
rect 22092 27234 22148 27244
rect 21756 27122 21812 27132
rect 21532 27020 21700 27076
rect 21308 26898 21364 26908
rect 21644 26908 21700 27020
rect 21532 26852 21588 26862
rect 21644 26852 21812 26908
rect 21532 26758 21588 26796
rect 21756 26740 21812 26852
rect 21756 26674 21812 26684
rect 22204 26516 22260 35532
rect 22652 35140 22708 36206
rect 22764 35924 22820 37214
rect 23100 37266 23156 37278
rect 23100 37214 23102 37266
rect 23154 37214 23156 37266
rect 23100 37044 23156 37214
rect 23100 36978 23156 36988
rect 22764 35858 22820 35868
rect 23100 36370 23156 36382
rect 23100 36318 23102 36370
rect 23154 36318 23156 36370
rect 23100 35922 23156 36318
rect 23100 35870 23102 35922
rect 23154 35870 23156 35922
rect 23100 35858 23156 35870
rect 22988 35810 23044 35822
rect 22988 35758 22990 35810
rect 23042 35758 23044 35810
rect 22764 35700 22820 35710
rect 22988 35700 23044 35758
rect 23100 35700 23156 35710
rect 22988 35644 23100 35700
rect 22764 35606 22820 35644
rect 22652 35074 22708 35084
rect 22764 35028 22820 35038
rect 23100 35028 23156 35644
rect 22820 34972 22932 35028
rect 22764 34962 22820 34972
rect 22876 34914 22932 34972
rect 22876 34862 22878 34914
rect 22930 34862 22932 34914
rect 22876 34850 22932 34862
rect 22988 34972 23156 35028
rect 22316 34804 22372 34814
rect 22988 34804 23044 34972
rect 23212 34916 23268 37998
rect 23324 36484 23380 36494
rect 23324 36390 23380 36428
rect 23436 35588 23492 40684
rect 23548 40404 23604 40414
rect 23548 40310 23604 40348
rect 24108 39618 24164 40910
rect 24556 40852 24612 40862
rect 24108 39566 24110 39618
rect 24162 39566 24164 39618
rect 24108 39554 24164 39566
rect 24220 40290 24276 40302
rect 24220 40238 24222 40290
rect 24274 40238 24276 40290
rect 23772 38722 23828 38734
rect 23772 38670 23774 38722
rect 23826 38670 23828 38722
rect 23772 38164 23828 38670
rect 24108 38724 24164 38762
rect 24108 38658 24164 38668
rect 24220 38612 24276 40238
rect 24332 39396 24388 39406
rect 24332 38836 24388 39340
rect 24332 38742 24388 38780
rect 23772 38098 23828 38108
rect 24108 38388 24164 38398
rect 24108 38162 24164 38332
rect 24108 38110 24110 38162
rect 24162 38110 24164 38162
rect 24108 38098 24164 38110
rect 24220 38052 24276 38556
rect 24220 37986 24276 37996
rect 24556 37938 24612 40796
rect 25340 40626 25396 41020
rect 25340 40574 25342 40626
rect 25394 40574 25396 40626
rect 25340 40562 25396 40574
rect 24668 40290 24724 40302
rect 24668 40238 24670 40290
rect 24722 40238 24724 40290
rect 24668 38836 24724 40238
rect 25116 40292 25172 40302
rect 24668 38770 24724 38780
rect 24780 39620 24836 39630
rect 24780 38668 24836 39564
rect 24668 38610 24724 38622
rect 24780 38612 24948 38668
rect 24668 38558 24670 38610
rect 24722 38558 24724 38610
rect 24668 38276 24724 38558
rect 24668 38220 24836 38276
rect 24780 38052 24836 38220
rect 24780 37986 24836 37996
rect 24556 37886 24558 37938
rect 24610 37886 24612 37938
rect 24556 37874 24612 37886
rect 24668 37940 24724 37950
rect 24668 37846 24724 37884
rect 23548 37828 23604 37838
rect 24332 37828 24388 37838
rect 23548 37826 24052 37828
rect 23548 37774 23550 37826
rect 23602 37774 24052 37826
rect 23548 37772 24052 37774
rect 23548 37762 23604 37772
rect 23884 37266 23940 37278
rect 23884 37214 23886 37266
rect 23938 37214 23940 37266
rect 23772 37156 23828 37166
rect 23548 37154 23828 37156
rect 23548 37102 23774 37154
rect 23826 37102 23828 37154
rect 23548 37100 23828 37102
rect 23548 36482 23604 37100
rect 23772 37090 23828 37100
rect 23548 36430 23550 36482
rect 23602 36430 23604 36482
rect 23548 36418 23604 36430
rect 23884 37044 23940 37214
rect 23996 37268 24052 37772
rect 24220 37826 24388 37828
rect 24220 37774 24334 37826
rect 24386 37774 24388 37826
rect 24220 37772 24388 37774
rect 24108 37268 24164 37278
rect 23996 37266 24164 37268
rect 23996 37214 24110 37266
rect 24162 37214 24164 37266
rect 23996 37212 24164 37214
rect 24220 37268 24276 37772
rect 24332 37762 24388 37772
rect 24444 37828 24500 37838
rect 24332 37492 24388 37502
rect 24444 37492 24500 37772
rect 24892 37716 24948 38612
rect 24332 37490 24500 37492
rect 24332 37438 24334 37490
rect 24386 37438 24500 37490
rect 24332 37436 24500 37438
rect 24556 37660 24948 37716
rect 25004 38164 25060 38174
rect 24556 37490 24612 37660
rect 24556 37438 24558 37490
rect 24610 37438 24612 37490
rect 24332 37426 24388 37436
rect 24556 37426 24612 37438
rect 24220 37212 24388 37268
rect 24108 37202 24164 37212
rect 23884 36484 23940 36988
rect 24332 36484 24388 37212
rect 25004 37044 25060 38108
rect 25004 36978 25060 36988
rect 24780 36932 24836 36942
rect 24780 36596 24836 36876
rect 24892 36708 24948 36718
rect 24892 36614 24948 36652
rect 24780 36530 24836 36540
rect 23884 36428 24052 36484
rect 23772 36370 23828 36382
rect 23772 36318 23774 36370
rect 23826 36318 23828 36370
rect 23772 36260 23828 36318
rect 23772 36194 23828 36204
rect 23884 36258 23940 36270
rect 23884 36206 23886 36258
rect 23938 36206 23940 36258
rect 23660 35924 23716 35934
rect 23660 35698 23716 35868
rect 23660 35646 23662 35698
rect 23714 35646 23716 35698
rect 23660 35634 23716 35646
rect 23436 35522 23492 35532
rect 23548 35586 23604 35598
rect 23548 35534 23550 35586
rect 23602 35534 23604 35586
rect 23324 35476 23380 35486
rect 23324 35382 23380 35420
rect 23548 35252 23604 35534
rect 23548 35186 23604 35196
rect 22316 34802 22596 34804
rect 22316 34750 22318 34802
rect 22370 34750 22596 34802
rect 22316 34748 22596 34750
rect 22316 34738 22372 34748
rect 22540 33570 22596 34748
rect 22988 34738 23044 34748
rect 23100 34860 23268 34916
rect 23884 34916 23940 36206
rect 23996 35812 24052 36428
rect 24332 36418 24388 36428
rect 24444 36428 24724 36484
rect 24220 36260 24276 36270
rect 24444 36260 24500 36428
rect 24668 36372 24724 36428
rect 25116 36482 25172 40236
rect 25564 40180 25620 42028
rect 25676 41746 25732 44044
rect 25676 41694 25678 41746
rect 25730 41694 25732 41746
rect 25676 40404 25732 41694
rect 25788 41636 25844 44828
rect 25788 41580 25956 41636
rect 25676 40338 25732 40348
rect 25676 40180 25732 40190
rect 25564 40178 25732 40180
rect 25564 40126 25678 40178
rect 25730 40126 25732 40178
rect 25564 40124 25732 40126
rect 25452 38724 25508 38762
rect 25452 38658 25508 38668
rect 25228 38500 25284 38510
rect 25228 37604 25284 38444
rect 25340 38388 25396 38398
rect 25340 38050 25396 38332
rect 25564 38276 25620 40124
rect 25676 40114 25732 40124
rect 25788 38724 25844 38762
rect 25788 38658 25844 38668
rect 25900 38668 25956 41580
rect 26012 38834 26068 45612
rect 26124 45106 26180 46622
rect 26124 45054 26126 45106
rect 26178 45054 26180 45106
rect 26124 41970 26180 45054
rect 26236 45218 26292 45230
rect 26236 45166 26238 45218
rect 26290 45166 26292 45218
rect 26236 44100 26292 45166
rect 26348 44884 26404 46734
rect 26908 46116 26964 48076
rect 27692 48020 27748 48030
rect 27692 47124 27748 47964
rect 27692 47068 28084 47124
rect 27804 46788 27860 46798
rect 27580 46786 27860 46788
rect 27580 46734 27806 46786
rect 27858 46734 27860 46786
rect 27580 46732 27860 46734
rect 27468 46676 27524 46686
rect 26908 46002 26964 46060
rect 27356 46674 27524 46676
rect 27356 46622 27470 46674
rect 27522 46622 27524 46674
rect 27356 46620 27524 46622
rect 27356 46114 27412 46620
rect 27468 46610 27524 46620
rect 27356 46062 27358 46114
rect 27410 46062 27412 46114
rect 27356 46050 27412 46062
rect 26908 45950 26910 46002
rect 26962 45950 26964 46002
rect 26908 45938 26964 45950
rect 27020 45108 27076 45118
rect 27020 45014 27076 45052
rect 27580 45106 27636 46732
rect 27804 46722 27860 46732
rect 27692 46116 27748 46126
rect 27692 46022 27748 46060
rect 27580 45054 27582 45106
rect 27634 45054 27636 45106
rect 27580 45042 27636 45054
rect 26348 44818 26404 44828
rect 27916 44996 27972 45006
rect 27916 44210 27972 44940
rect 27916 44158 27918 44210
rect 27970 44158 27972 44210
rect 27916 44146 27972 44158
rect 26460 44100 26516 44110
rect 26292 44098 26516 44100
rect 26292 44046 26462 44098
rect 26514 44046 26516 44098
rect 26292 44044 26516 44046
rect 26236 44034 26292 44044
rect 26460 44034 26516 44044
rect 27356 44100 27412 44110
rect 27580 44100 27636 44110
rect 27356 44098 27636 44100
rect 27356 44046 27358 44098
rect 27410 44046 27582 44098
rect 27634 44046 27636 44098
rect 27356 44044 27636 44046
rect 27356 44034 27412 44044
rect 26908 42530 26964 42542
rect 26908 42478 26910 42530
rect 26962 42478 26964 42530
rect 26236 42084 26292 42094
rect 26236 41990 26292 42028
rect 26908 42084 26964 42478
rect 26908 42018 26964 42028
rect 26124 41918 26126 41970
rect 26178 41918 26180 41970
rect 26124 41860 26180 41918
rect 26124 41804 26740 41860
rect 26348 40402 26404 41804
rect 26684 41298 26740 41804
rect 27580 41412 27636 44044
rect 28028 43708 28084 47068
rect 28476 47012 28532 48190
rect 28700 47460 28756 48972
rect 29260 48934 29316 48972
rect 29708 48962 29764 48972
rect 29820 48468 29876 49758
rect 32620 49812 32676 49822
rect 32620 49810 32788 49812
rect 32620 49758 32622 49810
rect 32674 49758 32788 49810
rect 32620 49756 32788 49758
rect 32620 49746 32676 49756
rect 32396 49028 32452 49038
rect 32620 49028 32676 49038
rect 32452 49026 32676 49028
rect 32452 48974 32622 49026
rect 32674 48974 32676 49026
rect 32452 48972 32676 48974
rect 32172 48802 32228 48814
rect 32172 48750 32174 48802
rect 32226 48750 32228 48802
rect 29932 48468 29988 48478
rect 29820 48466 29988 48468
rect 29820 48414 29934 48466
rect 29986 48414 29988 48466
rect 29820 48412 29988 48414
rect 29932 48402 29988 48412
rect 30828 48356 30884 48366
rect 30268 48244 30324 48254
rect 30268 48150 30324 48188
rect 30716 48242 30772 48254
rect 30716 48190 30718 48242
rect 30770 48190 30772 48242
rect 30716 48132 30772 48190
rect 28700 47404 29428 47460
rect 28476 46946 28532 46956
rect 28364 45890 28420 45902
rect 28364 45838 28366 45890
rect 28418 45838 28420 45890
rect 28364 44884 28420 45838
rect 28476 45778 28532 45790
rect 28476 45726 28478 45778
rect 28530 45726 28532 45778
rect 28476 45332 28532 45726
rect 28476 45266 28532 45276
rect 29036 45332 29092 45342
rect 28364 44818 28420 44828
rect 28028 43652 28196 43708
rect 28028 43540 28084 43550
rect 28028 43446 28084 43484
rect 27804 41970 27860 41982
rect 27804 41918 27806 41970
rect 27858 41918 27860 41970
rect 26684 41246 26686 41298
rect 26738 41246 26740 41298
rect 26684 41234 26740 41246
rect 27132 41356 27748 41412
rect 26460 40516 26516 40526
rect 26460 40514 26628 40516
rect 26460 40462 26462 40514
rect 26514 40462 26628 40514
rect 26460 40460 26628 40462
rect 26460 40450 26516 40460
rect 26348 40350 26350 40402
rect 26402 40350 26404 40402
rect 26348 40338 26404 40350
rect 26460 39396 26516 39406
rect 26572 39396 26628 40460
rect 27132 39396 27188 41356
rect 27692 41298 27748 41356
rect 27692 41246 27694 41298
rect 27746 41246 27748 41298
rect 27692 41234 27748 41246
rect 27356 41188 27412 41198
rect 26516 39340 26628 39396
rect 26908 39394 27188 39396
rect 26908 39342 27134 39394
rect 27186 39342 27188 39394
rect 26908 39340 27188 39342
rect 26460 39302 26516 39340
rect 26012 38782 26014 38834
rect 26066 38782 26068 38834
rect 26012 38770 26068 38782
rect 26236 38892 26628 38948
rect 26236 38668 26292 38892
rect 25900 38612 26292 38668
rect 26348 38610 26404 38622
rect 26348 38558 26350 38610
rect 26402 38558 26404 38610
rect 25564 38220 26180 38276
rect 25340 37998 25342 38050
rect 25394 37998 25396 38050
rect 25340 37986 25396 37998
rect 25676 38052 25732 38062
rect 25676 37958 25732 37996
rect 25900 37828 25956 37838
rect 25900 37734 25956 37772
rect 26012 37826 26068 37838
rect 26012 37774 26014 37826
rect 26066 37774 26068 37826
rect 25788 37716 25844 37726
rect 25228 37538 25284 37548
rect 25564 37660 25788 37716
rect 25564 37490 25620 37660
rect 25788 37650 25844 37660
rect 25564 37438 25566 37490
rect 25618 37438 25620 37490
rect 25564 37426 25620 37438
rect 25788 37492 25844 37502
rect 26012 37492 26068 37774
rect 26124 37826 26180 38220
rect 26348 38052 26404 38558
rect 26348 37986 26404 37996
rect 26572 37938 26628 38892
rect 26796 38722 26852 38734
rect 26796 38670 26798 38722
rect 26850 38670 26852 38722
rect 26796 38668 26852 38670
rect 26572 37886 26574 37938
rect 26626 37886 26628 37938
rect 26572 37874 26628 37886
rect 26684 38612 26852 38668
rect 26684 38276 26740 38612
rect 26684 38050 26740 38220
rect 26684 37998 26686 38050
rect 26738 37998 26740 38050
rect 26124 37774 26126 37826
rect 26178 37774 26180 37826
rect 26124 37762 26180 37774
rect 26348 37826 26404 37838
rect 26348 37774 26350 37826
rect 26402 37774 26404 37826
rect 26348 37716 26404 37774
rect 26348 37650 26404 37660
rect 25788 37490 26068 37492
rect 25788 37438 25790 37490
rect 25842 37438 26068 37490
rect 25788 37436 26068 37438
rect 26124 37604 26180 37614
rect 25788 37426 25844 37436
rect 26124 37380 26180 37548
rect 26460 37604 26516 37614
rect 26460 37490 26516 37548
rect 26460 37438 26462 37490
rect 26514 37438 26516 37490
rect 26460 37426 26516 37438
rect 26012 37324 26180 37380
rect 25340 37266 25396 37278
rect 25340 37214 25342 37266
rect 25394 37214 25396 37266
rect 25340 36708 25396 37214
rect 26012 37266 26068 37324
rect 26012 37214 26014 37266
rect 26066 37214 26068 37266
rect 26012 37202 26068 37214
rect 26124 37154 26180 37166
rect 26124 37102 26126 37154
rect 26178 37102 26180 37154
rect 25340 36642 25396 36652
rect 26012 36932 26068 36942
rect 25116 36430 25118 36482
rect 25170 36430 25172 36482
rect 25116 36418 25172 36430
rect 26012 36482 26068 36876
rect 26012 36430 26014 36482
rect 26066 36430 26068 36482
rect 26012 36418 26068 36430
rect 26124 36484 26180 37102
rect 26236 36484 26292 36494
rect 26124 36482 26292 36484
rect 26124 36430 26238 36482
rect 26290 36430 26292 36482
rect 26124 36428 26292 36430
rect 26236 36418 26292 36428
rect 26460 36484 26516 36494
rect 24780 36372 24836 36382
rect 24668 36370 24836 36372
rect 24668 36318 24782 36370
rect 24834 36318 24836 36370
rect 24668 36316 24836 36318
rect 24780 36306 24836 36316
rect 24220 36258 24500 36260
rect 24220 36206 24222 36258
rect 24274 36206 24500 36258
rect 24220 36204 24500 36206
rect 24556 36258 24612 36270
rect 24556 36206 24558 36258
rect 24610 36206 24612 36258
rect 24108 35812 24164 35822
rect 23996 35756 24108 35812
rect 24108 35718 24164 35756
rect 22540 33518 22542 33570
rect 22594 33518 22596 33570
rect 22540 33506 22596 33518
rect 22876 33348 22932 33358
rect 22652 33346 22932 33348
rect 22652 33294 22878 33346
rect 22930 33294 22932 33346
rect 22652 33292 22932 33294
rect 22652 31892 22708 33292
rect 22876 33282 22932 33292
rect 22540 31780 22596 31790
rect 22540 31686 22596 31724
rect 22652 31668 22708 31836
rect 22652 31666 22820 31668
rect 22652 31614 22654 31666
rect 22706 31614 22820 31666
rect 22652 31612 22820 31614
rect 22652 31602 22708 31612
rect 22764 31218 22820 31612
rect 22764 31166 22766 31218
rect 22818 31166 22820 31218
rect 22764 31154 22820 31166
rect 23100 30996 23156 34860
rect 23884 34850 23940 34860
rect 23212 34690 23268 34702
rect 23212 34638 23214 34690
rect 23266 34638 23268 34690
rect 23212 34468 23268 34638
rect 23212 34402 23268 34412
rect 24108 33348 24164 33358
rect 24108 33254 24164 33292
rect 23212 33234 23268 33246
rect 23212 33182 23214 33234
rect 23266 33182 23268 33234
rect 23212 31780 23268 33182
rect 23660 33234 23716 33246
rect 23660 33182 23662 33234
rect 23714 33182 23716 33234
rect 23660 32228 23716 33182
rect 24220 32900 24276 36204
rect 24556 35700 24612 36206
rect 24556 35634 24612 35644
rect 25452 36258 25508 36270
rect 26348 36260 26404 36270
rect 25452 36206 25454 36258
rect 25506 36206 25508 36258
rect 25452 35812 25508 36206
rect 24892 35364 24948 35374
rect 24556 34692 24612 34702
rect 24556 34598 24612 34636
rect 24444 34018 24500 34030
rect 24444 33966 24446 34018
rect 24498 33966 24500 34018
rect 24332 33460 24388 33470
rect 24332 33366 24388 33404
rect 24108 32844 24276 32900
rect 23660 32172 24052 32228
rect 23660 31892 23716 31902
rect 23660 31798 23716 31836
rect 23212 31714 23268 31724
rect 23884 31666 23940 31678
rect 23884 31614 23886 31666
rect 23938 31614 23940 31666
rect 23324 31556 23380 31566
rect 23884 31556 23940 31614
rect 23324 31554 23828 31556
rect 23324 31502 23326 31554
rect 23378 31502 23828 31554
rect 23324 31500 23828 31502
rect 23324 31490 23380 31500
rect 23772 31108 23828 31500
rect 23884 31490 23940 31500
rect 23884 31108 23940 31118
rect 23772 31106 23940 31108
rect 23772 31054 23886 31106
rect 23938 31054 23940 31106
rect 23772 31052 23940 31054
rect 23884 31042 23940 31052
rect 22204 26450 22260 26460
rect 22316 30940 23156 30996
rect 21644 26290 21700 26302
rect 21644 26238 21646 26290
rect 21698 26238 21700 26290
rect 21308 25396 21364 25406
rect 21308 25302 21364 25340
rect 20300 24444 20468 24500
rect 20188 24220 20356 24276
rect 20188 23940 20244 23950
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23380 20244 23884
rect 19740 23156 19796 23166
rect 18956 23090 19012 23100
rect 19628 23100 19740 23156
rect 17724 21812 17780 21822
rect 17724 21586 17780 21756
rect 18172 21698 18228 22204
rect 18172 21646 18174 21698
rect 18226 21646 18228 21698
rect 18172 21634 18228 21646
rect 18284 22372 18340 22382
rect 17724 21534 17726 21586
rect 17778 21534 17780 21586
rect 17724 21522 17780 21534
rect 18284 21252 18340 22316
rect 19516 22260 19572 22270
rect 18284 21186 18340 21196
rect 18396 22148 18452 22158
rect 18172 20916 18228 20926
rect 18060 20802 18116 20814
rect 18060 20750 18062 20802
rect 18114 20750 18116 20802
rect 18060 20244 18116 20750
rect 17612 19908 17668 19918
rect 17612 19906 17780 19908
rect 17612 19854 17614 19906
rect 17666 19854 17780 19906
rect 17612 19852 17780 19854
rect 17612 19842 17668 19852
rect 17164 19516 17332 19572
rect 16828 19282 16884 19292
rect 17052 19460 17108 19470
rect 17052 18452 17108 19404
rect 17052 18386 17108 18396
rect 16100 17836 16324 17892
rect 16604 18004 16660 18014
rect 16044 17798 16100 17836
rect 16604 17780 16660 17948
rect 16604 17714 16660 17724
rect 16716 17892 16772 17902
rect 15820 17666 15876 17678
rect 15820 17614 15822 17666
rect 15874 17614 15876 17666
rect 15484 17444 15540 17454
rect 15372 17108 15428 17118
rect 15372 17014 15428 17052
rect 15484 16994 15540 17388
rect 15484 16942 15486 16994
rect 15538 16942 15540 16994
rect 15484 16930 15540 16942
rect 15820 16996 15876 17614
rect 16156 17668 16212 17678
rect 16716 17668 16772 17836
rect 17052 17780 17108 17790
rect 16716 17612 16884 17668
rect 16156 17574 16212 17612
rect 16156 17444 16212 17454
rect 16156 17350 16212 17388
rect 16716 17442 16772 17454
rect 16716 17390 16718 17442
rect 16770 17390 16772 17442
rect 16044 16996 16100 17006
rect 15820 16940 16044 16996
rect 16044 16902 16100 16940
rect 16492 16996 16548 17006
rect 16716 16996 16772 17390
rect 16492 16994 16660 16996
rect 16492 16942 16494 16994
rect 16546 16942 16660 16994
rect 16492 16940 16660 16942
rect 16492 16930 16548 16940
rect 16604 16884 16660 16940
rect 16716 16930 16772 16940
rect 16828 16994 16884 17612
rect 17052 17666 17108 17724
rect 17052 17614 17054 17666
rect 17106 17614 17108 17666
rect 17052 17602 17108 17614
rect 16828 16942 16830 16994
rect 16882 16942 16884 16994
rect 16828 16930 16884 16942
rect 15372 16660 15428 16670
rect 15372 16658 15652 16660
rect 15372 16606 15374 16658
rect 15426 16606 15652 16658
rect 15372 16604 15652 16606
rect 15372 16594 15428 16604
rect 15260 16380 15540 16436
rect 14700 16098 14868 16100
rect 14700 16046 14702 16098
rect 14754 16046 14868 16098
rect 14700 16044 14868 16046
rect 15372 16100 15428 16110
rect 14476 15596 14644 15652
rect 14364 15250 14420 15260
rect 14476 15202 14532 15214
rect 14476 15150 14478 15202
rect 14530 15150 14532 15202
rect 14476 15148 14532 15150
rect 14252 15092 14532 15148
rect 13132 15026 13188 15036
rect 12908 14420 12964 14430
rect 12908 14418 13412 14420
rect 12908 14366 12910 14418
rect 12962 14366 13412 14418
rect 12908 14364 13412 14366
rect 12908 14354 12964 14364
rect 13356 13076 13412 14364
rect 14364 14308 14420 14318
rect 14364 14214 14420 14252
rect 14588 13860 14644 15596
rect 14028 13804 14644 13860
rect 14700 14644 14756 16044
rect 15372 15986 15428 16044
rect 15372 15934 15374 15986
rect 15426 15934 15428 15986
rect 14924 15876 14980 15886
rect 14924 15874 15092 15876
rect 14924 15822 14926 15874
rect 14978 15822 15092 15874
rect 14924 15820 15092 15822
rect 14924 15810 14980 15820
rect 14924 15316 14980 15326
rect 15036 15316 15092 15820
rect 15260 15540 15316 15550
rect 15260 15316 15316 15484
rect 15036 15260 15316 15316
rect 15372 15314 15428 15934
rect 15372 15262 15374 15314
rect 15426 15262 15428 15314
rect 14924 15222 14980 15260
rect 15372 15250 15428 15262
rect 15484 15148 15540 16380
rect 15596 15764 15652 16604
rect 15820 16658 15876 16670
rect 15820 16606 15822 16658
rect 15874 16606 15876 16658
rect 15820 16098 15876 16606
rect 16156 16660 16212 16670
rect 16156 16566 16212 16604
rect 16268 16212 16324 16222
rect 16268 16100 16324 16156
rect 15820 16046 15822 16098
rect 15874 16046 15876 16098
rect 15820 15764 15876 16046
rect 15596 15708 15764 15764
rect 15596 15540 15652 15550
rect 15596 15314 15652 15484
rect 15596 15262 15598 15314
rect 15650 15262 15652 15314
rect 15596 15250 15652 15262
rect 15708 15148 15764 15708
rect 15820 15698 15876 15708
rect 15932 16098 16324 16100
rect 15932 16046 16270 16098
rect 16322 16046 16324 16098
rect 15932 16044 16324 16046
rect 15820 15316 15876 15326
rect 15932 15316 15988 16044
rect 16268 16034 16324 16044
rect 16268 15874 16324 15886
rect 16268 15822 16270 15874
rect 16322 15822 16324 15874
rect 15820 15314 15988 15316
rect 15820 15262 15822 15314
rect 15874 15262 15988 15314
rect 15820 15260 15988 15262
rect 16044 15314 16100 15326
rect 16044 15262 16046 15314
rect 16098 15262 16100 15314
rect 15820 15250 15876 15260
rect 15260 15092 15316 15102
rect 13468 13076 13524 13086
rect 12796 13074 13188 13076
rect 12796 13022 12798 13074
rect 12850 13022 13188 13074
rect 12796 13020 13188 13022
rect 13356 13074 13524 13076
rect 13356 13022 13470 13074
rect 13522 13022 13524 13074
rect 13356 13020 13524 13022
rect 12796 13010 12852 13020
rect 12908 11508 12964 13020
rect 13132 12402 13188 13020
rect 13468 13010 13524 13020
rect 14028 12964 14084 13804
rect 14140 13636 14196 13646
rect 14700 13636 14756 14588
rect 15148 15090 15316 15092
rect 15148 15038 15262 15090
rect 15314 15038 15316 15090
rect 15148 15036 15316 15038
rect 14140 13634 14756 13636
rect 14140 13582 14142 13634
rect 14194 13582 14756 13634
rect 14140 13580 14756 13582
rect 15036 13636 15092 13646
rect 14140 13570 14196 13580
rect 15036 13542 15092 13580
rect 14252 13300 14308 13310
rect 14140 12964 14196 12974
rect 14028 12962 14196 12964
rect 14028 12910 14142 12962
rect 14194 12910 14196 12962
rect 14028 12908 14196 12910
rect 14140 12740 14196 12908
rect 14140 12674 14196 12684
rect 13132 12350 13134 12402
rect 13186 12350 13188 12402
rect 13132 12338 13188 12350
rect 14140 11844 14196 11854
rect 14252 11844 14308 13244
rect 15148 13188 15204 15036
rect 15260 15026 15316 15036
rect 15372 15092 15540 15148
rect 15596 15092 15764 15148
rect 16044 15204 16100 15262
rect 16268 15148 16324 15822
rect 16492 15540 16548 15550
rect 16492 15426 16548 15484
rect 16492 15374 16494 15426
rect 16546 15374 16548 15426
rect 16492 15362 16548 15374
rect 16044 15138 16100 15148
rect 16156 15092 16324 15148
rect 16604 15148 16660 16828
rect 16716 16436 16772 16446
rect 16716 15988 16772 16380
rect 16828 15988 16884 15998
rect 16716 15986 16884 15988
rect 16716 15934 16830 15986
rect 16882 15934 16884 15986
rect 16716 15932 16884 15934
rect 16828 15922 16884 15932
rect 15260 13860 15316 13870
rect 15260 13766 15316 13804
rect 14924 13132 15204 13188
rect 15260 13524 15316 13534
rect 14364 13076 14420 13086
rect 14364 12982 14420 13020
rect 14812 13076 14868 13086
rect 14812 12982 14868 13020
rect 14588 12292 14644 12302
rect 14588 12290 14868 12292
rect 14588 12238 14590 12290
rect 14642 12238 14868 12290
rect 14588 12236 14868 12238
rect 14588 12226 14644 12236
rect 14364 12178 14420 12190
rect 14364 12126 14366 12178
rect 14418 12126 14420 12178
rect 14364 11956 14420 12126
rect 14364 11890 14420 11900
rect 14476 12066 14532 12078
rect 14476 12014 14478 12066
rect 14530 12014 14532 12066
rect 14196 11788 14308 11844
rect 14140 11778 14196 11788
rect 14476 11620 14532 12014
rect 14700 12068 14756 12078
rect 14700 11732 14756 12012
rect 14028 11564 14532 11620
rect 14588 11676 14756 11732
rect 12908 11394 12964 11452
rect 13916 11508 13972 11518
rect 13916 11414 13972 11452
rect 12908 11342 12910 11394
rect 12962 11342 12964 11394
rect 12908 11330 12964 11342
rect 14028 10948 14084 11564
rect 14252 11396 14308 11406
rect 14252 11302 14308 11340
rect 14476 11396 14532 11406
rect 14588 11396 14644 11676
rect 14476 11394 14644 11396
rect 14476 11342 14478 11394
rect 14530 11342 14644 11394
rect 14476 11340 14644 11342
rect 14700 11508 14756 11518
rect 13916 10892 14084 10948
rect 13916 10610 13972 10892
rect 14140 10836 14196 10846
rect 13916 10558 13918 10610
rect 13970 10558 13972 10610
rect 13916 10546 13972 10558
rect 14028 10722 14084 10734
rect 14028 10670 14030 10722
rect 14082 10670 14084 10722
rect 13132 10500 13188 10510
rect 13188 10444 13300 10500
rect 13132 10434 13188 10444
rect 12908 10388 12964 10398
rect 12908 10294 12964 10332
rect 13244 10386 13300 10444
rect 13244 10334 13246 10386
rect 13298 10334 13300 10386
rect 13244 10322 13300 10334
rect 13580 10388 13636 10398
rect 13132 10276 13188 10286
rect 12684 10108 12852 10164
rect 12572 10050 12628 10062
rect 12572 9998 12574 10050
rect 12626 9998 12628 10050
rect 12572 9828 12628 9998
rect 12684 9940 12740 9950
rect 12684 9846 12740 9884
rect 12572 9042 12628 9772
rect 12572 8990 12574 9042
rect 12626 8990 12628 9042
rect 12572 8978 12628 8990
rect 12460 8878 12462 8930
rect 12514 8878 12516 8930
rect 12460 8866 12516 8878
rect 12236 8082 12292 8092
rect 12572 8148 12628 8158
rect 12572 8054 12628 8092
rect 12796 8146 12852 10108
rect 12796 8094 12798 8146
rect 12850 8094 12852 8146
rect 12684 8034 12740 8046
rect 12684 7982 12686 8034
rect 12738 7982 12740 8034
rect 12684 7476 12740 7982
rect 12796 7924 12852 8094
rect 12796 7858 12852 7868
rect 12908 8596 12964 8606
rect 12124 7422 12126 7474
rect 12178 7422 12180 7474
rect 12124 7252 12180 7422
rect 12124 7186 12180 7196
rect 12460 7420 12740 7476
rect 12796 7586 12852 7598
rect 12796 7534 12798 7586
rect 12850 7534 12852 7586
rect 12460 7028 12516 7420
rect 12460 6962 12516 6972
rect 12572 7252 12628 7262
rect 12796 7252 12852 7534
rect 12908 7474 12964 8540
rect 12908 7422 12910 7474
rect 12962 7422 12964 7474
rect 12908 7410 12964 7422
rect 13132 7252 13188 10220
rect 13580 9828 13636 10332
rect 14028 10050 14084 10670
rect 14028 9998 14030 10050
rect 14082 9998 14084 10050
rect 14028 9986 14084 9998
rect 13580 9734 13636 9772
rect 14140 9714 14196 10780
rect 14364 10498 14420 10510
rect 14364 10446 14366 10498
rect 14418 10446 14420 10498
rect 14364 10050 14420 10446
rect 14364 9998 14366 10050
rect 14418 9998 14420 10050
rect 14364 9986 14420 9998
rect 14140 9662 14142 9714
rect 14194 9662 14196 9714
rect 14140 9650 14196 9662
rect 13468 9604 13524 9614
rect 13468 7588 13524 9548
rect 14476 9268 14532 11340
rect 14700 10498 14756 11452
rect 14812 10836 14868 12236
rect 14924 11618 14980 13132
rect 15036 12962 15092 12974
rect 15036 12910 15038 12962
rect 15090 12910 15092 12962
rect 15036 12404 15092 12910
rect 15036 12338 15092 12348
rect 15148 12628 15204 12638
rect 14924 11566 14926 11618
rect 14978 11566 14980 11618
rect 14924 11554 14980 11566
rect 15036 12178 15092 12190
rect 15036 12126 15038 12178
rect 15090 12126 15092 12178
rect 15036 11620 15092 12126
rect 15036 11554 15092 11564
rect 15148 11172 15204 12572
rect 15036 11116 15204 11172
rect 14812 10770 14868 10780
rect 14924 11060 14980 11070
rect 14700 10446 14702 10498
rect 14754 10446 14756 10498
rect 14700 10434 14756 10446
rect 14812 10610 14868 10622
rect 14812 10558 14814 10610
rect 14866 10558 14868 10610
rect 14700 9268 14756 9278
rect 14476 9266 14756 9268
rect 14476 9214 14478 9266
rect 14530 9214 14702 9266
rect 14754 9214 14756 9266
rect 14476 9212 14756 9214
rect 14476 9202 14532 9212
rect 13692 8932 13748 8942
rect 13692 8930 13860 8932
rect 13692 8878 13694 8930
rect 13746 8878 13860 8930
rect 13692 8876 13860 8878
rect 13692 8866 13748 8876
rect 13692 8372 13748 8382
rect 13692 8278 13748 8316
rect 13580 8146 13636 8158
rect 13580 8094 13582 8146
rect 13634 8094 13636 8146
rect 13580 7812 13636 8094
rect 13580 7746 13636 7756
rect 13580 7588 13636 7598
rect 13468 7586 13636 7588
rect 13468 7534 13582 7586
rect 13634 7534 13636 7586
rect 13468 7532 13636 7534
rect 12796 7196 13188 7252
rect 12572 6914 12628 7196
rect 12572 6862 12574 6914
rect 12626 6862 12628 6914
rect 12572 6850 12628 6862
rect 12684 7028 12740 7038
rect 12236 6468 12292 6478
rect 12236 6374 12292 6412
rect 12348 5348 12404 5358
rect 12348 5254 12404 5292
rect 12684 5346 12740 6972
rect 12796 6692 12852 6702
rect 13580 6692 13636 7532
rect 12796 6690 13636 6692
rect 12796 6638 12798 6690
rect 12850 6638 13636 6690
rect 12796 6636 13636 6638
rect 12796 6626 12852 6636
rect 12684 5294 12686 5346
rect 12738 5294 12740 5346
rect 12684 5282 12740 5294
rect 12908 5124 12964 6636
rect 13580 6468 13636 6478
rect 12908 5030 12964 5068
rect 13468 6466 13636 6468
rect 13468 6414 13582 6466
rect 13634 6414 13636 6466
rect 13468 6412 13636 6414
rect 11228 4274 11284 4284
rect 10668 4226 10836 4228
rect 10668 4174 10670 4226
rect 10722 4174 10836 4226
rect 10668 4172 10836 4174
rect 10668 4162 10724 4172
rect 11452 4116 11508 4126
rect 10892 4114 11508 4116
rect 10892 4062 11454 4114
rect 11506 4062 11508 4114
rect 10892 4060 11508 4062
rect 10668 3444 10724 3454
rect 10892 3444 10948 4060
rect 11452 4050 11508 4060
rect 11116 3892 11172 3902
rect 11116 3666 11172 3836
rect 11116 3614 11118 3666
rect 11170 3614 11172 3666
rect 11116 3602 11172 3614
rect 10668 3442 10948 3444
rect 10668 3390 10670 3442
rect 10722 3390 10948 3442
rect 10668 3388 10948 3390
rect 11900 3388 11956 4956
rect 13468 4900 13524 6412
rect 13580 6402 13636 6412
rect 13468 4834 13524 4844
rect 13580 5012 13636 5022
rect 13580 4450 13636 4956
rect 13580 4398 13582 4450
rect 13634 4398 13636 4450
rect 13580 4386 13636 4398
rect 13804 4228 13860 8876
rect 14588 8370 14644 9212
rect 14700 9202 14756 9212
rect 14588 8318 14590 8370
rect 14642 8318 14644 8370
rect 14588 8260 14644 8318
rect 14812 8372 14868 10558
rect 14812 8306 14868 8316
rect 14924 9602 14980 11004
rect 15036 10836 15092 11116
rect 15260 11060 15316 13468
rect 15372 13186 15428 15092
rect 15484 13636 15540 13646
rect 15484 13542 15540 13580
rect 15372 13134 15374 13186
rect 15426 13134 15428 13186
rect 15372 13122 15428 13134
rect 15596 12292 15652 15092
rect 16044 14308 16100 14318
rect 15932 14252 16044 14308
rect 15708 13972 15764 13982
rect 15708 13878 15764 13916
rect 15932 13860 15988 14252
rect 16044 14242 16100 14252
rect 16156 13972 16212 15092
rect 15820 13858 15988 13860
rect 15820 13806 15934 13858
rect 15986 13806 15988 13858
rect 15820 13804 15988 13806
rect 15708 13524 15764 13534
rect 15708 13430 15764 13468
rect 15708 12964 15764 12974
rect 15820 12964 15876 13804
rect 15932 13794 15988 13804
rect 16044 13916 16212 13972
rect 16380 15090 16436 15102
rect 16604 15092 16772 15148
rect 16380 15038 16382 15090
rect 16434 15038 16436 15090
rect 16044 13300 16100 13916
rect 16268 13860 16324 13870
rect 16380 13860 16436 15038
rect 16604 14308 16660 14318
rect 16604 14214 16660 14252
rect 16716 13860 16772 15092
rect 17164 14980 17220 19516
rect 17276 19348 17332 19358
rect 17276 19254 17332 19292
rect 17724 19124 17780 19852
rect 18060 19234 18116 20188
rect 18172 20018 18228 20860
rect 18396 20804 18452 22092
rect 19068 21700 19124 21710
rect 19068 21606 19124 21644
rect 18508 21476 18564 21486
rect 18508 21382 18564 21420
rect 19516 20916 19572 22204
rect 19628 21586 19684 23100
rect 19740 23090 19796 23100
rect 20188 23154 20244 23324
rect 20188 23102 20190 23154
rect 20242 23102 20244 23154
rect 20188 23090 20244 23102
rect 20076 22372 20132 22382
rect 20300 22372 20356 24220
rect 20412 23604 20468 24444
rect 20412 23538 20468 23548
rect 20636 24444 21028 24500
rect 21420 25282 21476 25294
rect 21420 25230 21422 25282
rect 21474 25230 21476 25282
rect 20636 23268 20692 24444
rect 21420 24164 21476 25230
rect 21532 25284 21588 25322
rect 21532 25218 21588 25228
rect 20636 23202 20692 23212
rect 20748 24108 21476 24164
rect 21532 25060 21588 25070
rect 20748 23154 20804 24108
rect 20748 23102 20750 23154
rect 20802 23102 20804 23154
rect 20748 23090 20804 23102
rect 20860 23940 20916 23950
rect 20076 22370 20356 22372
rect 20076 22318 20078 22370
rect 20130 22318 20356 22370
rect 20076 22316 20356 22318
rect 20860 22370 20916 23884
rect 21532 23716 21588 25004
rect 21644 23940 21700 26238
rect 22204 26290 22260 26302
rect 22204 26238 22206 26290
rect 22258 26238 22260 26290
rect 22204 25620 22260 26238
rect 22204 25554 22260 25564
rect 22316 25394 22372 30940
rect 23548 30882 23604 30894
rect 23548 30830 23550 30882
rect 23602 30830 23604 30882
rect 23548 30548 23604 30830
rect 22764 30492 23044 30548
rect 22652 30436 22708 30446
rect 22764 30436 22820 30492
rect 22652 30434 22820 30436
rect 22652 30382 22654 30434
rect 22706 30382 22820 30434
rect 22652 30380 22820 30382
rect 22652 30370 22708 30380
rect 22876 30324 22932 30334
rect 22764 30268 22876 30324
rect 22428 29986 22484 29998
rect 22428 29934 22430 29986
rect 22482 29934 22484 29986
rect 22428 29876 22484 29934
rect 22428 29810 22484 29820
rect 22428 29652 22484 29662
rect 22428 29540 22484 29596
rect 22540 29540 22596 29550
rect 22428 29538 22596 29540
rect 22428 29486 22542 29538
rect 22594 29486 22596 29538
rect 22428 29484 22596 29486
rect 22428 28642 22484 29484
rect 22540 29474 22596 29484
rect 22428 28590 22430 28642
rect 22482 28590 22484 28642
rect 22428 28578 22484 28590
rect 22652 28756 22708 28766
rect 22652 28530 22708 28700
rect 22652 28478 22654 28530
rect 22706 28478 22708 28530
rect 22652 28466 22708 28478
rect 22428 28084 22484 28094
rect 22428 27990 22484 28028
rect 22540 27300 22596 27310
rect 22428 25508 22484 25518
rect 22428 25414 22484 25452
rect 22316 25342 22318 25394
rect 22370 25342 22372 25394
rect 22316 25330 22372 25342
rect 21756 25284 21812 25294
rect 22092 25284 22148 25294
rect 21756 25282 22148 25284
rect 21756 25230 21758 25282
rect 21810 25230 22094 25282
rect 22146 25230 22148 25282
rect 21756 25228 22148 25230
rect 21756 25218 21812 25228
rect 22092 25218 22148 25228
rect 22204 25284 22260 25294
rect 21644 23874 21700 23884
rect 21756 25060 21812 25070
rect 21532 23660 21700 23716
rect 20860 22318 20862 22370
rect 20914 22318 20916 22370
rect 20076 22306 20132 22316
rect 20860 22260 20916 22318
rect 20860 22194 20916 22204
rect 21308 22484 21364 22494
rect 20636 22148 20692 22158
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20300 21700 20356 21710
rect 19628 21534 19630 21586
rect 19682 21534 19684 21586
rect 19628 21522 19684 21534
rect 20188 21644 20300 21700
rect 20188 21586 20244 21644
rect 20300 21634 20356 21644
rect 20188 21534 20190 21586
rect 20242 21534 20244 21586
rect 20188 21522 20244 21534
rect 20524 21476 20580 21486
rect 20524 21382 20580 21420
rect 20636 20916 20692 22092
rect 21084 21700 21140 21710
rect 21084 21606 21140 21644
rect 19516 20822 19572 20860
rect 20412 20914 20692 20916
rect 20412 20862 20638 20914
rect 20690 20862 20692 20914
rect 20412 20860 20692 20862
rect 18396 20738 18452 20748
rect 18172 19966 18174 20018
rect 18226 19966 18228 20018
rect 18172 19954 18228 19966
rect 18396 20580 18452 20590
rect 18060 19182 18062 19234
rect 18114 19182 18116 19234
rect 18060 19170 18116 19182
rect 18284 19348 18340 19358
rect 17836 19124 17892 19134
rect 17724 19068 17836 19124
rect 17836 19058 17892 19068
rect 17948 18450 18004 18462
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17724 18226 17780 18238
rect 17724 18174 17726 18226
rect 17778 18174 17780 18226
rect 17388 17668 17444 17678
rect 17388 17574 17444 17612
rect 17612 17666 17668 17678
rect 17612 17614 17614 17666
rect 17666 17614 17668 17666
rect 17500 17332 17556 17342
rect 17500 16996 17556 17276
rect 17612 17220 17668 17614
rect 17612 17154 17668 17164
rect 17612 16996 17668 17006
rect 17500 16994 17668 16996
rect 17500 16942 17614 16994
rect 17666 16942 17668 16994
rect 17500 16940 17668 16942
rect 17612 16930 17668 16940
rect 17612 16548 17668 16558
rect 17612 16100 17668 16492
rect 17724 16324 17780 18174
rect 17948 17890 18004 18398
rect 18284 18450 18340 19292
rect 18284 18398 18286 18450
rect 18338 18398 18340 18450
rect 18284 18386 18340 18398
rect 18396 18338 18452 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20412 20244 20468 20860
rect 20636 20850 20692 20860
rect 18396 18286 18398 18338
rect 18450 18286 18452 18338
rect 18396 18116 18452 18286
rect 18396 18050 18452 18060
rect 18844 19906 18900 19918
rect 18844 19854 18846 19906
rect 18898 19854 18900 19906
rect 17948 17838 17950 17890
rect 18002 17838 18004 17890
rect 17948 17826 18004 17838
rect 18284 17668 18340 17678
rect 18172 17612 18284 17668
rect 18060 16996 18116 17006
rect 17836 16884 17892 16894
rect 17836 16790 17892 16828
rect 18060 16882 18116 16940
rect 18060 16830 18062 16882
rect 18114 16830 18116 16882
rect 17724 16258 17780 16268
rect 17612 16006 17668 16044
rect 17948 15988 18004 15998
rect 17948 15894 18004 15932
rect 18060 15148 18116 16830
rect 18172 16884 18228 17612
rect 18284 17602 18340 17612
rect 18732 17666 18788 17678
rect 18732 17614 18734 17666
rect 18786 17614 18788 17666
rect 18284 17444 18340 17454
rect 18284 17442 18452 17444
rect 18284 17390 18286 17442
rect 18338 17390 18452 17442
rect 18284 17388 18452 17390
rect 18284 17378 18340 17388
rect 18284 17108 18340 17118
rect 18284 17014 18340 17052
rect 18284 16884 18340 16894
rect 18172 16828 18284 16884
rect 18396 16884 18452 17388
rect 18732 17332 18788 17614
rect 18732 17266 18788 17276
rect 18844 16996 18900 19854
rect 19964 19346 20020 19358
rect 19964 19294 19966 19346
rect 20018 19294 20020 19346
rect 19964 19124 20020 19294
rect 19964 19058 20020 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19292 18562 19348 18574
rect 19292 18510 19294 18562
rect 19346 18510 19348 18562
rect 18956 17892 19012 17902
rect 18956 17798 19012 17836
rect 19180 17780 19236 17790
rect 19180 17686 19236 17724
rect 19292 17668 19348 18510
rect 19628 18452 19684 18462
rect 19404 18396 19628 18452
rect 19404 17778 19460 18396
rect 19628 18358 19684 18396
rect 20412 18450 20468 20188
rect 21308 20020 21364 22428
rect 21532 20578 21588 20590
rect 21532 20526 21534 20578
rect 21586 20526 21588 20578
rect 21532 20356 21588 20526
rect 21644 20580 21700 23660
rect 21756 21812 21812 25004
rect 21868 24948 21924 24958
rect 21868 22372 21924 24892
rect 22092 24164 22148 24174
rect 22204 24164 22260 25228
rect 22092 24162 22260 24164
rect 22092 24110 22094 24162
rect 22146 24110 22260 24162
rect 22092 24108 22260 24110
rect 22092 24098 22148 24108
rect 22204 23826 22260 23838
rect 22204 23774 22206 23826
rect 22258 23774 22260 23826
rect 22204 23380 22260 23774
rect 22540 23716 22596 27244
rect 22764 26908 22820 30268
rect 22876 30258 22932 30268
rect 22876 30100 22932 30110
rect 22988 30100 23044 30492
rect 23548 30482 23604 30492
rect 23996 30324 24052 32172
rect 24108 30994 24164 32844
rect 24108 30942 24110 30994
rect 24162 30942 24164 30994
rect 24108 30548 24164 30942
rect 24108 30482 24164 30492
rect 24220 31668 24276 31678
rect 24444 31668 24500 33966
rect 24556 33572 24612 33582
rect 24556 33478 24612 33516
rect 24892 33348 24948 35308
rect 25452 35252 25508 35756
rect 26012 36258 26404 36260
rect 26012 36206 26350 36258
rect 26402 36206 26404 36258
rect 26012 36204 26404 36206
rect 25452 35186 25508 35196
rect 25676 35586 25732 35598
rect 25676 35534 25678 35586
rect 25730 35534 25732 35586
rect 25004 35028 25060 35038
rect 25004 34914 25060 34972
rect 25004 34862 25006 34914
rect 25058 34862 25060 34914
rect 25004 34850 25060 34862
rect 25116 34916 25172 34926
rect 25116 34822 25172 34860
rect 25676 34916 25732 35534
rect 25676 34850 25732 34860
rect 25900 35028 25956 35038
rect 25452 34804 25508 34814
rect 25452 34710 25508 34748
rect 25340 34690 25396 34702
rect 25340 34638 25342 34690
rect 25394 34638 25396 34690
rect 25340 34580 25396 34638
rect 25788 34692 25844 34702
rect 25788 34598 25844 34636
rect 25340 34524 25732 34580
rect 25452 34244 25508 34254
rect 25452 34130 25508 34188
rect 25452 34078 25454 34130
rect 25506 34078 25508 34130
rect 25452 34066 25508 34078
rect 25564 34242 25620 34254
rect 25564 34190 25566 34242
rect 25618 34190 25620 34242
rect 25564 33796 25620 34190
rect 25004 33740 25620 33796
rect 25004 33570 25060 33740
rect 25004 33518 25006 33570
rect 25058 33518 25060 33570
rect 25004 33506 25060 33518
rect 25340 33348 25396 33358
rect 24892 33292 25060 33348
rect 24220 31666 24500 31668
rect 24220 31614 24222 31666
rect 24274 31614 24500 31666
rect 24220 31612 24500 31614
rect 24892 33124 24948 33134
rect 24220 30324 24276 31612
rect 24668 31220 24724 31230
rect 24668 31126 24724 31164
rect 24444 30994 24500 31006
rect 24444 30942 24446 30994
rect 24498 30942 24500 30994
rect 23996 30268 24276 30324
rect 24332 30770 24388 30782
rect 24332 30718 24334 30770
rect 24386 30718 24388 30770
rect 22876 30098 23044 30100
rect 22876 30046 22878 30098
rect 22930 30046 23044 30098
rect 22876 30044 23044 30046
rect 23100 30210 23156 30222
rect 23100 30158 23102 30210
rect 23154 30158 23156 30210
rect 22876 30034 22932 30044
rect 22876 29426 22932 29438
rect 22876 29374 22878 29426
rect 22930 29374 22932 29426
rect 22876 28756 22932 29374
rect 23100 28756 23156 30158
rect 23212 30212 23268 30222
rect 23212 29652 23268 30156
rect 23660 29988 23716 29998
rect 23660 29986 23828 29988
rect 23660 29934 23662 29986
rect 23714 29934 23828 29986
rect 23660 29932 23828 29934
rect 23660 29922 23716 29932
rect 23212 29558 23268 29596
rect 23436 29426 23492 29438
rect 23436 29374 23438 29426
rect 23490 29374 23492 29426
rect 23436 29092 23492 29374
rect 23436 29026 23492 29036
rect 23548 28868 23604 28878
rect 22876 28700 23380 28756
rect 23212 27300 23268 27310
rect 22764 26852 22932 26908
rect 22540 23650 22596 23660
rect 22204 23314 22260 23324
rect 21980 22372 22036 22382
rect 21868 22316 21980 22372
rect 21980 22278 22036 22316
rect 22540 22146 22596 22158
rect 22540 22094 22542 22146
rect 22594 22094 22596 22146
rect 22540 22036 22596 22094
rect 22540 21970 22596 21980
rect 21756 21756 22148 21812
rect 22092 20916 22148 21756
rect 22204 21700 22260 21710
rect 22204 21606 22260 21644
rect 22540 21586 22596 21598
rect 22540 21534 22542 21586
rect 22594 21534 22596 21586
rect 22092 20914 22372 20916
rect 22092 20862 22094 20914
rect 22146 20862 22372 20914
rect 22092 20860 22372 20862
rect 22092 20850 22148 20860
rect 22316 20802 22372 20860
rect 22316 20750 22318 20802
rect 22370 20750 22372 20802
rect 22316 20738 22372 20750
rect 22540 20804 22596 21534
rect 22876 21474 22932 26852
rect 23100 25620 23156 25630
rect 23100 25526 23156 25564
rect 23212 25506 23268 27244
rect 23212 25454 23214 25506
rect 23266 25454 23268 25506
rect 23212 25442 23268 25454
rect 22988 25396 23044 25406
rect 22988 25302 23044 25340
rect 23324 24164 23380 28700
rect 23548 28642 23604 28812
rect 23548 28590 23550 28642
rect 23602 28590 23604 28642
rect 23548 28578 23604 28590
rect 23660 28644 23716 28654
rect 23660 28550 23716 28588
rect 23660 28084 23716 28094
rect 23772 28084 23828 29932
rect 23884 29652 23940 29662
rect 23884 29426 23940 29596
rect 23884 29374 23886 29426
rect 23938 29374 23940 29426
rect 23884 29362 23940 29374
rect 23884 28530 23940 28542
rect 23884 28478 23886 28530
rect 23938 28478 23940 28530
rect 23884 28420 23940 28478
rect 23884 28354 23940 28364
rect 23716 28028 23828 28084
rect 23660 28018 23716 28028
rect 23996 27860 24052 30268
rect 24332 29650 24388 30718
rect 24444 30772 24500 30942
rect 24444 30706 24500 30716
rect 24892 30324 24948 33068
rect 24892 30258 24948 30268
rect 25004 30212 25060 33292
rect 25228 33292 25340 33348
rect 25004 30146 25060 30156
rect 25116 31554 25172 31566
rect 25116 31502 25118 31554
rect 25170 31502 25172 31554
rect 25116 30772 25172 31502
rect 25228 31108 25284 33292
rect 25340 33254 25396 33292
rect 25452 31556 25508 31566
rect 25452 31462 25508 31500
rect 25228 30994 25284 31052
rect 25228 30942 25230 30994
rect 25282 30942 25284 30994
rect 25228 30930 25284 30942
rect 25452 31220 25508 31230
rect 25676 31220 25732 34524
rect 25900 34356 25956 34972
rect 25900 34290 25956 34300
rect 25900 34020 25956 34030
rect 25676 31164 25844 31220
rect 25452 30994 25508 31164
rect 25452 30942 25454 30994
rect 25506 30942 25508 30994
rect 25452 30930 25508 30942
rect 24332 29598 24334 29650
rect 24386 29598 24388 29650
rect 24332 29586 24388 29598
rect 24556 29988 24612 29998
rect 24892 29988 24948 29998
rect 24612 29986 24948 29988
rect 24612 29934 24894 29986
rect 24946 29934 24948 29986
rect 24612 29932 24948 29934
rect 24332 29428 24388 29438
rect 24556 29428 24612 29932
rect 24892 29922 24948 29932
rect 24332 29426 24612 29428
rect 24332 29374 24334 29426
rect 24386 29374 24612 29426
rect 24332 29372 24612 29374
rect 24668 29426 24724 29438
rect 24668 29374 24670 29426
rect 24722 29374 24724 29426
rect 24220 29204 24276 29214
rect 24220 29110 24276 29148
rect 24332 28868 24388 29372
rect 24220 28812 24388 28868
rect 24108 28532 24164 28542
rect 24108 28438 24164 28476
rect 24108 28084 24164 28094
rect 24108 27990 24164 28028
rect 23660 27804 24052 27860
rect 23660 26962 23716 27804
rect 23660 26910 23662 26962
rect 23714 26910 23716 26962
rect 23660 26898 23716 26910
rect 23772 26962 23828 26974
rect 23772 26910 23774 26962
rect 23826 26910 23828 26962
rect 23436 26852 23492 26862
rect 23436 26850 23604 26852
rect 23436 26798 23438 26850
rect 23490 26798 23604 26850
rect 23436 26796 23604 26798
rect 23436 26786 23492 26796
rect 23548 25506 23604 26796
rect 23548 25454 23550 25506
rect 23602 25454 23604 25506
rect 23548 25442 23604 25454
rect 23772 25508 23828 26910
rect 24220 26908 24276 28812
rect 24332 28642 24388 28654
rect 24332 28590 24334 28642
rect 24386 28590 24388 28642
rect 24332 28084 24388 28590
rect 24668 28420 24724 29374
rect 25004 28644 25060 28654
rect 25004 28550 25060 28588
rect 25116 28420 25172 30716
rect 25676 30770 25732 30782
rect 25676 30718 25678 30770
rect 25730 30718 25732 30770
rect 25676 30660 25732 30718
rect 25676 30594 25732 30604
rect 25228 29428 25284 29466
rect 25228 29362 25284 29372
rect 25228 29204 25284 29214
rect 25564 29204 25620 29214
rect 25228 29110 25284 29148
rect 25340 29148 25564 29204
rect 24332 28018 24388 28028
rect 24444 28364 24668 28420
rect 24444 27300 24500 28364
rect 24668 28354 24724 28364
rect 25004 28364 25172 28420
rect 24444 27206 24500 27244
rect 23772 25442 23828 25452
rect 24108 26852 24276 26908
rect 24556 26962 24612 26974
rect 24556 26910 24558 26962
rect 24610 26910 24612 26962
rect 23996 25396 24052 25406
rect 23996 24946 24052 25340
rect 24108 25284 24164 26852
rect 24556 26516 24612 26910
rect 24668 26516 24724 26526
rect 24556 26514 24724 26516
rect 24556 26462 24670 26514
rect 24722 26462 24724 26514
rect 24556 26460 24724 26462
rect 24668 26450 24724 26460
rect 24556 25732 24612 25742
rect 24220 25620 24276 25630
rect 24556 25620 24612 25676
rect 24220 25618 24612 25620
rect 24220 25566 24222 25618
rect 24274 25566 24612 25618
rect 24220 25564 24612 25566
rect 24220 25554 24276 25564
rect 24444 25396 24500 25406
rect 24444 25302 24500 25340
rect 24556 25394 24612 25564
rect 24556 25342 24558 25394
rect 24610 25342 24612 25394
rect 24556 25330 24612 25342
rect 24780 25284 24836 25294
rect 24108 25228 24388 25284
rect 23996 24894 23998 24946
rect 24050 24894 24052 24946
rect 23996 24882 24052 24894
rect 24220 24836 24276 24874
rect 24220 24770 24276 24780
rect 23212 24108 23380 24164
rect 24108 24610 24164 24622
rect 24108 24558 24110 24610
rect 24162 24558 24164 24610
rect 23100 23380 23156 23390
rect 23100 23286 23156 23324
rect 22988 22370 23044 22382
rect 22988 22318 22990 22370
rect 23042 22318 23044 22370
rect 22988 22036 23044 22318
rect 22988 21970 23044 21980
rect 22876 21422 22878 21474
rect 22930 21422 22932 21474
rect 22876 21364 22932 21422
rect 22876 21298 22932 21308
rect 22988 20804 23044 20814
rect 23212 20804 23268 24108
rect 23324 23940 23380 23950
rect 23324 23846 23380 23884
rect 24108 23938 24164 24558
rect 24332 23940 24388 25228
rect 24668 25282 24836 25284
rect 24668 25230 24782 25282
rect 24834 25230 24836 25282
rect 24668 25228 24836 25230
rect 24668 24722 24724 25228
rect 24780 25218 24836 25228
rect 24668 24670 24670 24722
rect 24722 24670 24724 24722
rect 24668 24658 24724 24670
rect 25004 24724 25060 28364
rect 25340 28082 25396 29148
rect 25564 29110 25620 29148
rect 25564 28756 25620 28766
rect 25340 28030 25342 28082
rect 25394 28030 25396 28082
rect 25340 28018 25396 28030
rect 25452 28532 25508 28542
rect 25452 28082 25508 28476
rect 25452 28030 25454 28082
rect 25506 28030 25508 28082
rect 25452 28018 25508 28030
rect 25564 27634 25620 28700
rect 25564 27582 25566 27634
rect 25618 27582 25620 27634
rect 25564 27300 25620 27582
rect 25676 27300 25732 27310
rect 25564 27244 25676 27300
rect 25676 27234 25732 27244
rect 25116 26962 25172 26974
rect 25116 26910 25118 26962
rect 25170 26910 25172 26962
rect 25116 26908 25172 26910
rect 25788 26908 25844 31164
rect 25116 26852 25284 26908
rect 25228 26290 25284 26852
rect 25228 26238 25230 26290
rect 25282 26238 25284 26290
rect 25228 26068 25284 26238
rect 25228 26002 25284 26012
rect 25340 26852 25844 26908
rect 25340 25506 25396 26852
rect 25340 25454 25342 25506
rect 25394 25454 25396 25506
rect 25340 25442 25396 25454
rect 25564 25956 25620 25966
rect 25564 25506 25620 25900
rect 25564 25454 25566 25506
rect 25618 25454 25620 25506
rect 25564 25442 25620 25454
rect 25900 25730 25956 33964
rect 26012 31778 26068 36204
rect 26348 36194 26404 36204
rect 26460 35924 26516 36428
rect 26572 36372 26628 36382
rect 26572 36278 26628 36316
rect 26460 35810 26516 35868
rect 26684 35812 26740 37998
rect 26908 36596 26964 39340
rect 27132 39330 27188 39340
rect 27244 40962 27300 40974
rect 27244 40910 27246 40962
rect 27298 40910 27300 40962
rect 27244 39396 27300 40910
rect 27356 40402 27412 41132
rect 27804 41188 27860 41918
rect 27804 41122 27860 41132
rect 27356 40350 27358 40402
rect 27410 40350 27412 40402
rect 27356 40338 27412 40350
rect 27916 40402 27972 40414
rect 27916 40350 27918 40402
rect 27970 40350 27972 40402
rect 27916 39506 27972 40350
rect 28140 39844 28196 43652
rect 28252 43650 28308 43662
rect 28252 43598 28254 43650
rect 28306 43598 28308 43650
rect 28252 41970 28308 43598
rect 28700 43540 28756 43550
rect 28700 43446 28756 43484
rect 28252 41918 28254 41970
rect 28306 41918 28308 41970
rect 28252 41906 28308 41918
rect 29036 43314 29092 45276
rect 29260 44884 29316 44894
rect 29260 43650 29316 44828
rect 29260 43598 29262 43650
rect 29314 43598 29316 43650
rect 29260 43586 29316 43598
rect 29036 43262 29038 43314
rect 29090 43262 29092 43314
rect 29036 41076 29092 43262
rect 29372 41188 29428 47404
rect 30716 47012 30772 48076
rect 30828 48020 30884 48300
rect 32172 48356 32228 48750
rect 32172 48290 32228 48300
rect 30828 47954 30884 47964
rect 32396 48130 32452 48972
rect 32620 48962 32676 48972
rect 32732 48916 32788 49756
rect 32844 49028 32900 49870
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 33292 49028 33348 49038
rect 32844 49026 33348 49028
rect 32844 48974 33294 49026
rect 33346 48974 33348 49026
rect 32844 48972 33348 48974
rect 33292 48962 33348 48972
rect 37100 49026 37156 49038
rect 37100 48974 37102 49026
rect 37154 48974 37156 49026
rect 32732 48860 33236 48916
rect 33180 48466 33236 48860
rect 33180 48414 33182 48466
rect 33234 48414 33236 48466
rect 33180 48402 33236 48414
rect 35756 48802 35812 48814
rect 35756 48750 35758 48802
rect 35810 48750 35812 48802
rect 32396 48078 32398 48130
rect 32450 48078 32452 48130
rect 32284 47460 32340 47470
rect 32172 47404 32284 47460
rect 32396 47460 32452 48078
rect 33740 48354 33796 48366
rect 33740 48302 33742 48354
rect 33794 48302 33796 48354
rect 33740 48132 33796 48302
rect 34076 48354 34132 48366
rect 34076 48302 34078 48354
rect 34130 48302 34132 48354
rect 34076 48244 34132 48302
rect 34076 48178 34132 48188
rect 35756 48244 35812 48750
rect 33516 48020 33572 48030
rect 33404 48018 33572 48020
rect 33404 47966 33518 48018
rect 33570 47966 33572 48018
rect 33404 47964 33572 47966
rect 32620 47460 32676 47470
rect 32396 47458 32676 47460
rect 32396 47406 32622 47458
rect 32674 47406 32676 47458
rect 32396 47404 32676 47406
rect 31836 47348 31892 47358
rect 30716 46946 30772 46956
rect 31276 47346 31892 47348
rect 31276 47294 31838 47346
rect 31890 47294 31892 47346
rect 31276 47292 31892 47294
rect 31276 46898 31332 47292
rect 31836 47282 31892 47292
rect 32172 47346 32228 47404
rect 32284 47394 32340 47404
rect 32172 47294 32174 47346
rect 32226 47294 32228 47346
rect 32172 47282 32228 47294
rect 32620 47236 32676 47404
rect 33068 47460 33124 47470
rect 33068 47366 33124 47404
rect 32620 47170 32676 47180
rect 31276 46846 31278 46898
rect 31330 46846 31332 46898
rect 31276 46834 31332 46846
rect 30156 46788 30212 46798
rect 30156 46562 30212 46732
rect 31948 46788 32004 46798
rect 31948 46694 32004 46732
rect 32396 46788 32452 46798
rect 32396 46694 32452 46732
rect 33404 46788 33460 47964
rect 33516 47954 33572 47964
rect 33404 46722 33460 46732
rect 33516 47236 33572 47246
rect 30156 46510 30158 46562
rect 30210 46510 30212 46562
rect 30156 46498 30212 46510
rect 30604 46674 30660 46686
rect 30604 46622 30606 46674
rect 30658 46622 30660 46674
rect 29932 45332 29988 45342
rect 29932 45238 29988 45276
rect 30268 45220 30324 45230
rect 30156 45108 30212 45118
rect 30156 44436 30212 45052
rect 30268 45106 30324 45164
rect 30604 45220 30660 46622
rect 31612 46450 31668 46462
rect 31612 46398 31614 46450
rect 31666 46398 31668 46450
rect 31500 45332 31556 45342
rect 30604 45154 30660 45164
rect 31164 45330 31556 45332
rect 31164 45278 31502 45330
rect 31554 45278 31556 45330
rect 31164 45276 31556 45278
rect 30268 45054 30270 45106
rect 30322 45054 30324 45106
rect 30268 44996 30324 45054
rect 30268 44930 30324 44940
rect 30716 44994 30772 45006
rect 30716 44942 30718 44994
rect 30770 44942 30772 44994
rect 30716 44884 30772 44942
rect 30156 44434 30548 44436
rect 30156 44382 30158 44434
rect 30210 44382 30548 44434
rect 30156 44380 30548 44382
rect 30156 44370 30212 44380
rect 30492 44322 30548 44380
rect 30492 44270 30494 44322
rect 30546 44270 30548 44322
rect 30492 44258 30548 44270
rect 30716 44324 30772 44828
rect 30716 44258 30772 44268
rect 31164 44322 31220 45276
rect 31500 45266 31556 45276
rect 31164 44270 31166 44322
rect 31218 44270 31220 44322
rect 31164 44258 31220 44270
rect 31276 45106 31332 45118
rect 31276 45054 31278 45106
rect 31330 45054 31332 45106
rect 30604 43764 30660 43774
rect 29820 43650 29876 43662
rect 29820 43598 29822 43650
rect 29874 43598 29876 43650
rect 29820 43316 29876 43598
rect 29820 41860 29876 43260
rect 30044 41860 30100 41870
rect 29820 41804 30044 41860
rect 29596 41188 29652 41198
rect 29372 41132 29596 41188
rect 29036 41020 29428 41076
rect 28140 39788 28308 39844
rect 27916 39454 27918 39506
rect 27970 39454 27972 39506
rect 27916 39442 27972 39454
rect 28140 39618 28196 39630
rect 28140 39566 28142 39618
rect 28194 39566 28196 39618
rect 27468 39396 27524 39406
rect 27244 39340 27468 39396
rect 27244 38834 27300 39340
rect 27468 39302 27524 39340
rect 28140 39058 28196 39566
rect 28140 39006 28142 39058
rect 28194 39006 28196 39058
rect 28140 38994 28196 39006
rect 27244 38782 27246 38834
rect 27298 38782 27300 38834
rect 27244 38770 27300 38782
rect 27692 38724 27748 38734
rect 27804 38724 27860 38734
rect 27692 38722 27804 38724
rect 27692 38670 27694 38722
rect 27746 38670 27804 38722
rect 27692 38668 27804 38670
rect 28252 38668 28308 39788
rect 27692 38658 27748 38668
rect 27804 38612 28084 38668
rect 27468 38388 27524 38398
rect 27468 38050 27524 38332
rect 27804 38162 27860 38174
rect 27804 38110 27806 38162
rect 27858 38110 27860 38162
rect 27468 37998 27470 38050
rect 27522 37998 27524 38050
rect 27020 37268 27076 37278
rect 27020 37174 27076 37212
rect 27468 37268 27524 37998
rect 27692 38052 27748 38062
rect 27692 37958 27748 37996
rect 27468 37202 27524 37212
rect 27580 37492 27636 37502
rect 27356 37044 27412 37054
rect 26908 36530 26964 36540
rect 27020 36932 27076 36942
rect 27020 36260 27076 36876
rect 27020 36258 27188 36260
rect 27020 36206 27022 36258
rect 27074 36206 27188 36258
rect 27020 36204 27188 36206
rect 27020 36194 27076 36204
rect 26460 35758 26462 35810
rect 26514 35758 26516 35810
rect 26460 35746 26516 35758
rect 26572 35756 26740 35812
rect 26124 35586 26180 35598
rect 26124 35534 26126 35586
rect 26178 35534 26180 35586
rect 26124 35252 26180 35534
rect 26124 35028 26180 35196
rect 26236 35028 26292 35038
rect 26124 35026 26292 35028
rect 26124 34974 26238 35026
rect 26290 34974 26292 35026
rect 26124 34972 26292 34974
rect 26236 34962 26292 34972
rect 26572 34468 26628 35756
rect 26684 35588 26740 35598
rect 26684 35494 26740 35532
rect 27020 35474 27076 35486
rect 27020 35422 27022 35474
rect 27074 35422 27076 35474
rect 26684 35252 26740 35262
rect 26684 34914 26740 35196
rect 26684 34862 26686 34914
rect 26738 34862 26740 34914
rect 26684 34850 26740 34862
rect 26908 34916 26964 34926
rect 26572 34412 26852 34468
rect 26236 34244 26292 34254
rect 26684 34244 26740 34254
rect 26236 34242 26628 34244
rect 26236 34190 26238 34242
rect 26290 34190 26628 34242
rect 26236 34188 26628 34190
rect 26236 34178 26292 34188
rect 26236 34020 26292 34030
rect 26236 33926 26292 33964
rect 26236 32564 26292 32574
rect 26236 32470 26292 32508
rect 26012 31726 26014 31778
rect 26066 31726 26068 31778
rect 26012 31714 26068 31726
rect 26124 31666 26180 31678
rect 26124 31614 26126 31666
rect 26178 31614 26180 31666
rect 26124 31218 26180 31614
rect 26124 31166 26126 31218
rect 26178 31166 26180 31218
rect 26124 31154 26180 31166
rect 26460 31108 26516 31118
rect 26460 31014 26516 31052
rect 26572 30322 26628 34188
rect 26684 34130 26740 34188
rect 26684 34078 26686 34130
rect 26738 34078 26740 34130
rect 26684 34066 26740 34078
rect 26796 34132 26852 34412
rect 26908 34356 26964 34860
rect 27020 34914 27076 35422
rect 27020 34862 27022 34914
rect 27074 34862 27076 34914
rect 27020 34850 27076 34862
rect 27132 34580 27188 36204
rect 27356 35308 27412 36988
rect 27580 37044 27636 37436
rect 27580 36482 27636 36988
rect 27580 36430 27582 36482
rect 27634 36430 27636 36482
rect 27468 35588 27524 35598
rect 27468 35494 27524 35532
rect 27244 35252 27524 35308
rect 27244 34858 27300 35252
rect 27468 35186 27524 35196
rect 27244 34806 27246 34858
rect 27298 34806 27300 34858
rect 27468 34916 27524 34926
rect 27468 34822 27524 34860
rect 27244 34794 27300 34806
rect 27356 34802 27412 34814
rect 27356 34750 27358 34802
rect 27410 34750 27412 34802
rect 27132 34524 27300 34580
rect 26908 34290 26964 34300
rect 26796 34076 26964 34132
rect 26796 33122 26852 33134
rect 26796 33070 26798 33122
rect 26850 33070 26852 33122
rect 26796 32562 26852 33070
rect 26796 32510 26798 32562
rect 26850 32510 26852 32562
rect 26796 32498 26852 32510
rect 26908 32340 26964 34076
rect 27132 33460 27188 33470
rect 26796 32284 26964 32340
rect 27020 33404 27132 33460
rect 26572 30270 26574 30322
rect 26626 30270 26628 30322
rect 26572 30258 26628 30270
rect 26684 31666 26740 31678
rect 26684 31614 26686 31666
rect 26738 31614 26740 31666
rect 26684 30210 26740 31614
rect 26684 30158 26686 30210
rect 26738 30158 26740 30210
rect 26684 30146 26740 30158
rect 26236 29988 26292 29998
rect 26236 29894 26292 29932
rect 26012 29428 26068 29438
rect 26012 29334 26068 29372
rect 26012 28868 26068 28878
rect 26012 27970 26068 28812
rect 26012 27918 26014 27970
rect 26066 27918 26068 27970
rect 26012 27906 26068 27918
rect 26348 27858 26404 27870
rect 26348 27806 26350 27858
rect 26402 27806 26404 27858
rect 26124 27748 26180 27758
rect 26124 27654 26180 27692
rect 25900 25678 25902 25730
rect 25954 25678 25956 25730
rect 25452 25284 25508 25294
rect 25004 24658 25060 24668
rect 25340 25282 25508 25284
rect 25340 25230 25454 25282
rect 25506 25230 25508 25282
rect 25340 25228 25508 25230
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 24108 23874 24164 23886
rect 24220 23884 24388 23940
rect 22540 20802 23268 20804
rect 22540 20750 22990 20802
rect 23042 20750 23268 20802
rect 22540 20748 23268 20750
rect 23324 23604 23380 23614
rect 21756 20580 21812 20590
rect 21644 20524 21756 20580
rect 21756 20514 21812 20524
rect 22428 20578 22484 20590
rect 22428 20526 22430 20578
rect 22482 20526 22484 20578
rect 21532 20290 21588 20300
rect 22428 20356 22484 20526
rect 22428 20290 22484 20300
rect 22652 20578 22708 20590
rect 22652 20526 22654 20578
rect 22706 20526 22708 20578
rect 22540 20020 22596 20030
rect 21084 20018 21364 20020
rect 21084 19966 21310 20018
rect 21362 19966 21364 20018
rect 21084 19964 21364 19966
rect 20972 19908 21028 19918
rect 20972 19814 21028 19852
rect 21084 19684 21140 19964
rect 21308 19954 21364 19964
rect 21980 20018 22596 20020
rect 21980 19966 22542 20018
rect 22594 19966 22596 20018
rect 21980 19964 22596 19966
rect 20748 19628 21140 19684
rect 21980 19908 22036 19964
rect 22540 19954 22596 19964
rect 22652 20020 22708 20526
rect 22652 19954 22708 19964
rect 22764 20580 22820 20590
rect 20748 19346 20804 19628
rect 20748 19294 20750 19346
rect 20802 19294 20804 19346
rect 20748 19282 20804 19294
rect 20412 18398 20414 18450
rect 20466 18398 20468 18450
rect 20412 18386 20468 18398
rect 21420 19234 21476 19246
rect 21420 19182 21422 19234
rect 21474 19182 21476 19234
rect 20860 18338 20916 18350
rect 20860 18286 20862 18338
rect 20914 18286 20916 18338
rect 20860 18116 20916 18286
rect 20860 18050 20916 18060
rect 19404 17726 19406 17778
rect 19458 17726 19460 17778
rect 19404 17714 19460 17726
rect 19292 17602 19348 17612
rect 20412 17668 20468 17678
rect 21196 17668 21252 17678
rect 20412 17666 21252 17668
rect 20412 17614 20414 17666
rect 20466 17614 21198 17666
rect 21250 17614 21252 17666
rect 20412 17612 21252 17614
rect 20412 17602 20468 17612
rect 21196 17602 21252 17612
rect 20076 17554 20132 17566
rect 20076 17502 20078 17554
rect 20130 17502 20132 17554
rect 20076 17444 20132 17502
rect 20076 17378 20132 17388
rect 20188 17442 20244 17454
rect 20188 17390 20190 17442
rect 20242 17390 20244 17442
rect 19628 17332 19684 17342
rect 20188 17332 20244 17390
rect 19068 17108 19124 17118
rect 19068 17014 19124 17052
rect 18844 16940 19012 16996
rect 18396 16828 18788 16884
rect 18284 16790 18340 16828
rect 18732 16772 18788 16828
rect 18844 16772 18900 16782
rect 18732 16770 18900 16772
rect 18732 16718 18846 16770
rect 18898 16718 18900 16770
rect 18732 16716 18900 16718
rect 18844 16706 18900 16716
rect 18508 16660 18564 16670
rect 18508 15986 18564 16604
rect 18620 16658 18676 16670
rect 18620 16606 18622 16658
rect 18674 16606 18676 16658
rect 18620 16436 18676 16606
rect 18620 16370 18676 16380
rect 18956 16212 19012 16940
rect 18508 15934 18510 15986
rect 18562 15934 18564 15986
rect 18508 15922 18564 15934
rect 18620 16156 19012 16212
rect 19068 16884 19124 16894
rect 18620 15148 18676 16156
rect 18956 15988 19012 15998
rect 18060 15092 18228 15148
rect 17164 14914 17220 14924
rect 17276 14644 17332 14654
rect 17164 14532 17220 14542
rect 17164 14438 17220 14476
rect 17276 14530 17332 14588
rect 17276 14478 17278 14530
rect 17330 14478 17332 14530
rect 17276 14466 17332 14478
rect 17724 14532 17780 14542
rect 17724 14438 17780 14476
rect 17052 14420 17108 14430
rect 17052 14326 17108 14364
rect 17388 14420 17444 14430
rect 16324 13804 16436 13860
rect 16604 13804 16772 13860
rect 17388 13858 17444 14364
rect 18060 14306 18116 14318
rect 18060 14254 18062 14306
rect 18114 14254 18116 14306
rect 17388 13806 17390 13858
rect 17442 13806 17444 13858
rect 16268 13794 16324 13804
rect 16044 13234 16100 13244
rect 16156 13748 16212 13758
rect 16156 12964 16212 13692
rect 16380 13076 16436 13086
rect 16380 12982 16436 13020
rect 15708 12962 15820 12964
rect 15708 12910 15710 12962
rect 15762 12910 15820 12962
rect 15708 12908 15820 12910
rect 15708 12898 15764 12908
rect 15820 12870 15876 12908
rect 16044 12908 16212 12964
rect 15932 12852 15988 12862
rect 15932 12758 15988 12796
rect 15932 12516 15988 12526
rect 15932 12402 15988 12460
rect 15932 12350 15934 12402
rect 15986 12350 15988 12402
rect 15932 12338 15988 12350
rect 16044 12292 16100 12908
rect 16492 12852 16548 12862
rect 16604 12852 16660 13804
rect 17388 13794 17444 13806
rect 17836 13860 17892 13870
rect 18060 13860 18116 14254
rect 17836 13858 18116 13860
rect 17836 13806 17838 13858
rect 17890 13806 18116 13858
rect 17836 13804 18116 13806
rect 17612 13748 17668 13758
rect 17612 13654 17668 13692
rect 17500 13636 17556 13646
rect 17500 13542 17556 13580
rect 17836 13524 17892 13804
rect 17836 13458 17892 13468
rect 16940 12964 16996 12974
rect 16940 12870 16996 12908
rect 17388 12964 17444 12974
rect 17388 12870 17444 12908
rect 17836 12962 17892 12974
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 16548 12796 16660 12852
rect 17724 12850 17780 12862
rect 17724 12798 17726 12850
rect 17778 12798 17780 12850
rect 16492 12758 16548 12796
rect 16156 12740 16212 12750
rect 16156 12646 16212 12684
rect 16268 12740 16324 12750
rect 16268 12738 16436 12740
rect 16268 12686 16270 12738
rect 16322 12686 16436 12738
rect 16268 12684 16436 12686
rect 16268 12674 16324 12684
rect 16268 12292 16324 12302
rect 15596 12236 15876 12292
rect 16044 12236 16268 12292
rect 15596 12068 15652 12078
rect 15596 11974 15652 12012
rect 15372 11620 15428 11630
rect 15372 11526 15428 11564
rect 15820 11396 15876 12236
rect 16268 12198 16324 12236
rect 16044 11732 16100 11742
rect 16044 11506 16100 11676
rect 16044 11454 16046 11506
rect 16098 11454 16100 11506
rect 16044 11442 16100 11454
rect 15932 11396 15988 11406
rect 15260 10994 15316 11004
rect 15372 11394 15988 11396
rect 15372 11342 15934 11394
rect 15986 11342 15988 11394
rect 15372 11340 15988 11342
rect 15148 10836 15204 10846
rect 15036 10834 15204 10836
rect 15036 10782 15150 10834
rect 15202 10782 15204 10834
rect 15036 10780 15204 10782
rect 15148 10770 15204 10780
rect 15260 10836 15316 10846
rect 15260 10742 15316 10780
rect 15372 10834 15428 11340
rect 15932 11330 15988 11340
rect 15372 10782 15374 10834
rect 15426 10782 15428 10834
rect 15372 10770 15428 10782
rect 15708 11170 15764 11182
rect 15708 11118 15710 11170
rect 15762 11118 15764 11170
rect 15708 10500 15764 11118
rect 16156 11170 16212 11182
rect 16156 11118 16158 11170
rect 16210 11118 16212 11170
rect 16156 10836 16212 11118
rect 16156 10770 16212 10780
rect 15820 10500 15876 10510
rect 15708 10498 15876 10500
rect 15708 10446 15822 10498
rect 15874 10446 15876 10498
rect 15708 10444 15876 10446
rect 15820 10388 15876 10444
rect 15820 10322 15876 10332
rect 16268 10052 16324 10062
rect 15484 9714 15540 9726
rect 15484 9662 15486 9714
rect 15538 9662 15540 9714
rect 14924 9550 14926 9602
rect 14978 9550 14980 9602
rect 14924 9492 14980 9550
rect 15260 9604 15316 9614
rect 15260 9510 15316 9548
rect 15372 9602 15428 9614
rect 15372 9550 15374 9602
rect 15426 9550 15428 9602
rect 14924 9156 14980 9436
rect 15036 9156 15092 9166
rect 15372 9156 15428 9550
rect 14924 9154 15092 9156
rect 14924 9102 15038 9154
rect 15090 9102 15092 9154
rect 14924 9100 15092 9102
rect 14588 8194 14644 8204
rect 14028 8034 14084 8046
rect 14028 7982 14030 8034
rect 14082 7982 14084 8034
rect 14028 7812 14084 7982
rect 14028 7746 14084 7756
rect 13916 7476 13972 7486
rect 13916 7382 13972 7420
rect 14588 7362 14644 7374
rect 14588 7310 14590 7362
rect 14642 7310 14644 7362
rect 14588 6804 14644 7310
rect 14924 7140 14980 9100
rect 15036 9090 15092 9100
rect 15148 9100 15428 9156
rect 15484 9156 15540 9662
rect 16044 9602 16100 9614
rect 16044 9550 16046 9602
rect 16098 9550 16100 9602
rect 16044 9492 16100 9550
rect 16044 9426 16100 9436
rect 16268 9268 16324 9996
rect 16380 9268 16436 12684
rect 16716 12738 16772 12750
rect 16716 12686 16718 12738
rect 16770 12686 16772 12738
rect 16492 12516 16548 12526
rect 16716 12516 16772 12686
rect 16548 12460 16772 12516
rect 16492 12450 16548 12460
rect 16716 10052 16772 12460
rect 17612 12738 17668 12750
rect 17612 12686 17614 12738
rect 17666 12686 17668 12738
rect 17612 12290 17668 12686
rect 17724 12628 17780 12798
rect 17836 12852 17892 12910
rect 17836 12786 17892 12796
rect 17724 12572 18116 12628
rect 17724 12404 17780 12414
rect 17724 12310 17780 12348
rect 17612 12238 17614 12290
rect 17666 12238 17668 12290
rect 17612 12226 17668 12238
rect 17948 12178 18004 12190
rect 17948 12126 17950 12178
rect 18002 12126 18004 12178
rect 17948 12068 18004 12126
rect 17948 12002 18004 12012
rect 17612 11506 17668 11518
rect 17612 11454 17614 11506
rect 17666 11454 17668 11506
rect 16716 9996 17220 10052
rect 16604 9714 16660 9726
rect 16604 9662 16606 9714
rect 16658 9662 16660 9714
rect 16604 9604 16660 9662
rect 17164 9714 17220 9996
rect 17164 9662 17166 9714
rect 17218 9662 17220 9714
rect 16380 9212 16548 9268
rect 16268 9202 16324 9212
rect 15484 9100 15988 9156
rect 15148 7588 15204 9100
rect 15372 8932 15428 8942
rect 15372 8838 15428 8876
rect 15484 8818 15540 8830
rect 15484 8766 15486 8818
rect 15538 8766 15540 8818
rect 15484 8372 15540 8766
rect 15484 8306 15540 8316
rect 15260 8148 15316 8158
rect 15260 8054 15316 8092
rect 15596 8036 15652 8046
rect 15596 8034 15764 8036
rect 15596 7982 15598 8034
rect 15650 7982 15764 8034
rect 15596 7980 15764 7982
rect 15596 7970 15652 7980
rect 15596 7588 15652 7598
rect 14924 7074 14980 7084
rect 15036 7532 15204 7588
rect 15260 7586 15652 7588
rect 15260 7534 15598 7586
rect 15650 7534 15652 7586
rect 15260 7532 15652 7534
rect 14588 6738 14644 6748
rect 13916 6690 13972 6702
rect 13916 6638 13918 6690
rect 13970 6638 13972 6690
rect 13916 5794 13972 6638
rect 14140 6692 14196 6702
rect 14140 6578 14196 6636
rect 14140 6526 14142 6578
rect 14194 6526 14196 6578
rect 14140 6514 14196 6526
rect 14476 6580 14532 6590
rect 14476 6486 14532 6524
rect 15036 6580 15092 7532
rect 15148 6916 15204 6926
rect 15260 6916 15316 7532
rect 15596 7522 15652 7532
rect 15708 7252 15764 7980
rect 15932 7364 15988 9100
rect 16156 9044 16212 9054
rect 16044 9042 16212 9044
rect 16044 8990 16158 9042
rect 16210 8990 16212 9042
rect 16044 8988 16212 8990
rect 16044 8372 16100 8988
rect 16156 8978 16212 8988
rect 16492 8932 16548 9212
rect 16268 8930 16548 8932
rect 16268 8878 16494 8930
rect 16546 8878 16548 8930
rect 16268 8876 16548 8878
rect 16156 8484 16212 8494
rect 16268 8484 16324 8876
rect 16492 8866 16548 8876
rect 16156 8482 16324 8484
rect 16156 8430 16158 8482
rect 16210 8430 16324 8482
rect 16156 8428 16324 8430
rect 16492 8484 16548 8494
rect 16156 8418 16212 8428
rect 16492 8390 16548 8428
rect 16044 8306 16100 8316
rect 16380 8372 16436 8382
rect 16380 8146 16436 8316
rect 16380 8094 16382 8146
rect 16434 8094 16436 8146
rect 16380 8082 16436 8094
rect 16492 8036 16548 8046
rect 16380 7700 16436 7710
rect 16492 7700 16548 7980
rect 16436 7644 16548 7700
rect 16380 7606 16436 7644
rect 16044 7364 16100 7374
rect 15932 7308 16044 7364
rect 16044 7298 16100 7308
rect 15820 7252 15876 7262
rect 15708 7196 15820 7252
rect 15820 7186 15876 7196
rect 15148 6914 15316 6916
rect 15148 6862 15150 6914
rect 15202 6862 15316 6914
rect 15148 6860 15316 6862
rect 15372 7140 15428 7150
rect 15148 6850 15204 6860
rect 15260 6692 15316 6702
rect 15372 6692 15428 7084
rect 15260 6690 15428 6692
rect 15260 6638 15262 6690
rect 15314 6638 15428 6690
rect 15260 6636 15428 6638
rect 15484 6916 15540 6926
rect 15260 6626 15316 6636
rect 15036 6514 15092 6524
rect 15148 6356 15204 6366
rect 15036 6020 15092 6030
rect 15036 5926 15092 5964
rect 14812 5906 14868 5918
rect 14812 5854 14814 5906
rect 14866 5854 14868 5906
rect 13916 5742 13918 5794
rect 13970 5742 13972 5794
rect 13916 5730 13972 5742
rect 14364 5796 14420 5806
rect 14364 5702 14420 5740
rect 14812 5236 14868 5854
rect 14812 5170 14868 5180
rect 15148 5234 15204 6300
rect 15484 6020 15540 6860
rect 15596 6804 15652 6814
rect 16156 6804 16212 6814
rect 15596 6802 16212 6804
rect 15596 6750 15598 6802
rect 15650 6750 16158 6802
rect 16210 6750 16212 6802
rect 15596 6748 16212 6750
rect 15596 6738 15652 6748
rect 16156 6738 16212 6748
rect 15484 5964 15652 6020
rect 15148 5182 15150 5234
rect 15202 5182 15204 5234
rect 15148 5170 15204 5182
rect 15372 5794 15428 5806
rect 15372 5742 15374 5794
rect 15426 5742 15428 5794
rect 14364 5124 14420 5134
rect 13244 4172 13860 4228
rect 14140 5010 14196 5022
rect 14140 4958 14142 5010
rect 14194 4958 14196 5010
rect 13244 3668 13300 4172
rect 14140 3780 14196 4958
rect 14140 3714 14196 3724
rect 12460 3444 12516 3482
rect 9660 3332 9940 3388
rect 10444 3332 10612 3388
rect 10668 3378 10724 3388
rect 11900 3332 12180 3388
rect 12460 3378 12516 3388
rect 7756 2930 7812 2940
rect 9884 800 9940 3332
rect 10556 1092 10612 3332
rect 10556 1036 11060 1092
rect 11004 800 11060 1036
rect 12124 800 12180 3332
rect 13244 800 13300 3612
rect 13468 3668 13524 3678
rect 13468 3666 13748 3668
rect 13468 3614 13470 3666
rect 13522 3614 13748 3666
rect 13468 3612 13748 3614
rect 13468 3602 13524 3612
rect 13692 3556 13748 3612
rect 14364 3556 14420 5068
rect 14476 4450 14532 4462
rect 14476 4398 14478 4450
rect 14530 4398 14532 4450
rect 14476 4004 14532 4398
rect 14476 3938 14532 3948
rect 15372 3892 15428 5742
rect 15484 5796 15540 5806
rect 15484 5122 15540 5740
rect 15596 5572 15652 5964
rect 15596 5506 15652 5516
rect 16380 6018 16436 6030
rect 16380 5966 16382 6018
rect 16434 5966 16436 6018
rect 16268 5460 16324 5470
rect 16268 5234 16324 5404
rect 16268 5182 16270 5234
rect 16322 5182 16324 5234
rect 16268 5170 16324 5182
rect 15484 5070 15486 5122
rect 15538 5070 15540 5122
rect 15484 5058 15540 5070
rect 16380 5124 16436 5966
rect 16380 5058 16436 5068
rect 16604 4226 16660 9548
rect 16716 9602 16772 9614
rect 16716 9550 16718 9602
rect 16770 9550 16772 9602
rect 16716 9156 16772 9550
rect 16940 9604 16996 9614
rect 16940 9602 17108 9604
rect 16940 9550 16942 9602
rect 16994 9550 17108 9602
rect 16940 9548 17108 9550
rect 16940 9538 16996 9548
rect 16716 9100 16996 9156
rect 16828 8932 16884 8942
rect 16828 8838 16884 8876
rect 16716 7700 16772 7710
rect 16716 7140 16772 7644
rect 16716 7074 16772 7084
rect 16940 6132 16996 9100
rect 17052 7924 17108 9548
rect 17164 9268 17220 9662
rect 17500 9716 17556 9726
rect 17500 9622 17556 9660
rect 17612 9492 17668 11454
rect 18060 11508 18116 12572
rect 17836 11396 17892 11406
rect 17836 11302 17892 11340
rect 18060 10834 18116 11452
rect 18060 10782 18062 10834
rect 18114 10782 18116 10834
rect 18060 10770 18116 10782
rect 17836 10610 17892 10622
rect 17836 10558 17838 10610
rect 17890 10558 17892 10610
rect 17836 9716 17892 10558
rect 18172 10052 18228 15092
rect 18508 15092 18676 15148
rect 18732 15932 18956 15988
rect 18508 12402 18564 15092
rect 18732 14418 18788 15932
rect 18956 15894 19012 15932
rect 19068 15148 19124 16828
rect 19292 16882 19348 16894
rect 19292 16830 19294 16882
rect 19346 16830 19348 16882
rect 19180 16770 19236 16782
rect 19180 16718 19182 16770
rect 19234 16718 19236 16770
rect 19180 16100 19236 16718
rect 19292 16772 19348 16830
rect 19292 16706 19348 16716
rect 19516 16436 19572 16446
rect 19404 16100 19460 16110
rect 19180 16098 19460 16100
rect 19180 16046 19406 16098
rect 19458 16046 19460 16098
rect 19180 16044 19460 16046
rect 19404 16034 19460 16044
rect 18732 14366 18734 14418
rect 18786 14366 18788 14418
rect 18620 14306 18676 14318
rect 18620 14254 18622 14306
rect 18674 14254 18676 14306
rect 18620 12628 18676 14254
rect 18620 12562 18676 12572
rect 18508 12350 18510 12402
rect 18562 12350 18564 12402
rect 18508 12338 18564 12350
rect 18620 12290 18676 12302
rect 18620 12238 18622 12290
rect 18674 12238 18676 12290
rect 18620 12068 18676 12238
rect 18396 11954 18452 11966
rect 18396 11902 18398 11954
rect 18450 11902 18452 11954
rect 18396 11506 18452 11902
rect 18396 11454 18398 11506
rect 18450 11454 18452 11506
rect 18396 11442 18452 11454
rect 18172 9986 18228 9996
rect 17836 9650 17892 9660
rect 18396 9714 18452 9726
rect 18396 9662 18398 9714
rect 18450 9662 18452 9714
rect 17164 9202 17220 9212
rect 17500 9436 17668 9492
rect 18060 9602 18116 9614
rect 18284 9604 18340 9614
rect 18060 9550 18062 9602
rect 18114 9550 18116 9602
rect 17276 9044 17332 9054
rect 17276 8484 17332 8988
rect 17500 8930 17556 9436
rect 18060 9380 18116 9550
rect 18172 9602 18340 9604
rect 18172 9550 18286 9602
rect 18338 9550 18340 9602
rect 18172 9548 18340 9550
rect 18172 9492 18228 9548
rect 18284 9538 18340 9548
rect 18172 9426 18228 9436
rect 17724 9324 18116 9380
rect 18284 9380 18340 9390
rect 17612 9268 17668 9278
rect 17612 9174 17668 9212
rect 17724 9044 17780 9324
rect 17500 8878 17502 8930
rect 17554 8878 17556 8930
rect 17500 8866 17556 8878
rect 17612 8988 17780 9044
rect 17836 9154 17892 9166
rect 17836 9102 17838 9154
rect 17890 9102 17892 9154
rect 17836 9044 17892 9102
rect 18172 9154 18228 9166
rect 18172 9102 18174 9154
rect 18226 9102 18228 9154
rect 18172 9044 18228 9102
rect 17836 8988 18228 9044
rect 17276 8418 17332 8428
rect 17388 8372 17444 8382
rect 17612 8372 17668 8988
rect 17388 8370 17668 8372
rect 17388 8318 17390 8370
rect 17442 8318 17668 8370
rect 17388 8316 17668 8318
rect 17388 8306 17444 8316
rect 17052 7858 17108 7868
rect 17724 8260 17780 8270
rect 17836 8260 17892 8988
rect 17724 8258 17892 8260
rect 17724 8206 17726 8258
rect 17778 8206 17892 8258
rect 17724 8204 17892 8206
rect 17948 8820 18004 8830
rect 17724 7588 17780 8204
rect 17724 7522 17780 7532
rect 17948 7586 18004 8764
rect 18284 8820 18340 9324
rect 18396 9044 18452 9662
rect 18620 9268 18676 12012
rect 18732 11396 18788 14366
rect 18956 15092 19124 15148
rect 19292 15874 19348 15886
rect 19292 15822 19294 15874
rect 19346 15822 19348 15874
rect 18956 14308 19012 15092
rect 18732 11330 18788 11340
rect 18844 14306 19012 14308
rect 18844 14254 18958 14306
rect 19010 14254 19012 14306
rect 18844 14252 19012 14254
rect 18844 11172 18900 14252
rect 18956 14242 19012 14252
rect 19180 14306 19236 14318
rect 19180 14254 19182 14306
rect 19234 14254 19236 14306
rect 19180 13972 19236 14254
rect 19180 13906 19236 13916
rect 19068 13858 19124 13870
rect 19068 13806 19070 13858
rect 19122 13806 19124 13858
rect 19068 13524 19124 13806
rect 19068 13458 19124 13468
rect 19180 11620 19236 11630
rect 19292 11620 19348 15822
rect 19516 15540 19572 16380
rect 19628 15988 19684 17276
rect 19836 17276 20100 17286
rect 20188 17276 20580 17332
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 19852 17014 19908 17052
rect 20188 16994 20244 17006
rect 20188 16942 20190 16994
rect 20242 16942 20244 16994
rect 20076 16772 20132 16782
rect 20076 16678 20132 16716
rect 19628 15922 19684 15932
rect 20188 15876 20244 16942
rect 20412 16882 20468 16894
rect 20412 16830 20414 16882
rect 20466 16830 20468 16882
rect 20412 16100 20468 16830
rect 20524 16884 20580 17276
rect 20972 16994 21028 17006
rect 20972 16942 20974 16994
rect 21026 16942 21028 16994
rect 20748 16884 20804 16894
rect 20524 16882 20804 16884
rect 20524 16830 20750 16882
rect 20802 16830 20804 16882
rect 20524 16828 20804 16830
rect 20748 16772 20804 16828
rect 20860 16772 20916 16782
rect 20748 16716 20860 16772
rect 20860 16706 20916 16716
rect 20412 16034 20468 16044
rect 20636 16660 20692 16670
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19516 15474 19572 15484
rect 20076 15540 20132 15550
rect 20188 15540 20244 15820
rect 20412 15876 20468 15886
rect 20636 15876 20692 16604
rect 20972 16100 21028 16942
rect 21308 16996 21364 17006
rect 21308 16902 21364 16940
rect 21420 16436 21476 19182
rect 21980 19234 22036 19852
rect 22764 19796 22820 20524
rect 22988 20580 23044 20748
rect 23324 20692 23380 23548
rect 24220 22596 24276 23884
rect 24668 23716 24724 23726
rect 23436 22484 23492 22494
rect 23436 22390 23492 22428
rect 24220 22482 24276 22540
rect 24220 22430 24222 22482
rect 24274 22430 24276 22482
rect 24220 22418 24276 22430
rect 24332 23604 24388 23614
rect 23436 22036 23492 22046
rect 23436 21810 23492 21980
rect 23436 21758 23438 21810
rect 23490 21758 23492 21810
rect 23436 21746 23492 21758
rect 23772 21700 23828 21710
rect 23772 21606 23828 21644
rect 24332 21586 24388 23548
rect 24668 21700 24724 23660
rect 25228 22820 25284 22830
rect 25228 22484 25284 22764
rect 24780 22482 25284 22484
rect 24780 22430 25230 22482
rect 25282 22430 25284 22482
rect 24780 22428 25284 22430
rect 24780 22370 24836 22428
rect 25228 22418 25284 22428
rect 24780 22318 24782 22370
rect 24834 22318 24836 22370
rect 24780 22306 24836 22318
rect 24668 21634 24724 21644
rect 24332 21534 24334 21586
rect 24386 21534 24388 21586
rect 24332 21522 24388 21534
rect 25340 21026 25396 25228
rect 25452 25218 25508 25228
rect 25788 22146 25844 22158
rect 25788 22094 25790 22146
rect 25842 22094 25844 22146
rect 25788 21812 25844 22094
rect 25564 21756 25844 21812
rect 25452 21700 25508 21710
rect 25452 21606 25508 21644
rect 25564 21252 25620 21756
rect 25788 21588 25844 21598
rect 25340 20974 25342 21026
rect 25394 20974 25396 21026
rect 25340 20962 25396 20974
rect 25452 21196 25620 21252
rect 25676 21586 25844 21588
rect 25676 21534 25790 21586
rect 25842 21534 25844 21586
rect 25676 21532 25844 21534
rect 23996 20916 24052 20926
rect 23996 20914 24276 20916
rect 23996 20862 23998 20914
rect 24050 20862 24276 20914
rect 23996 20860 24276 20862
rect 23996 20850 24052 20860
rect 23436 20692 23492 20702
rect 23324 20690 23492 20692
rect 23324 20638 23438 20690
rect 23490 20638 23492 20690
rect 23324 20636 23492 20638
rect 22988 20514 23044 20524
rect 23436 20468 23492 20636
rect 23436 20402 23492 20412
rect 23660 20580 23716 20590
rect 23436 20020 23492 20030
rect 23436 19926 23492 19964
rect 22652 19740 22820 19796
rect 21980 19182 21982 19234
rect 22034 19182 22036 19234
rect 21980 19170 22036 19182
rect 22428 19234 22484 19246
rect 22428 19182 22430 19234
rect 22482 19182 22484 19234
rect 21868 19124 21924 19134
rect 21868 18788 21924 19068
rect 21868 18732 22036 18788
rect 21756 18452 21812 18462
rect 21532 17668 21588 17678
rect 21532 17574 21588 17612
rect 21756 17554 21812 18396
rect 21756 17502 21758 17554
rect 21810 17502 21812 17554
rect 21756 17490 21812 17502
rect 21868 17556 21924 17566
rect 21868 17462 21924 17500
rect 21980 17332 22036 18732
rect 22092 18340 22148 18350
rect 22428 18340 22484 19182
rect 22092 18338 22596 18340
rect 22092 18286 22094 18338
rect 22146 18286 22596 18338
rect 22092 18284 22596 18286
rect 22092 18004 22148 18284
rect 22092 17938 22148 17948
rect 22092 17556 22148 17566
rect 22092 17462 22148 17500
rect 22204 17442 22260 17454
rect 22428 17444 22484 17454
rect 22204 17390 22206 17442
rect 22258 17390 22260 17442
rect 21980 17276 22148 17332
rect 21756 16994 21812 17006
rect 21756 16942 21758 16994
rect 21810 16942 21812 16994
rect 21756 16884 21812 16942
rect 21756 16818 21812 16828
rect 21980 16996 22036 17006
rect 21644 16772 21700 16782
rect 21644 16678 21700 16716
rect 21980 16770 22036 16940
rect 21980 16718 21982 16770
rect 22034 16718 22036 16770
rect 21980 16706 22036 16718
rect 21420 16370 21476 16380
rect 20412 15874 20692 15876
rect 20412 15822 20414 15874
rect 20466 15822 20692 15874
rect 20412 15820 20692 15822
rect 20412 15810 20468 15820
rect 20076 15538 20244 15540
rect 20076 15486 20078 15538
rect 20130 15486 20244 15538
rect 20076 15484 20244 15486
rect 20076 15474 20132 15484
rect 20412 15426 20468 15438
rect 20412 15374 20414 15426
rect 20466 15374 20468 15426
rect 19628 15314 19684 15326
rect 19628 15262 19630 15314
rect 19682 15262 19684 15314
rect 19628 14756 19684 15262
rect 19852 15314 19908 15326
rect 19852 15262 19854 15314
rect 19906 15262 19908 15314
rect 19740 15204 19796 15242
rect 19740 15138 19796 15148
rect 19740 14756 19796 14766
rect 19404 14754 19796 14756
rect 19404 14702 19742 14754
rect 19794 14702 19796 14754
rect 19404 14700 19796 14702
rect 19404 14530 19460 14700
rect 19740 14690 19796 14700
rect 19852 14756 19908 15262
rect 20412 15148 20468 15374
rect 20636 15314 20692 15820
rect 20748 16044 21028 16100
rect 21756 16100 21812 16110
rect 20748 15652 20804 16044
rect 20860 15876 20916 15886
rect 20860 15874 21364 15876
rect 20860 15822 20862 15874
rect 20914 15822 21364 15874
rect 20860 15820 21364 15822
rect 20860 15810 20916 15820
rect 20748 15596 21028 15652
rect 20636 15262 20638 15314
rect 20690 15262 20692 15314
rect 20636 15250 20692 15262
rect 20300 15092 20468 15148
rect 20972 15204 21028 15596
rect 19852 14690 19908 14700
rect 20076 14868 20132 14878
rect 19404 14478 19406 14530
rect 19458 14478 19460 14530
rect 19404 14466 19460 14478
rect 20076 14530 20132 14812
rect 20076 14478 20078 14530
rect 20130 14478 20132 14530
rect 20076 14420 20132 14478
rect 20300 14532 20356 15092
rect 20300 14466 20356 14476
rect 20636 14756 20692 14766
rect 19516 14364 20132 14420
rect 19516 13746 19572 14364
rect 20188 14308 20244 14318
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19516 13694 19518 13746
rect 19570 13694 19572 13746
rect 19516 13682 19572 13694
rect 20076 13748 20132 13758
rect 20188 13748 20244 14252
rect 20636 13972 20692 14700
rect 20860 14644 20916 14654
rect 20524 13916 20692 13972
rect 20748 14418 20804 14430
rect 20748 14366 20750 14418
rect 20802 14366 20804 14418
rect 20524 13858 20580 13916
rect 20524 13806 20526 13858
rect 20578 13806 20580 13858
rect 20524 13794 20580 13806
rect 20748 13748 20804 14366
rect 20076 13746 20356 13748
rect 20076 13694 20078 13746
rect 20130 13694 20356 13746
rect 20076 13692 20356 13694
rect 20076 13682 20132 13692
rect 19628 13634 19684 13646
rect 19628 13582 19630 13634
rect 19682 13582 19684 13634
rect 19180 11618 19460 11620
rect 19180 11566 19182 11618
rect 19234 11566 19460 11618
rect 19180 11564 19460 11566
rect 19180 11554 19236 11564
rect 18620 9202 18676 9212
rect 18732 11116 18900 11172
rect 18956 11508 19012 11518
rect 18956 11172 19012 11452
rect 18396 8978 18452 8988
rect 18508 9044 18564 9054
rect 18732 9044 18788 11116
rect 18956 11106 19012 11116
rect 19068 11396 19124 11406
rect 18956 10836 19012 10846
rect 18956 10742 19012 10780
rect 19068 10834 19124 11340
rect 19068 10782 19070 10834
rect 19122 10782 19124 10834
rect 19068 10770 19124 10782
rect 19068 10612 19124 10622
rect 18844 9940 18900 9950
rect 18844 9602 18900 9884
rect 18844 9550 18846 9602
rect 18898 9550 18900 9602
rect 18844 9380 18900 9550
rect 18844 9314 18900 9324
rect 19068 9266 19124 10556
rect 19292 10610 19348 10622
rect 19292 10558 19294 10610
rect 19346 10558 19348 10610
rect 19068 9214 19070 9266
rect 19122 9214 19124 9266
rect 19068 9202 19124 9214
rect 19180 10052 19236 10062
rect 19180 9268 19236 9996
rect 19292 9940 19348 10558
rect 19404 10388 19460 11564
rect 19516 11170 19572 11182
rect 19516 11118 19518 11170
rect 19570 11118 19572 11170
rect 19516 10612 19572 11118
rect 19516 10546 19572 10556
rect 19628 10610 19684 13582
rect 20188 13524 20244 13534
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10948 20244 13468
rect 20300 12516 20356 13692
rect 20748 13682 20804 13692
rect 20300 12460 20580 12516
rect 20300 11956 20356 11966
rect 20300 11394 20356 11900
rect 20300 11342 20302 11394
rect 20354 11342 20356 11394
rect 20300 11330 20356 11342
rect 20524 11394 20580 12460
rect 20860 12178 20916 14588
rect 20860 12126 20862 12178
rect 20914 12126 20916 12178
rect 20748 11956 20804 11966
rect 20860 11956 20916 12126
rect 20804 11900 20916 11956
rect 20748 11890 20804 11900
rect 20860 11396 20916 11406
rect 20524 11342 20526 11394
rect 20578 11342 20580 11394
rect 20524 11330 20580 11342
rect 20636 11394 20916 11396
rect 20636 11342 20862 11394
rect 20914 11342 20916 11394
rect 20636 11340 20916 11342
rect 20188 10882 20244 10892
rect 19964 10722 20020 10734
rect 19964 10670 19966 10722
rect 20018 10670 20020 10722
rect 19628 10558 19630 10610
rect 19682 10558 19684 10610
rect 19628 10546 19684 10558
rect 19740 10612 19796 10622
rect 19740 10518 19796 10556
rect 19964 10388 20020 10670
rect 20076 10724 20132 10734
rect 20412 10724 20468 10734
rect 20636 10724 20692 11340
rect 20860 11330 20916 11340
rect 20748 11172 20804 11182
rect 20972 11172 21028 15148
rect 21196 15540 21252 15550
rect 21196 14754 21252 15484
rect 21308 15148 21364 15820
rect 21644 15874 21700 15886
rect 21644 15822 21646 15874
rect 21698 15822 21700 15874
rect 21420 15428 21476 15438
rect 21420 15334 21476 15372
rect 21532 15204 21588 15214
rect 21308 15092 21476 15148
rect 21196 14702 21198 14754
rect 21250 14702 21252 14754
rect 21196 14690 21252 14702
rect 21308 14532 21364 14542
rect 21308 14418 21364 14476
rect 21308 14366 21310 14418
rect 21362 14366 21364 14418
rect 21308 14354 21364 14366
rect 21084 14308 21140 14318
rect 21084 12628 21140 14252
rect 21420 14308 21476 15092
rect 21532 14530 21588 15148
rect 21532 14478 21534 14530
rect 21586 14478 21588 14530
rect 21532 14466 21588 14478
rect 21644 14308 21700 15822
rect 21756 15204 21812 16044
rect 21980 15876 22036 15886
rect 21980 15316 22036 15820
rect 21980 15222 22036 15260
rect 21868 15204 21924 15214
rect 21756 15202 21924 15204
rect 21756 15150 21870 15202
rect 21922 15150 21924 15202
rect 21756 15148 21924 15150
rect 22092 15148 22148 17276
rect 22204 16772 22260 17390
rect 22204 15540 22260 16716
rect 22316 17442 22484 17444
rect 22316 17390 22430 17442
rect 22482 17390 22484 17442
rect 22316 17388 22484 17390
rect 22316 15986 22372 17388
rect 22428 17378 22484 17388
rect 22540 17220 22596 18284
rect 22540 17154 22596 17164
rect 22428 16884 22484 16894
rect 22428 16790 22484 16828
rect 22428 16436 22484 16446
rect 22428 16098 22484 16380
rect 22428 16046 22430 16098
rect 22482 16046 22484 16098
rect 22428 16034 22484 16046
rect 22316 15934 22318 15986
rect 22370 15934 22372 15986
rect 22316 15922 22372 15934
rect 22204 15474 22260 15484
rect 21756 14644 21812 15148
rect 21868 15138 21924 15148
rect 21756 14578 21812 14588
rect 21980 15092 22148 15148
rect 22204 15314 22260 15326
rect 22204 15262 22206 15314
rect 22258 15262 22260 15314
rect 22204 15204 22260 15262
rect 22204 15138 22260 15148
rect 22316 15316 22372 15326
rect 22316 15148 22372 15260
rect 22316 15092 22484 15148
rect 21420 14252 21700 14308
rect 21756 14418 21812 14430
rect 21756 14366 21758 14418
rect 21810 14366 21812 14418
rect 21420 14196 21476 14252
rect 21196 14140 21476 14196
rect 21196 13858 21252 14140
rect 21308 13972 21364 13982
rect 21756 13972 21812 14366
rect 21364 13916 21812 13972
rect 21308 13878 21364 13916
rect 21196 13806 21198 13858
rect 21250 13806 21252 13858
rect 21196 13076 21252 13806
rect 21420 13748 21476 13758
rect 21420 13654 21476 13692
rect 21868 13748 21924 13758
rect 21980 13748 22036 15092
rect 22428 14530 22484 15092
rect 22428 14478 22430 14530
rect 22482 14478 22484 14530
rect 22428 14466 22484 14478
rect 22540 14644 22596 14654
rect 22652 14644 22708 19740
rect 22988 19122 23044 19134
rect 22988 19070 22990 19122
rect 23042 19070 23044 19122
rect 22988 17892 23044 19070
rect 22988 17826 23044 17836
rect 23660 17778 23716 20524
rect 23884 20132 23940 20142
rect 23772 18338 23828 18350
rect 23772 18286 23774 18338
rect 23826 18286 23828 18338
rect 23772 18004 23828 18286
rect 23772 17938 23828 17948
rect 23660 17726 23662 17778
rect 23714 17726 23716 17778
rect 23660 17714 23716 17726
rect 23212 17666 23268 17678
rect 23212 17614 23214 17666
rect 23266 17614 23268 17666
rect 22876 17442 22932 17454
rect 22876 17390 22878 17442
rect 22930 17390 22932 17442
rect 22764 16770 22820 16782
rect 22764 16718 22766 16770
rect 22818 16718 22820 16770
rect 22764 14868 22820 16718
rect 22876 16772 22932 17390
rect 23212 17108 23268 17614
rect 23212 17052 23828 17108
rect 23772 16996 23828 17052
rect 23324 16884 23380 16894
rect 22876 16706 22932 16716
rect 23212 16882 23380 16884
rect 23212 16830 23326 16882
rect 23378 16830 23380 16882
rect 23212 16828 23380 16830
rect 22988 16660 23044 16670
rect 22988 16212 23044 16604
rect 22988 16146 23044 16156
rect 23212 15202 23268 16828
rect 23324 16818 23380 16828
rect 23772 16882 23828 16940
rect 23772 16830 23774 16882
rect 23826 16830 23828 16882
rect 23772 16818 23828 16830
rect 23884 16436 23940 20076
rect 23996 19346 24052 19358
rect 23996 19294 23998 19346
rect 24050 19294 24052 19346
rect 23996 16660 24052 19294
rect 24108 19234 24164 19246
rect 24108 19182 24110 19234
rect 24162 19182 24164 19234
rect 24108 18338 24164 19182
rect 24108 18286 24110 18338
rect 24162 18286 24164 18338
rect 24108 17668 24164 18286
rect 24220 19122 24276 20860
rect 24780 20804 24836 20814
rect 25452 20804 25508 21196
rect 24780 20710 24836 20748
rect 25116 20748 25508 20804
rect 25564 20802 25620 20814
rect 25564 20750 25566 20802
rect 25618 20750 25620 20802
rect 25004 20690 25060 20702
rect 25004 20638 25006 20690
rect 25058 20638 25060 20690
rect 24220 19070 24222 19122
rect 24274 19070 24276 19122
rect 24220 18228 24276 19070
rect 24444 20578 24500 20590
rect 24444 20526 24446 20578
rect 24498 20526 24500 20578
rect 24444 18676 24500 20526
rect 24556 19796 24612 19806
rect 24556 19702 24612 19740
rect 24444 18610 24500 18620
rect 25004 18564 25060 20638
rect 25116 20132 25172 20748
rect 25564 20692 25620 20750
rect 25564 20626 25620 20636
rect 25228 20580 25284 20590
rect 25228 20578 25508 20580
rect 25228 20526 25230 20578
rect 25282 20526 25508 20578
rect 25228 20524 25508 20526
rect 25228 20514 25284 20524
rect 25116 20066 25172 20076
rect 25340 20132 25396 20142
rect 25340 20038 25396 20076
rect 25004 18498 25060 18508
rect 25228 18562 25284 18574
rect 25228 18510 25230 18562
rect 25282 18510 25284 18562
rect 24556 18450 24612 18462
rect 24556 18398 24558 18450
rect 24610 18398 24612 18450
rect 24444 18228 24500 18238
rect 24220 18172 24444 18228
rect 24108 17602 24164 17612
rect 24444 17554 24500 18172
rect 24556 18004 24612 18398
rect 25228 18452 25284 18510
rect 25228 18386 25284 18396
rect 24780 18340 24836 18350
rect 24780 18116 24836 18284
rect 24780 18050 24836 18060
rect 24556 17938 24612 17948
rect 24444 17502 24446 17554
rect 24498 17502 24500 17554
rect 24444 17490 24500 17502
rect 24668 17668 24724 17678
rect 23996 16594 24052 16604
rect 24332 16882 24388 16894
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 23884 16370 23940 16380
rect 23996 16098 24052 16110
rect 23996 16046 23998 16098
rect 24050 16046 24052 16098
rect 23548 15988 23604 15998
rect 23548 15316 23604 15932
rect 23548 15250 23604 15260
rect 23212 15150 23214 15202
rect 23266 15150 23268 15202
rect 23212 15138 23268 15150
rect 23996 15148 24052 16046
rect 23436 15092 24052 15148
rect 23436 15090 23492 15092
rect 23436 15038 23438 15090
rect 23490 15038 23492 15090
rect 23436 15026 23492 15038
rect 22764 14812 23156 14868
rect 23100 14644 23156 14812
rect 23212 14644 23268 14654
rect 22652 14588 22932 14644
rect 23100 14588 23212 14644
rect 22540 14420 22596 14588
rect 22764 14420 22820 14430
rect 22540 14418 22820 14420
rect 22540 14366 22766 14418
rect 22818 14366 22820 14418
rect 22540 14364 22820 14366
rect 22764 14354 22820 14364
rect 22092 14308 22148 14318
rect 22092 14214 22148 14252
rect 22876 14196 22932 14588
rect 23212 14578 23268 14588
rect 21868 13746 22036 13748
rect 21868 13694 21870 13746
rect 21922 13694 22036 13746
rect 21868 13692 22036 13694
rect 22764 14140 22932 14196
rect 22988 14530 23044 14542
rect 22988 14478 22990 14530
rect 23042 14478 23044 14530
rect 22988 14420 23044 14478
rect 23548 14532 23604 14542
rect 23548 14438 23604 14476
rect 24332 14530 24388 16830
rect 24668 16884 24724 17612
rect 25228 16996 25284 17006
rect 25452 16996 25508 20524
rect 25564 19124 25620 19134
rect 25564 18676 25620 19068
rect 25564 18582 25620 18620
rect 25676 18452 25732 21532
rect 25788 21522 25844 21532
rect 25900 21364 25956 25678
rect 26012 27636 26068 27646
rect 26012 22932 26068 27580
rect 26124 25506 26180 25518
rect 26124 25454 26126 25506
rect 26178 25454 26180 25506
rect 26124 25284 26180 25454
rect 26124 25218 26180 25228
rect 26236 25396 26292 25406
rect 26236 25060 26292 25340
rect 26012 22866 26068 22876
rect 26124 25004 26292 25060
rect 26348 25172 26404 27806
rect 26572 27860 26628 27870
rect 26572 27858 26740 27860
rect 26572 27806 26574 27858
rect 26626 27806 26740 27858
rect 26572 27804 26740 27806
rect 26572 27794 26628 27804
rect 26572 27300 26628 27310
rect 26572 27206 26628 27244
rect 26684 27186 26740 27804
rect 26684 27134 26686 27186
rect 26738 27134 26740 27186
rect 26684 27122 26740 27134
rect 26796 26964 26852 32284
rect 27020 31778 27076 33404
rect 27132 33394 27188 33404
rect 27020 31726 27022 31778
rect 27074 31726 27076 31778
rect 27020 31714 27076 31726
rect 27132 33234 27188 33246
rect 27132 33182 27134 33234
rect 27186 33182 27188 33234
rect 27132 31218 27188 33182
rect 27132 31166 27134 31218
rect 27186 31166 27188 31218
rect 27132 31154 27188 31166
rect 27020 30210 27076 30222
rect 27020 30158 27022 30210
rect 27074 30158 27076 30210
rect 27020 29876 27076 30158
rect 27020 29810 27076 29820
rect 27244 28532 27300 34524
rect 27356 34356 27412 34750
rect 27580 34580 27636 36430
rect 27692 37380 27748 37390
rect 27692 35924 27748 37324
rect 27804 36482 27860 38110
rect 27916 37828 27972 37838
rect 27916 37380 27972 37772
rect 27916 37314 27972 37324
rect 27804 36430 27806 36482
rect 27858 36430 27860 36482
rect 27804 36418 27860 36430
rect 27916 36372 27972 36382
rect 27916 36278 27972 36316
rect 27692 35812 27748 35868
rect 27804 35812 27860 35822
rect 27692 35810 27860 35812
rect 27692 35758 27806 35810
rect 27858 35758 27860 35810
rect 27692 35756 27860 35758
rect 27804 35364 27860 35756
rect 28028 35308 28084 38612
rect 28140 38612 28308 38668
rect 28700 38946 28756 38958
rect 28700 38894 28702 38946
rect 28754 38894 28756 38946
rect 28700 38724 28756 38894
rect 29036 38948 29092 38958
rect 29036 38668 29092 38892
rect 28700 38658 28756 38668
rect 28140 38050 28196 38612
rect 28140 37998 28142 38050
rect 28194 37998 28196 38050
rect 28140 37986 28196 37998
rect 28476 38610 28532 38622
rect 28476 38558 28478 38610
rect 28530 38558 28532 38610
rect 28252 37154 28308 37166
rect 28252 37102 28254 37154
rect 28306 37102 28308 37154
rect 28252 37044 28308 37102
rect 28252 36978 28308 36988
rect 28364 36932 28420 36942
rect 28140 36482 28196 36494
rect 28140 36430 28142 36482
rect 28194 36430 28196 36482
rect 28140 35922 28196 36430
rect 28140 35870 28142 35922
rect 28194 35870 28196 35922
rect 28140 35858 28196 35870
rect 28364 35810 28420 36876
rect 28364 35758 28366 35810
rect 28418 35758 28420 35810
rect 28364 35746 28420 35758
rect 28140 35698 28196 35710
rect 28140 35646 28142 35698
rect 28194 35646 28196 35698
rect 28140 35476 28196 35646
rect 28140 35410 28196 35420
rect 27804 35298 27860 35308
rect 27916 35252 28084 35308
rect 27804 34690 27860 34702
rect 27804 34638 27806 34690
rect 27858 34638 27860 34690
rect 27580 34524 27748 34580
rect 27356 34300 27636 34356
rect 27580 34242 27636 34300
rect 27580 34190 27582 34242
rect 27634 34190 27636 34242
rect 27580 34178 27636 34190
rect 27468 34130 27524 34142
rect 27468 34078 27470 34130
rect 27522 34078 27524 34130
rect 27468 34020 27524 34078
rect 27692 34020 27748 34524
rect 27804 34244 27860 34638
rect 27804 34178 27860 34188
rect 27468 33964 27748 34020
rect 27804 34020 27860 34030
rect 27468 33124 27524 33964
rect 27804 33926 27860 33964
rect 27580 33124 27636 33134
rect 27468 33122 27636 33124
rect 27468 33070 27582 33122
rect 27634 33070 27636 33122
rect 27468 33068 27636 33070
rect 27580 32340 27636 33068
rect 27916 32676 27972 35252
rect 28252 35140 28308 35150
rect 28028 34914 28084 34926
rect 28028 34862 28030 34914
rect 28082 34862 28084 34914
rect 28028 34356 28084 34862
rect 28028 34290 28084 34300
rect 28140 34914 28196 34926
rect 28140 34862 28142 34914
rect 28194 34862 28196 34914
rect 28028 34132 28084 34142
rect 28028 34038 28084 34076
rect 28140 33572 28196 34862
rect 28252 34914 28308 35084
rect 28252 34862 28254 34914
rect 28306 34862 28308 34914
rect 28252 34850 28308 34862
rect 28476 34692 28532 38558
rect 28924 38612 29092 38668
rect 29372 38668 29428 41020
rect 29596 40404 29652 41132
rect 29596 40338 29652 40348
rect 29372 38612 29652 38668
rect 28700 37268 28756 37278
rect 28700 37154 28756 37212
rect 28924 37266 28980 38612
rect 29484 38388 29540 38398
rect 29372 38332 29484 38388
rect 29260 37268 29316 37278
rect 28924 37214 28926 37266
rect 28978 37214 28980 37266
rect 28924 37202 28980 37214
rect 29036 37266 29316 37268
rect 29036 37214 29262 37266
rect 29314 37214 29316 37266
rect 29036 37212 29316 37214
rect 28700 37102 28702 37154
rect 28754 37102 28756 37154
rect 28588 36260 28644 36270
rect 28588 35476 28644 36204
rect 28700 35476 28756 37102
rect 29036 36820 29092 37212
rect 29260 37202 29316 37212
rect 28924 36260 28980 36270
rect 29036 36260 29092 36764
rect 28980 36204 29092 36260
rect 29148 37042 29204 37054
rect 29148 36990 29150 37042
rect 29202 36990 29204 37042
rect 28924 36194 28980 36204
rect 29148 36036 29204 36990
rect 29372 36596 29428 38332
rect 29484 38322 29540 38332
rect 29484 37378 29540 37390
rect 29484 37326 29486 37378
rect 29538 37326 29540 37378
rect 29484 37268 29540 37326
rect 29484 37202 29540 37212
rect 29148 35970 29204 35980
rect 29260 36540 29428 36596
rect 29260 35924 29316 36540
rect 29596 36484 29652 38612
rect 29708 37826 29764 37838
rect 29708 37774 29710 37826
rect 29762 37774 29764 37826
rect 29708 36820 29764 37774
rect 30044 37266 30100 41804
rect 30156 41636 30212 41646
rect 30156 41186 30212 41580
rect 30156 41134 30158 41186
rect 30210 41134 30212 41186
rect 30156 41122 30212 41134
rect 30492 40404 30548 40414
rect 30268 40290 30324 40302
rect 30268 40238 30270 40290
rect 30322 40238 30324 40290
rect 30268 40180 30324 40238
rect 30268 38948 30324 40124
rect 30492 39730 30548 40348
rect 30492 39678 30494 39730
rect 30546 39678 30548 39730
rect 30492 39666 30548 39678
rect 30604 39060 30660 43708
rect 31164 43764 31220 43774
rect 31276 43764 31332 45054
rect 31612 44548 31668 46398
rect 31612 44482 31668 44492
rect 33404 45108 33460 45118
rect 33404 44996 33460 45052
rect 33516 44996 33572 47180
rect 33740 47012 33796 48076
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35532 47234 35588 47246
rect 35532 47182 35534 47234
rect 35586 47182 35588 47234
rect 35532 47124 35588 47182
rect 35532 47058 35588 47068
rect 33740 46946 33796 46956
rect 35196 46788 35252 46798
rect 34860 46786 35252 46788
rect 34860 46734 35198 46786
rect 35250 46734 35252 46786
rect 34860 46732 35252 46734
rect 34636 46450 34692 46462
rect 34636 46398 34638 46450
rect 34690 46398 34692 46450
rect 34300 45106 34356 45118
rect 34300 45054 34302 45106
rect 34354 45054 34356 45106
rect 33852 44996 33908 45006
rect 34300 44996 34356 45054
rect 33404 44994 34356 44996
rect 33404 44942 33406 44994
rect 33458 44942 33854 44994
rect 33906 44942 34356 44994
rect 33404 44940 34356 44942
rect 31164 43762 31332 43764
rect 31164 43710 31166 43762
rect 31218 43710 31332 43762
rect 31164 43708 31332 43710
rect 31948 44324 32004 44334
rect 31164 43698 31220 43708
rect 31948 43540 32004 44268
rect 32956 43764 33012 43774
rect 32284 43652 32340 43662
rect 32508 43652 32564 43662
rect 32284 43650 32508 43652
rect 32284 43598 32286 43650
rect 32338 43598 32508 43650
rect 32284 43596 32508 43598
rect 32284 43586 32340 43596
rect 32508 43586 32564 43596
rect 32060 43540 32116 43550
rect 31948 43484 32060 43540
rect 32060 43446 32116 43484
rect 31500 43316 31556 43326
rect 31500 43222 31556 43260
rect 31052 42082 31108 42094
rect 31052 42030 31054 42082
rect 31106 42030 31108 42082
rect 30716 41860 30772 41870
rect 30716 41766 30772 41804
rect 31052 41636 31108 42030
rect 31276 41972 31332 41982
rect 31052 41570 31108 41580
rect 31164 41970 31332 41972
rect 31164 41918 31278 41970
rect 31330 41918 31332 41970
rect 31164 41916 31332 41918
rect 31164 41076 31220 41916
rect 31276 41906 31332 41916
rect 32956 41970 33012 43708
rect 33404 43764 33460 44940
rect 33852 44930 33908 44940
rect 34412 44322 34468 44334
rect 34412 44270 34414 44322
rect 34466 44270 34468 44322
rect 34300 44212 34356 44222
rect 33404 43698 33460 43708
rect 33628 44098 33684 44110
rect 34076 44100 34132 44110
rect 33628 44046 33630 44098
rect 33682 44046 33684 44098
rect 33628 43652 33684 44046
rect 33628 43586 33684 43596
rect 33964 44098 34132 44100
rect 33964 44046 34078 44098
rect 34130 44046 34132 44098
rect 33964 44044 34132 44046
rect 33628 41972 33684 41982
rect 32956 41918 32958 41970
rect 33010 41918 33012 41970
rect 30716 41020 31220 41076
rect 31836 41858 31892 41870
rect 31836 41806 31838 41858
rect 31890 41806 31892 41858
rect 30716 40626 30772 41020
rect 31724 40964 31780 40974
rect 30716 40574 30718 40626
rect 30770 40574 30772 40626
rect 30716 40562 30772 40574
rect 31612 40908 31724 40964
rect 31612 40514 31668 40908
rect 31724 40898 31780 40908
rect 31612 40462 31614 40514
rect 31666 40462 31668 40514
rect 31052 40180 31108 40190
rect 31052 40086 31108 40124
rect 30268 38882 30324 38892
rect 30492 39004 30660 39060
rect 30044 37214 30046 37266
rect 30098 37214 30100 37266
rect 30044 37202 30100 37214
rect 29708 36754 29764 36764
rect 29820 37154 29876 37166
rect 29820 37102 29822 37154
rect 29874 37102 29876 37154
rect 29708 36484 29764 36494
rect 29596 36482 29764 36484
rect 29596 36430 29710 36482
rect 29762 36430 29764 36482
rect 29596 36428 29764 36430
rect 29708 36418 29764 36428
rect 29820 36484 29876 37102
rect 29820 36418 29876 36428
rect 29932 37044 29988 37054
rect 30380 37044 30436 37054
rect 29372 36372 29428 36382
rect 29372 36278 29428 36316
rect 29932 36372 29988 36988
rect 29932 36278 29988 36316
rect 30044 37042 30436 37044
rect 30044 36990 30382 37042
rect 30434 36990 30436 37042
rect 30044 36988 30436 36990
rect 30044 36370 30100 36988
rect 30380 36978 30436 36988
rect 30492 36932 30548 39004
rect 30828 38948 30884 38958
rect 30828 38946 31444 38948
rect 30828 38894 30830 38946
rect 30882 38894 31444 38946
rect 30828 38892 31444 38894
rect 30828 38882 30884 38892
rect 30604 38834 30660 38846
rect 30604 38782 30606 38834
rect 30658 38782 30660 38834
rect 30604 38724 30660 38782
rect 31276 38724 31332 38734
rect 30604 38722 31332 38724
rect 30604 38670 31278 38722
rect 31330 38670 31332 38722
rect 30604 38668 31332 38670
rect 31276 38658 31332 38668
rect 30940 38050 30996 38062
rect 30940 37998 30942 38050
rect 30994 37998 30996 38050
rect 30940 37828 30996 37998
rect 31388 38050 31444 38892
rect 31612 38836 31668 40462
rect 31724 40402 31780 40414
rect 31724 40350 31726 40402
rect 31778 40350 31780 40402
rect 31724 40292 31780 40350
rect 31836 40404 31892 41806
rect 32508 40964 32564 40974
rect 32508 40870 32564 40908
rect 31836 40338 31892 40348
rect 32508 40404 32564 40414
rect 32564 40348 32676 40404
rect 32508 40310 32564 40348
rect 31724 40226 31780 40236
rect 31948 40292 32004 40302
rect 31948 38946 32004 40236
rect 31948 38894 31950 38946
rect 32002 38894 32004 38946
rect 31948 38882 32004 38894
rect 32284 38946 32340 38958
rect 32284 38894 32286 38946
rect 32338 38894 32340 38946
rect 31612 38742 31668 38780
rect 31388 37998 31390 38050
rect 31442 37998 31444 38050
rect 31388 37986 31444 37998
rect 32284 38500 32340 38894
rect 30940 37762 30996 37772
rect 30828 37154 30884 37166
rect 30828 37102 30830 37154
rect 30882 37102 30884 37154
rect 30828 37044 30884 37102
rect 30828 36978 30884 36988
rect 31500 37156 31556 37166
rect 30492 36866 30548 36876
rect 30044 36318 30046 36370
rect 30098 36318 30100 36370
rect 30044 36306 30100 36318
rect 30156 36484 30212 36494
rect 29820 36258 29876 36270
rect 29820 36206 29822 36258
rect 29874 36206 29876 36258
rect 29820 36036 29876 36206
rect 30156 36148 30212 36428
rect 30380 36482 30436 36494
rect 30380 36430 30382 36482
rect 30434 36430 30436 36482
rect 30156 36092 30324 36148
rect 29820 35980 30212 36036
rect 29484 35924 29540 35934
rect 29260 35868 29428 35924
rect 29036 35812 29092 35822
rect 29036 35718 29092 35756
rect 29260 35700 29316 35710
rect 29148 35698 29316 35700
rect 29148 35646 29262 35698
rect 29314 35646 29316 35698
rect 29148 35644 29316 35646
rect 29372 35700 29428 35868
rect 29484 35922 29988 35924
rect 29484 35870 29486 35922
rect 29538 35870 29988 35922
rect 29484 35868 29988 35870
rect 29484 35858 29540 35868
rect 29932 35810 29988 35868
rect 29932 35758 29934 35810
rect 29986 35758 29988 35810
rect 29932 35746 29988 35758
rect 29596 35700 29652 35710
rect 29372 35698 29652 35700
rect 29372 35646 29598 35698
rect 29650 35646 29652 35698
rect 29372 35644 29652 35646
rect 29148 35476 29204 35644
rect 29260 35634 29316 35644
rect 29596 35634 29652 35644
rect 30156 35698 30212 35980
rect 30156 35646 30158 35698
rect 30210 35646 30212 35698
rect 30156 35634 30212 35646
rect 30044 35588 30100 35598
rect 29932 35586 30100 35588
rect 29932 35534 30046 35586
rect 30098 35534 30100 35586
rect 29932 35532 30100 35534
rect 28700 35420 29204 35476
rect 29596 35476 29652 35486
rect 28588 35410 28644 35420
rect 28700 35252 28756 35262
rect 28588 35196 28700 35252
rect 28588 34914 28644 35196
rect 28700 35186 28756 35196
rect 28588 34862 28590 34914
rect 28642 34862 28644 34914
rect 28588 34850 28644 34862
rect 29260 35140 29316 35150
rect 28252 34636 28532 34692
rect 28700 34804 28756 34814
rect 28252 33796 28308 34636
rect 28588 34468 28644 34478
rect 28588 34242 28644 34412
rect 28588 34190 28590 34242
rect 28642 34190 28644 34242
rect 28588 34178 28644 34190
rect 28252 33740 28532 33796
rect 28140 33506 28196 33516
rect 28364 33234 28420 33246
rect 28364 33182 28366 33234
rect 28418 33182 28420 33234
rect 28140 33124 28196 33134
rect 28364 33124 28420 33182
rect 28196 33068 28420 33124
rect 28476 33236 28532 33740
rect 28700 33346 28756 34748
rect 29260 34690 29316 35084
rect 29260 34638 29262 34690
rect 29314 34638 29316 34690
rect 29260 34580 29316 34638
rect 29260 34524 29540 34580
rect 28812 34468 28868 34478
rect 28868 34412 29428 34468
rect 28812 34402 28868 34412
rect 28700 33294 28702 33346
rect 28754 33294 28756 33346
rect 28700 33282 28756 33294
rect 28812 34244 28868 34254
rect 28140 33030 28196 33068
rect 27916 32610 27972 32620
rect 27580 32284 28196 32340
rect 27468 31778 27524 31790
rect 27468 31726 27470 31778
rect 27522 31726 27524 31778
rect 27468 31556 27524 31726
rect 27916 31780 27972 31790
rect 27972 31724 28084 31780
rect 27916 31714 27972 31724
rect 27916 31556 27972 31566
rect 27468 31554 27972 31556
rect 27468 31502 27918 31554
rect 27970 31502 27972 31554
rect 27468 31500 27972 31502
rect 27468 30770 27524 30782
rect 27468 30718 27470 30770
rect 27522 30718 27524 30770
rect 27468 29204 27524 30718
rect 27916 30100 27972 31500
rect 28028 30994 28084 31724
rect 28028 30942 28030 30994
rect 28082 30942 28084 30994
rect 28028 30930 28084 30942
rect 27916 30044 28084 30100
rect 27804 29876 27860 29886
rect 27860 29820 27972 29876
rect 27804 29810 27860 29820
rect 27468 28754 27524 29148
rect 27468 28702 27470 28754
rect 27522 28702 27524 28754
rect 27468 28690 27524 28702
rect 27244 28476 27524 28532
rect 27468 28308 27524 28476
rect 27468 28252 27860 28308
rect 27356 28196 27412 28206
rect 27020 28084 27076 28094
rect 27020 27858 27076 28028
rect 27020 27806 27022 27858
rect 27074 27806 27076 27858
rect 27020 27794 27076 27806
rect 27356 27188 27412 28140
rect 27692 27972 27748 27982
rect 27468 27860 27524 27870
rect 27468 27766 27524 27804
rect 26908 27186 27412 27188
rect 26908 27134 27358 27186
rect 27410 27134 27412 27186
rect 26908 27132 27412 27134
rect 26908 27074 26964 27132
rect 27356 27122 27412 27132
rect 27580 27748 27636 27758
rect 26908 27022 26910 27074
rect 26962 27022 26964 27074
rect 26908 27010 26964 27022
rect 26684 26908 26852 26964
rect 27580 26908 27636 27692
rect 26572 25844 26628 25854
rect 26572 25508 26628 25788
rect 26572 25414 26628 25452
rect 25788 21308 25956 21364
rect 26012 21698 26068 21710
rect 26012 21646 26014 21698
rect 26066 21646 26068 21698
rect 25788 19348 25844 21308
rect 25900 21028 25956 21038
rect 25900 20934 25956 20972
rect 25900 20244 25956 20254
rect 26012 20244 26068 21646
rect 26124 21026 26180 25004
rect 26348 24836 26404 25116
rect 26348 24742 26404 24780
rect 26460 24610 26516 24622
rect 26460 24558 26462 24610
rect 26514 24558 26516 24610
rect 26236 24500 26292 24510
rect 26236 23042 26292 24444
rect 26460 24050 26516 24558
rect 26460 23998 26462 24050
rect 26514 23998 26516 24050
rect 26460 23986 26516 23998
rect 26572 23156 26628 23166
rect 26236 22990 26238 23042
rect 26290 22990 26292 23042
rect 26236 22978 26292 22990
rect 26348 23154 26628 23156
rect 26348 23102 26574 23154
rect 26626 23102 26628 23154
rect 26348 23100 26628 23102
rect 26348 21588 26404 23100
rect 26572 23090 26628 23100
rect 26124 20974 26126 21026
rect 26178 20974 26180 21026
rect 26124 20962 26180 20974
rect 26236 21532 26404 21588
rect 26460 22932 26516 22942
rect 26460 21588 26516 22876
rect 26572 22484 26628 22494
rect 26684 22484 26740 26908
rect 27020 26852 27636 26908
rect 26908 25620 26964 25658
rect 26908 25554 26964 25564
rect 27020 25506 27076 26852
rect 27132 25732 27188 25742
rect 27692 25732 27748 27916
rect 27188 25676 27300 25732
rect 27132 25666 27188 25676
rect 27020 25454 27022 25506
rect 27074 25454 27076 25506
rect 27020 25442 27076 25454
rect 27132 25394 27188 25406
rect 27132 25342 27134 25394
rect 27186 25342 27188 25394
rect 26796 25282 26852 25294
rect 26796 25230 26798 25282
rect 26850 25230 26852 25282
rect 26796 25172 26852 25230
rect 26796 25106 26852 25116
rect 27020 25172 27076 25182
rect 26796 24948 26852 24958
rect 26796 24834 26852 24892
rect 26796 24782 26798 24834
rect 26850 24782 26852 24834
rect 26796 24770 26852 24782
rect 26796 24164 26852 24174
rect 26796 24050 26852 24108
rect 26796 23998 26798 24050
rect 26850 23998 26852 24050
rect 26796 23548 26852 23998
rect 27020 23940 27076 25116
rect 27132 24946 27188 25342
rect 27132 24894 27134 24946
rect 27186 24894 27188 24946
rect 27132 24882 27188 24894
rect 27132 24724 27188 24734
rect 27244 24724 27300 25676
rect 27468 25676 27748 25732
rect 27468 25172 27524 25676
rect 27468 25106 27524 25116
rect 27580 25508 27636 25518
rect 27132 24722 27300 24724
rect 27132 24670 27134 24722
rect 27186 24670 27300 24722
rect 27132 24668 27300 24670
rect 27468 24722 27524 24734
rect 27468 24670 27470 24722
rect 27522 24670 27524 24722
rect 27132 24658 27188 24668
rect 27468 24276 27524 24670
rect 27580 24612 27636 25452
rect 27804 25506 27860 28252
rect 27804 25454 27806 25506
rect 27858 25454 27860 25506
rect 27692 25284 27748 25294
rect 27692 25190 27748 25228
rect 27580 24546 27636 24556
rect 27804 24610 27860 25454
rect 27804 24558 27806 24610
rect 27858 24558 27860 24610
rect 27804 24500 27860 24558
rect 27804 24434 27860 24444
rect 27020 23874 27076 23884
rect 27356 24164 27412 24174
rect 27356 23714 27412 24108
rect 27468 23828 27524 24220
rect 27468 23772 27860 23828
rect 27356 23662 27358 23714
rect 27410 23662 27412 23714
rect 26796 23492 26964 23548
rect 26908 23044 26964 23492
rect 27020 23268 27076 23278
rect 27020 23266 27300 23268
rect 27020 23214 27022 23266
rect 27074 23214 27300 23266
rect 27020 23212 27300 23214
rect 27020 23202 27076 23212
rect 26908 22988 27076 23044
rect 26628 22428 26740 22484
rect 26572 22418 26628 22428
rect 26796 21700 26852 21710
rect 26796 21606 26852 21644
rect 26908 21700 26964 21710
rect 26236 21028 26292 21532
rect 26460 21522 26516 21532
rect 26684 21586 26740 21598
rect 26684 21534 26686 21586
rect 26738 21534 26740 21586
rect 26572 21474 26628 21486
rect 26572 21422 26574 21474
rect 26626 21422 26628 21474
rect 26572 21364 26628 21422
rect 25900 20242 26068 20244
rect 25900 20190 25902 20242
rect 25954 20190 26068 20242
rect 25900 20188 26068 20190
rect 26124 20356 26180 20366
rect 25900 20178 25956 20188
rect 25900 20018 25956 20030
rect 25900 19966 25902 20018
rect 25954 19966 25956 20018
rect 25900 19908 25956 19966
rect 26124 19908 26180 20300
rect 26236 20132 26292 20972
rect 26236 20066 26292 20076
rect 26348 21308 26628 21364
rect 26124 19852 26292 19908
rect 25900 19842 25956 19852
rect 26012 19348 26068 19358
rect 25788 19346 26068 19348
rect 25788 19294 26014 19346
rect 26066 19294 26068 19346
rect 25788 19292 26068 19294
rect 26012 19282 26068 19292
rect 25676 18386 25732 18396
rect 25452 16940 25620 16996
rect 25228 16902 25284 16940
rect 24668 16324 24724 16828
rect 25452 16772 25508 16782
rect 24332 14478 24334 14530
rect 24386 14478 24388 14530
rect 21196 13010 21252 13020
rect 21644 13076 21700 13086
rect 21644 12982 21700 13020
rect 21868 12740 21924 13692
rect 22540 13634 22596 13646
rect 22540 13582 22542 13634
rect 22594 13582 22596 13634
rect 22092 12740 22148 12750
rect 21868 12738 22148 12740
rect 21868 12686 22094 12738
rect 22146 12686 22148 12738
rect 21868 12684 22148 12686
rect 21084 12572 21476 12628
rect 21084 12290 21140 12302
rect 21084 12238 21086 12290
rect 21138 12238 21140 12290
rect 21084 11732 21140 12238
rect 21084 11666 21140 11676
rect 21420 12290 21476 12572
rect 21420 12238 21422 12290
rect 21474 12238 21476 12290
rect 21420 11394 21476 12238
rect 21980 12292 22036 12302
rect 21980 12198 22036 12236
rect 21756 12178 21812 12190
rect 21756 12126 21758 12178
rect 21810 12126 21812 12178
rect 21756 11732 21812 12126
rect 21644 11676 21756 11732
rect 21644 11620 21700 11676
rect 21756 11666 21812 11676
rect 21868 12066 21924 12078
rect 21868 12014 21870 12066
rect 21922 12014 21924 12066
rect 21420 11342 21422 11394
rect 21474 11342 21476 11394
rect 21420 11330 21476 11342
rect 21532 11564 21700 11620
rect 21868 11620 21924 12014
rect 22092 12068 22148 12684
rect 22540 12402 22596 13582
rect 22540 12350 22542 12402
rect 22594 12350 22596 12402
rect 22540 12338 22596 12350
rect 22316 12292 22372 12302
rect 22316 12198 22372 12236
rect 22092 12002 22148 12012
rect 22652 12178 22708 12190
rect 22652 12126 22654 12178
rect 22706 12126 22708 12178
rect 22652 11956 22708 12126
rect 22652 11890 22708 11900
rect 21532 11394 21588 11564
rect 21868 11554 21924 11564
rect 21532 11342 21534 11394
rect 21586 11342 21588 11394
rect 21532 11330 21588 11342
rect 22092 11396 22148 11406
rect 22652 11396 22708 11406
rect 22092 11394 22708 11396
rect 22092 11342 22094 11394
rect 22146 11342 22654 11394
rect 22706 11342 22708 11394
rect 22092 11340 22708 11342
rect 22092 11330 22148 11340
rect 21644 11282 21700 11294
rect 21644 11230 21646 11282
rect 21698 11230 21700 11282
rect 20748 11170 21028 11172
rect 20748 11118 20750 11170
rect 20802 11118 21028 11170
rect 20748 11116 21028 11118
rect 20748 11106 20804 11116
rect 20972 11060 21028 11116
rect 20972 10994 21028 11004
rect 21196 11172 21252 11182
rect 21644 11172 21700 11230
rect 21252 11116 21700 11172
rect 20076 10722 20692 10724
rect 20076 10670 20078 10722
rect 20130 10670 20414 10722
rect 20466 10670 20692 10722
rect 20076 10668 20692 10670
rect 20748 10948 20804 10958
rect 20076 10658 20132 10668
rect 20412 10658 20468 10668
rect 20748 10612 20804 10892
rect 21196 10834 21252 11116
rect 21196 10782 21198 10834
rect 21250 10782 21252 10834
rect 21196 10770 21252 10782
rect 22316 11060 22372 11070
rect 22316 10834 22372 11004
rect 22316 10782 22318 10834
rect 22370 10782 22372 10834
rect 22316 10770 22372 10782
rect 22540 10834 22596 11340
rect 22652 11330 22708 11340
rect 22540 10782 22542 10834
rect 22594 10782 22596 10834
rect 22540 10770 22596 10782
rect 19404 10332 20020 10388
rect 19292 9884 19684 9940
rect 19292 9716 19348 9726
rect 19292 9622 19348 9660
rect 19404 9602 19460 9614
rect 19404 9550 19406 9602
rect 19458 9550 19460 9602
rect 19292 9268 19348 9278
rect 19180 9266 19348 9268
rect 19180 9214 19294 9266
rect 19346 9214 19348 9266
rect 19180 9212 19348 9214
rect 19292 9202 19348 9212
rect 19404 9268 19460 9550
rect 19404 9174 19460 9212
rect 18956 9156 19012 9166
rect 18508 9042 18788 9044
rect 18508 8990 18510 9042
rect 18562 8990 18788 9042
rect 18508 8988 18788 8990
rect 18844 9042 18900 9054
rect 18844 8990 18846 9042
rect 18898 8990 18900 9042
rect 18284 8754 18340 8764
rect 18508 8820 18564 8988
rect 18844 8932 18900 8990
rect 18844 8866 18900 8876
rect 18508 8754 18564 8764
rect 18732 8372 18788 8382
rect 18732 8278 18788 8316
rect 18844 8260 18900 8270
rect 18956 8260 19012 9100
rect 19180 9044 19236 9054
rect 19180 8950 19236 8988
rect 18844 8258 19012 8260
rect 18844 8206 18846 8258
rect 18898 8206 19012 8258
rect 18844 8204 19012 8206
rect 19292 8820 19348 8830
rect 19292 8258 19348 8764
rect 19292 8206 19294 8258
rect 19346 8206 19348 8258
rect 18844 8194 18900 8204
rect 19292 8194 19348 8206
rect 19516 8260 19572 8270
rect 18172 8148 18228 8158
rect 18508 8148 18564 8158
rect 18172 8146 18564 8148
rect 18172 8094 18174 8146
rect 18226 8094 18510 8146
rect 18562 8094 18564 8146
rect 18172 8092 18564 8094
rect 18172 8082 18228 8092
rect 18508 8082 18564 8092
rect 17948 7534 17950 7586
rect 18002 7534 18004 7586
rect 17948 7522 18004 7534
rect 18060 7924 18116 7934
rect 18060 7476 18116 7868
rect 18284 7588 18340 7598
rect 18340 7532 18564 7588
rect 18172 7476 18228 7486
rect 18060 7474 18228 7476
rect 18060 7422 18174 7474
rect 18226 7422 18228 7474
rect 18060 7420 18228 7422
rect 18172 7410 18228 7420
rect 17276 7364 17332 7374
rect 17276 7252 17332 7308
rect 17388 7252 17444 7262
rect 17724 7252 17780 7262
rect 17276 7250 17444 7252
rect 17276 7198 17390 7250
rect 17442 7198 17444 7250
rect 17276 7196 17444 7198
rect 17164 6580 17220 6590
rect 17164 6486 17220 6524
rect 16940 6066 16996 6076
rect 16604 4174 16606 4226
rect 16658 4174 16660 4226
rect 16604 4162 16660 4174
rect 15372 3826 15428 3836
rect 16828 3780 16884 3790
rect 17276 3780 17332 7196
rect 17388 7186 17444 7196
rect 17612 7250 17780 7252
rect 17612 7198 17726 7250
rect 17778 7198 17780 7250
rect 17612 7196 17780 7198
rect 17388 5908 17444 5918
rect 17612 5908 17668 7196
rect 17724 7186 17780 7196
rect 18060 7252 18116 7262
rect 18284 7252 18340 7532
rect 18508 7474 18564 7532
rect 18844 7476 18900 7486
rect 18508 7422 18510 7474
rect 18562 7422 18564 7474
rect 18508 7410 18564 7422
rect 18732 7420 18844 7476
rect 18060 6690 18116 7196
rect 18060 6638 18062 6690
rect 18114 6638 18116 6690
rect 18060 6626 18116 6638
rect 18172 7196 18340 7252
rect 18396 7362 18452 7374
rect 18396 7310 18398 7362
rect 18450 7310 18452 7362
rect 18172 6468 18228 7196
rect 18396 7140 18452 7310
rect 18284 7084 18396 7140
rect 18284 6914 18340 7084
rect 18396 7074 18452 7084
rect 18284 6862 18286 6914
rect 18338 6862 18340 6914
rect 18284 6850 18340 6862
rect 18732 6916 18788 7420
rect 18844 7382 18900 7420
rect 19180 7474 19236 7486
rect 19180 7422 19182 7474
rect 19234 7422 19236 7474
rect 18732 6850 18788 6860
rect 18956 6804 19012 6814
rect 18956 6710 19012 6748
rect 18620 6692 18676 6702
rect 18620 6598 18676 6636
rect 18060 6412 18228 6468
rect 18396 6580 18452 6590
rect 17388 5906 17668 5908
rect 17388 5854 17390 5906
rect 17442 5854 17668 5906
rect 17388 5852 17668 5854
rect 17724 6132 17780 6142
rect 17388 5684 17444 5852
rect 17724 5796 17780 6076
rect 17388 5618 17444 5628
rect 17500 5740 17780 5796
rect 17500 5460 17556 5740
rect 17388 5404 17556 5460
rect 17388 4450 17444 5404
rect 17388 4398 17390 4450
rect 17442 4398 17444 4450
rect 17388 4386 17444 4398
rect 17500 4452 17556 4462
rect 17500 4358 17556 4396
rect 17724 4450 17780 4462
rect 17724 4398 17726 4450
rect 17778 4398 17780 4450
rect 17724 4340 17780 4398
rect 17836 4340 17892 4350
rect 17724 4338 17892 4340
rect 17724 4286 17838 4338
rect 17890 4286 17892 4338
rect 17724 4284 17892 4286
rect 18060 4340 18116 6412
rect 18396 6020 18452 6524
rect 19180 6356 19236 7422
rect 19180 6290 19236 6300
rect 18284 6018 18452 6020
rect 18284 5966 18398 6018
rect 18450 5966 18452 6018
rect 18284 5964 18452 5966
rect 18172 4564 18228 4574
rect 18284 4564 18340 5964
rect 18396 5954 18452 5964
rect 18732 6244 18788 6254
rect 18732 6018 18788 6188
rect 18732 5966 18734 6018
rect 18786 5966 18788 6018
rect 18732 5908 18788 5966
rect 18732 5842 18788 5852
rect 19068 6020 19124 6030
rect 18956 5684 19012 5694
rect 18396 5682 19012 5684
rect 18396 5630 18958 5682
rect 19010 5630 19012 5682
rect 18396 5628 19012 5630
rect 18396 5234 18452 5628
rect 18956 5618 19012 5628
rect 18396 5182 18398 5234
rect 18450 5182 18452 5234
rect 18396 5170 18452 5182
rect 18732 5236 18788 5246
rect 18732 5142 18788 5180
rect 18172 4562 18340 4564
rect 18172 4510 18174 4562
rect 18226 4510 18340 4562
rect 18172 4508 18340 4510
rect 18508 5012 18564 5022
rect 18172 4498 18228 4508
rect 18508 4450 18564 4956
rect 18508 4398 18510 4450
rect 18562 4398 18564 4450
rect 18508 4386 18564 4398
rect 19068 4450 19124 5964
rect 19292 5684 19348 5694
rect 19292 5590 19348 5628
rect 19516 5572 19572 8204
rect 19628 8146 19684 9884
rect 19852 9604 19908 9642
rect 19964 9604 20020 10332
rect 20636 10610 20804 10612
rect 20636 10558 20750 10610
rect 20802 10558 20804 10610
rect 20636 10556 20804 10558
rect 20636 10164 20692 10556
rect 20748 10546 20804 10556
rect 21084 10612 21140 10622
rect 21084 10518 21140 10556
rect 21420 10612 21476 10622
rect 21868 10612 21924 10622
rect 21420 10610 21924 10612
rect 21420 10558 21422 10610
rect 21474 10558 21870 10610
rect 21922 10558 21924 10610
rect 21420 10556 21924 10558
rect 21420 10546 21476 10556
rect 20636 10098 20692 10108
rect 20748 10386 20804 10398
rect 20748 10334 20750 10386
rect 20802 10334 20804 10386
rect 20748 9828 20804 10334
rect 21532 10164 21588 10174
rect 20748 9762 20804 9772
rect 21308 10052 21364 10062
rect 21308 9826 21364 9996
rect 21308 9774 21310 9826
rect 21362 9774 21364 9826
rect 21308 9762 21364 9774
rect 21532 9826 21588 10108
rect 21644 10052 21700 10556
rect 21868 10546 21924 10556
rect 21644 9986 21700 9996
rect 21980 10500 22036 10510
rect 21532 9774 21534 9826
rect 21586 9774 21588 9826
rect 21532 9762 21588 9774
rect 21644 9828 21700 9838
rect 21700 9772 21812 9828
rect 21644 9762 21700 9772
rect 21756 9714 21812 9772
rect 21980 9826 22036 10444
rect 22428 10498 22484 10510
rect 22428 10446 22430 10498
rect 22482 10446 22484 10498
rect 22428 10050 22484 10446
rect 22428 9998 22430 10050
rect 22482 9998 22484 10050
rect 22428 9986 22484 9998
rect 22652 9940 22708 9950
rect 22652 9846 22708 9884
rect 21980 9774 21982 9826
rect 22034 9774 22036 9826
rect 21980 9762 22036 9774
rect 21756 9662 21758 9714
rect 21810 9662 21812 9714
rect 21756 9650 21812 9662
rect 20636 9604 20692 9614
rect 19964 9548 20356 9604
rect 19852 9538 19908 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 9278
rect 19852 9156 19908 9166
rect 19852 9062 19908 9100
rect 20188 9042 20244 9212
rect 20188 8990 20190 9042
rect 20242 8990 20244 9042
rect 20188 8978 20244 8990
rect 20300 8930 20356 9548
rect 20300 8878 20302 8930
rect 20354 8878 20356 8930
rect 20300 8866 20356 8878
rect 20524 9602 20692 9604
rect 20524 9550 20638 9602
rect 20690 9550 20692 9602
rect 20524 9548 20692 9550
rect 20524 8260 20580 9548
rect 20636 9538 20692 9548
rect 21308 9604 21364 9614
rect 20748 9380 20804 9390
rect 20524 8194 20580 8204
rect 20636 9324 20748 9380
rect 19628 8094 19630 8146
rect 19682 8094 19684 8146
rect 19628 7588 19684 8094
rect 20188 8146 20244 8158
rect 20188 8094 20190 8146
rect 20242 8094 20244 8146
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19628 7522 19684 7532
rect 19740 7362 19796 7374
rect 19740 7310 19742 7362
rect 19794 7310 19796 7362
rect 19740 6468 19796 7310
rect 20188 6692 20244 8094
rect 20412 8036 20468 8046
rect 20412 7698 20468 7980
rect 20412 7646 20414 7698
rect 20466 7646 20468 7698
rect 20412 7634 20468 7646
rect 20524 8034 20580 8046
rect 20524 7982 20526 8034
rect 20578 7982 20580 8034
rect 20412 7364 20468 7374
rect 20412 7270 20468 7308
rect 20188 6626 20244 6636
rect 20300 6580 20356 6590
rect 20300 6486 20356 6524
rect 19740 6412 20244 6468
rect 20188 6356 20244 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20188 6290 20244 6300
rect 19836 6234 20100 6244
rect 20524 6018 20580 7982
rect 20636 7586 20692 9324
rect 20748 9314 20804 9324
rect 21196 9156 21252 9166
rect 21196 9044 21252 9100
rect 21084 9042 21252 9044
rect 21084 8990 21198 9042
rect 21250 8990 21252 9042
rect 21084 8988 21252 8990
rect 20636 7534 20638 7586
rect 20690 7534 20692 7586
rect 20636 7522 20692 7534
rect 20972 8148 21028 8158
rect 20972 7586 21028 8092
rect 20972 7534 20974 7586
rect 21026 7534 21028 7586
rect 20972 7522 21028 7534
rect 20748 7476 20804 7486
rect 20748 6692 20804 7420
rect 21084 7252 21140 8988
rect 21196 8978 21252 8988
rect 21308 8932 21364 9548
rect 21644 9602 21700 9614
rect 21644 9550 21646 9602
rect 21698 9550 21700 9602
rect 21644 9380 21700 9550
rect 21644 9314 21700 9324
rect 22652 9602 22708 9614
rect 22652 9550 22654 9602
rect 22706 9550 22708 9602
rect 21532 9268 21588 9278
rect 21532 9154 21588 9212
rect 21532 9102 21534 9154
rect 21586 9102 21588 9154
rect 21532 9090 21588 9102
rect 21644 9156 21700 9166
rect 21644 9062 21700 9100
rect 21308 8260 21364 8876
rect 22204 8932 22260 8942
rect 22204 8838 22260 8876
rect 21644 8818 21700 8830
rect 21644 8766 21646 8818
rect 21698 8766 21700 8818
rect 21644 8484 21700 8766
rect 21644 8418 21700 8428
rect 21084 7186 21140 7196
rect 21196 8258 21364 8260
rect 21196 8206 21310 8258
rect 21362 8206 21364 8258
rect 21196 8204 21364 8206
rect 20748 6626 20804 6636
rect 20524 5966 20526 6018
rect 20578 5966 20580 6018
rect 20524 5954 20580 5966
rect 19740 5906 19796 5918
rect 19740 5854 19742 5906
rect 19794 5854 19796 5906
rect 19740 5796 19796 5854
rect 19740 5730 19796 5740
rect 20636 5908 20692 5918
rect 19516 5516 19796 5572
rect 19068 4398 19070 4450
rect 19122 4398 19124 4450
rect 19068 4386 19124 4398
rect 19292 5124 19348 5134
rect 18172 4340 18228 4350
rect 18060 4338 18228 4340
rect 18060 4286 18174 4338
rect 18226 4286 18228 4338
rect 18060 4284 18228 4286
rect 17836 4274 17892 4284
rect 18172 4274 18228 4284
rect 17388 3780 17444 3790
rect 17276 3724 17388 3780
rect 16828 3686 16884 3724
rect 17388 3714 17444 3724
rect 13692 3500 14420 3556
rect 13580 3444 13636 3482
rect 13580 3378 13636 3388
rect 14364 800 14420 3500
rect 15708 3668 15764 3678
rect 15708 3442 15764 3612
rect 15708 3390 15710 3442
rect 15762 3390 15764 3442
rect 15708 3378 15764 3390
rect 19292 3442 19348 5068
rect 19740 5012 19796 5516
rect 19292 3390 19294 3442
rect 19346 3390 19348 3442
rect 19292 3388 19348 3390
rect 18844 3332 19348 3388
rect 19628 5010 19796 5012
rect 19628 4958 19742 5010
rect 19794 4958 19796 5010
rect 19628 4956 19796 4958
rect 18844 800 18900 3332
rect 19628 2996 19684 4956
rect 19740 4946 19796 4956
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20636 4564 20692 5852
rect 20748 5796 20804 5806
rect 20748 5234 20804 5740
rect 21196 5796 21252 8204
rect 21308 8194 21364 8204
rect 22092 8146 22148 8158
rect 22092 8094 22094 8146
rect 22146 8094 22148 8146
rect 21308 7700 21364 7710
rect 21308 7606 21364 7644
rect 21980 7586 22036 7598
rect 21980 7534 21982 7586
rect 22034 7534 22036 7586
rect 21420 7140 21476 7150
rect 21420 6578 21476 7084
rect 21420 6526 21422 6578
rect 21474 6526 21476 6578
rect 21420 6514 21476 6526
rect 21532 6690 21588 6702
rect 21532 6638 21534 6690
rect 21586 6638 21588 6690
rect 21196 5730 21252 5740
rect 20748 5182 20750 5234
rect 20802 5182 20804 5234
rect 20748 5170 20804 5182
rect 21420 5124 21476 5134
rect 21420 5030 21476 5068
rect 20748 4564 20804 4574
rect 20636 4562 20804 4564
rect 20636 4510 20750 4562
rect 20802 4510 20804 4562
rect 20636 4508 20804 4510
rect 20748 4498 20804 4508
rect 20188 4452 20244 4462
rect 20188 4226 20244 4396
rect 20188 4174 20190 4226
rect 20242 4174 20244 4226
rect 20188 4162 20244 4174
rect 20972 4452 21028 4462
rect 19964 4116 20020 4126
rect 19964 3554 20020 4060
rect 20748 3780 20804 3790
rect 20748 3686 20804 3724
rect 19964 3502 19966 3554
rect 20018 3502 20020 3554
rect 19964 3490 20020 3502
rect 20188 3444 20244 3482
rect 20188 3378 20244 3388
rect 20972 3442 21028 4396
rect 21308 4452 21364 4462
rect 21532 4452 21588 6638
rect 21756 5796 21812 5806
rect 21812 5740 21924 5796
rect 21756 5730 21812 5740
rect 21308 4450 21588 4452
rect 21308 4398 21310 4450
rect 21362 4398 21588 4450
rect 21308 4396 21588 4398
rect 21308 4386 21364 4396
rect 21532 4340 21588 4396
rect 21532 4274 21588 4284
rect 21868 4338 21924 5740
rect 21868 4286 21870 4338
rect 21922 4286 21924 4338
rect 21868 4274 21924 4286
rect 21084 3780 21140 3790
rect 21980 3780 22036 7534
rect 22092 7364 22148 8094
rect 22652 8036 22708 9550
rect 22652 7970 22708 7980
rect 22764 7924 22820 14140
rect 22988 13748 23044 14364
rect 23996 14420 24052 14430
rect 23996 14326 24052 14364
rect 24108 14418 24164 14430
rect 24108 14366 24110 14418
rect 24162 14366 24164 14418
rect 22988 13682 23044 13692
rect 23772 13188 23828 13198
rect 23100 12178 23156 12190
rect 23100 12126 23102 12178
rect 23154 12126 23156 12178
rect 22876 11956 22932 11966
rect 22876 11954 23044 11956
rect 22876 11902 22878 11954
rect 22930 11902 23044 11954
rect 22876 11900 23044 11902
rect 22876 11890 22932 11900
rect 22876 11620 22932 11630
rect 22876 11526 22932 11564
rect 22988 10834 23044 11900
rect 22988 10782 22990 10834
rect 23042 10782 23044 10834
rect 22988 10770 23044 10782
rect 23100 11394 23156 12126
rect 23548 12068 23604 12078
rect 23604 12012 23716 12068
rect 23548 11974 23604 12012
rect 23100 11342 23102 11394
rect 23154 11342 23156 11394
rect 22876 10500 22932 10510
rect 22876 10406 22932 10444
rect 22988 9044 23044 9054
rect 23100 9044 23156 11342
rect 23324 11732 23380 11742
rect 23212 11284 23268 11294
rect 23212 11190 23268 11228
rect 23212 10612 23268 10622
rect 23324 10612 23380 11676
rect 23212 10610 23380 10612
rect 23212 10558 23214 10610
rect 23266 10558 23380 10610
rect 23212 10556 23380 10558
rect 23660 11394 23716 12012
rect 23660 11342 23662 11394
rect 23714 11342 23716 11394
rect 23212 10546 23268 10556
rect 23660 9604 23716 11342
rect 23772 11060 23828 13132
rect 24108 13076 24164 14366
rect 24332 13636 24388 14478
rect 24332 13570 24388 13580
rect 24444 16268 24724 16324
rect 25340 16770 25508 16772
rect 25340 16718 25454 16770
rect 25506 16718 25508 16770
rect 25340 16716 25508 16718
rect 23884 12740 23940 12750
rect 24108 12740 24164 13020
rect 24220 12740 24276 12750
rect 24108 12738 24276 12740
rect 24108 12686 24222 12738
rect 24274 12686 24276 12738
rect 24108 12684 24276 12686
rect 23884 12180 23940 12684
rect 24220 12292 24276 12684
rect 24220 12226 24276 12236
rect 23884 12114 23940 12124
rect 24332 11284 24388 11294
rect 24332 11190 24388 11228
rect 23772 10994 23828 11004
rect 24108 9826 24164 9838
rect 24108 9774 24110 9826
rect 24162 9774 24164 9826
rect 23772 9604 23828 9614
rect 24108 9604 24164 9774
rect 23660 9602 24164 9604
rect 23660 9550 23774 9602
rect 23826 9550 24164 9602
rect 23660 9548 24164 9550
rect 24220 9828 24276 9838
rect 23324 9044 23380 9054
rect 23100 9042 23492 9044
rect 23100 8990 23326 9042
rect 23378 8990 23492 9042
rect 23100 8988 23492 8990
rect 22988 8950 23044 8988
rect 23324 8978 23380 8988
rect 22764 7858 22820 7868
rect 23324 8818 23380 8830
rect 23324 8766 23326 8818
rect 23378 8766 23380 8818
rect 22092 7298 22148 7308
rect 22988 7362 23044 7374
rect 22988 7310 22990 7362
rect 23042 7310 23044 7362
rect 22204 6692 22260 6702
rect 22204 6690 22708 6692
rect 22204 6638 22206 6690
rect 22258 6638 22708 6690
rect 22204 6636 22708 6638
rect 22204 6626 22260 6636
rect 22092 6468 22148 6478
rect 22540 6468 22596 6478
rect 22092 5122 22148 6412
rect 22092 5070 22094 5122
rect 22146 5070 22148 5122
rect 22092 5058 22148 5070
rect 22428 6466 22596 6468
rect 22428 6414 22542 6466
rect 22594 6414 22596 6466
rect 22428 6412 22596 6414
rect 22428 5124 22484 6412
rect 22540 6402 22596 6412
rect 22428 5058 22484 5068
rect 22540 6132 22596 6142
rect 22540 4450 22596 6076
rect 22652 5794 22708 6636
rect 22988 5906 23044 7310
rect 23212 7252 23268 7262
rect 22988 5854 22990 5906
rect 23042 5854 23044 5906
rect 22988 5842 23044 5854
rect 23100 7196 23212 7252
rect 23100 5908 23156 7196
rect 23212 7186 23268 7196
rect 23324 6804 23380 8766
rect 23324 6738 23380 6748
rect 23436 7700 23492 8988
rect 23772 8932 23828 9548
rect 24220 9492 24276 9772
rect 24108 9436 24276 9492
rect 23772 8866 23828 8876
rect 23884 9156 23940 9166
rect 23212 6690 23268 6702
rect 23212 6638 23214 6690
rect 23266 6638 23268 6690
rect 23212 6356 23268 6638
rect 23212 6290 23268 6300
rect 23212 5908 23268 5918
rect 23100 5906 23268 5908
rect 23100 5854 23214 5906
rect 23266 5854 23268 5906
rect 23100 5852 23268 5854
rect 22652 5742 22654 5794
rect 22706 5742 22708 5794
rect 22652 5730 22708 5742
rect 23212 5012 23268 5852
rect 23436 5906 23492 7644
rect 23660 8820 23716 8830
rect 23660 8148 23716 8764
rect 23660 7698 23716 8092
rect 23660 7646 23662 7698
rect 23714 7646 23716 7698
rect 23660 7634 23716 7646
rect 23548 6580 23604 6590
rect 23548 6018 23604 6524
rect 23772 6468 23828 6478
rect 23772 6374 23828 6412
rect 23884 6356 23940 9100
rect 24108 7698 24164 9436
rect 24220 8372 24276 8382
rect 24444 8372 24500 16268
rect 25340 15988 25396 16716
rect 25452 16706 25508 16716
rect 25228 15932 25396 15988
rect 24892 15874 24948 15886
rect 24892 15822 24894 15874
rect 24946 15822 24948 15874
rect 24556 15316 24612 15326
rect 24556 13074 24612 15260
rect 24668 15204 24724 15242
rect 24668 15138 24724 15148
rect 24668 14308 24724 14318
rect 24668 13634 24724 14252
rect 24668 13582 24670 13634
rect 24722 13582 24724 13634
rect 24668 13570 24724 13582
rect 24556 13022 24558 13074
rect 24610 13022 24612 13074
rect 24556 13010 24612 13022
rect 24892 10164 24948 15822
rect 25228 14868 25284 15932
rect 25564 15876 25620 16940
rect 25676 16772 25732 16782
rect 25676 15986 25732 16716
rect 25676 15934 25678 15986
rect 25730 15934 25732 15986
rect 25676 15922 25732 15934
rect 25340 15820 25620 15876
rect 25340 15314 25396 15820
rect 25900 15428 25956 15438
rect 25900 15334 25956 15372
rect 25340 15262 25342 15314
rect 25394 15262 25396 15314
rect 25340 15250 25396 15262
rect 25564 15316 25620 15326
rect 25564 15314 25844 15316
rect 25564 15262 25566 15314
rect 25618 15262 25844 15314
rect 25564 15260 25844 15262
rect 25564 15250 25620 15260
rect 25452 15204 25508 15214
rect 25228 14530 25284 14812
rect 25228 14478 25230 14530
rect 25282 14478 25284 14530
rect 25228 14466 25284 14478
rect 25340 15092 25508 15148
rect 25340 14980 25396 15092
rect 25340 14642 25396 14924
rect 25340 14590 25342 14642
rect 25394 14590 25396 14642
rect 25004 14420 25060 14430
rect 25060 14364 25172 14420
rect 25004 14354 25060 14364
rect 25116 13972 25172 14364
rect 25228 13972 25284 13982
rect 25116 13970 25284 13972
rect 25116 13918 25230 13970
rect 25282 13918 25284 13970
rect 25116 13916 25284 13918
rect 25228 13906 25284 13916
rect 25004 12962 25060 12974
rect 25004 12910 25006 12962
rect 25058 12910 25060 12962
rect 25004 12740 25060 12910
rect 25004 12674 25060 12684
rect 24892 10108 25060 10164
rect 24892 9940 24948 9950
rect 24892 9846 24948 9884
rect 24668 9156 24724 9166
rect 24668 9062 24724 9100
rect 24220 8370 24500 8372
rect 24220 8318 24222 8370
rect 24274 8318 24500 8370
rect 24220 8316 24500 8318
rect 24556 8932 24612 8942
rect 24220 8306 24276 8316
rect 24108 7646 24110 7698
rect 24162 7646 24164 7698
rect 23884 6290 23940 6300
rect 23996 6802 24052 6814
rect 23996 6750 23998 6802
rect 24050 6750 24052 6802
rect 23996 6132 24052 6750
rect 24108 6356 24164 7646
rect 24556 8260 24612 8876
rect 24892 8260 24948 8270
rect 24556 8258 24948 8260
rect 24556 8206 24894 8258
rect 24946 8206 24948 8258
rect 24556 8204 24948 8206
rect 24556 7698 24612 8204
rect 24892 8194 24948 8204
rect 24556 7646 24558 7698
rect 24610 7646 24612 7698
rect 24556 7634 24612 7646
rect 24108 6290 24164 6300
rect 24220 7588 24276 7598
rect 23996 6066 24052 6076
rect 24220 6130 24276 7532
rect 25004 7476 25060 10108
rect 25228 9156 25284 9166
rect 25340 9156 25396 14590
rect 25564 14308 25620 14318
rect 25564 13858 25620 14252
rect 25564 13806 25566 13858
rect 25618 13806 25620 13858
rect 25564 13794 25620 13806
rect 25676 14196 25732 14206
rect 25676 12964 25732 14140
rect 25788 13412 25844 15260
rect 26012 15090 26068 15102
rect 26012 15038 26014 15090
rect 26066 15038 26068 15090
rect 26012 14530 26068 15038
rect 26124 15090 26180 15102
rect 26124 15038 26126 15090
rect 26178 15038 26180 15090
rect 26124 14868 26180 15038
rect 26124 14802 26180 14812
rect 26012 14478 26014 14530
rect 26066 14478 26068 14530
rect 26012 14466 26068 14478
rect 26236 14530 26292 19852
rect 26348 19236 26404 21308
rect 26572 21140 26628 21150
rect 26460 20804 26516 20814
rect 26460 20710 26516 20748
rect 26572 20802 26628 21084
rect 26684 20914 26740 21534
rect 26684 20862 26686 20914
rect 26738 20862 26740 20914
rect 26684 20850 26740 20862
rect 26572 20750 26574 20802
rect 26626 20750 26628 20802
rect 26572 20738 26628 20750
rect 26348 19170 26404 19180
rect 26572 20580 26628 20590
rect 26796 20580 26852 20590
rect 26460 18452 26516 18462
rect 26460 18358 26516 18396
rect 26572 17892 26628 20524
rect 26684 20578 26852 20580
rect 26684 20526 26798 20578
rect 26850 20526 26852 20578
rect 26684 20524 26852 20526
rect 26684 20244 26740 20524
rect 26796 20514 26852 20524
rect 26908 20580 26964 21644
rect 26908 20514 26964 20524
rect 26684 20178 26740 20188
rect 26796 20130 26852 20142
rect 26796 20078 26798 20130
rect 26850 20078 26852 20130
rect 26796 19684 26852 20078
rect 26908 20020 26964 20030
rect 26908 19926 26964 19964
rect 27020 19908 27076 22988
rect 27132 22146 27188 22158
rect 27132 22094 27134 22146
rect 27186 22094 27188 22146
rect 27132 21812 27188 22094
rect 27244 22036 27300 23212
rect 27356 23266 27412 23662
rect 27804 23714 27860 23772
rect 27804 23662 27806 23714
rect 27858 23662 27860 23714
rect 27804 23650 27860 23662
rect 27356 23214 27358 23266
rect 27410 23214 27412 23266
rect 27356 23202 27412 23214
rect 27468 23044 27524 23054
rect 27468 22370 27524 22988
rect 27916 22708 27972 29820
rect 28028 27972 28084 30044
rect 28140 29650 28196 32284
rect 28252 31108 28308 31118
rect 28476 31108 28532 33180
rect 28812 33124 28868 34188
rect 28924 34130 28980 34142
rect 28924 34078 28926 34130
rect 28978 34078 28980 34130
rect 28924 34020 28980 34078
rect 29036 34132 29092 34142
rect 29036 34038 29092 34076
rect 29260 34132 29316 34142
rect 29260 34038 29316 34076
rect 28924 33954 28980 33964
rect 28252 31106 28532 31108
rect 28252 31054 28254 31106
rect 28306 31054 28532 31106
rect 28252 31052 28532 31054
rect 28700 33068 28868 33124
rect 28924 33684 28980 33694
rect 28924 33124 28980 33628
rect 29372 33460 29428 34412
rect 29260 33458 29428 33460
rect 29260 33406 29374 33458
rect 29426 33406 29428 33458
rect 29260 33404 29428 33406
rect 28252 31042 28308 31052
rect 28140 29598 28142 29650
rect 28194 29598 28196 29650
rect 28140 29586 28196 29598
rect 28476 30772 28532 30782
rect 28028 27906 28084 27916
rect 28364 29426 28420 29438
rect 28364 29374 28366 29426
rect 28418 29374 28420 29426
rect 28252 25732 28308 25742
rect 28028 25620 28084 25630
rect 28028 25526 28084 25564
rect 28140 25508 28196 25518
rect 28140 25414 28196 25452
rect 27916 22642 27972 22652
rect 28028 25284 28084 25294
rect 27916 22484 27972 22494
rect 28028 22484 28084 25228
rect 28252 24836 28308 25676
rect 28140 24780 28308 24836
rect 28140 24164 28196 24780
rect 28252 24612 28308 24622
rect 28252 24518 28308 24556
rect 28364 24276 28420 29374
rect 28476 26908 28532 30716
rect 28476 26852 28644 26908
rect 28476 26740 28532 26750
rect 28476 25506 28532 26684
rect 28476 25454 28478 25506
rect 28530 25454 28532 25506
rect 28476 25442 28532 25454
rect 28588 25508 28644 26852
rect 28588 25284 28644 25452
rect 28364 24210 28420 24220
rect 28476 25228 28644 25284
rect 28700 26178 28756 33068
rect 28812 30212 28868 30222
rect 28812 29426 28868 30156
rect 28812 29374 28814 29426
rect 28866 29374 28868 29426
rect 28812 29362 28868 29374
rect 28700 26126 28702 26178
rect 28754 26126 28756 26178
rect 28140 24108 28308 24164
rect 28252 24052 28308 24108
rect 28364 24052 28420 24062
rect 28252 24050 28420 24052
rect 28252 23998 28366 24050
rect 28418 23998 28420 24050
rect 28252 23996 28420 23998
rect 28364 23986 28420 23996
rect 27916 22482 28084 22484
rect 27916 22430 27918 22482
rect 27970 22430 28084 22482
rect 27916 22428 28084 22430
rect 28140 22932 28196 22942
rect 27916 22418 27972 22428
rect 27468 22318 27470 22370
rect 27522 22318 27524 22370
rect 27468 22306 27524 22318
rect 27244 21970 27300 21980
rect 27804 22036 27860 22046
rect 27132 21746 27188 21756
rect 27580 21812 27636 21822
rect 27580 21698 27636 21756
rect 27804 21810 27860 21980
rect 27804 21758 27806 21810
rect 27858 21758 27860 21810
rect 27804 21746 27860 21758
rect 27580 21646 27582 21698
rect 27634 21646 27636 21698
rect 27580 21634 27636 21646
rect 28028 21588 28084 21598
rect 28028 21494 28084 21532
rect 28140 20916 28196 22876
rect 28252 22370 28308 22382
rect 28252 22318 28254 22370
rect 28306 22318 28308 22370
rect 28252 21698 28308 22318
rect 28252 21646 28254 21698
rect 28306 21646 28308 21698
rect 28252 21364 28308 21646
rect 28364 21476 28420 21486
rect 28364 21382 28420 21420
rect 28252 21298 28308 21308
rect 27916 20860 28196 20916
rect 28252 21140 28308 21150
rect 28252 20914 28308 21084
rect 28252 20862 28254 20914
rect 28306 20862 28308 20914
rect 27244 20804 27300 20814
rect 27244 20242 27300 20748
rect 27804 20802 27860 20814
rect 27804 20750 27806 20802
rect 27858 20750 27860 20802
rect 27804 20356 27860 20750
rect 27804 20290 27860 20300
rect 27244 20190 27246 20242
rect 27298 20190 27300 20242
rect 27244 20178 27300 20190
rect 27468 20132 27860 20188
rect 27916 20132 27972 20860
rect 28252 20850 28308 20862
rect 28028 20692 28084 20702
rect 28084 20636 28196 20692
rect 28028 20626 28084 20636
rect 27356 20018 27412 20030
rect 27356 19966 27358 20018
rect 27410 19966 27412 20018
rect 27132 19908 27188 19918
rect 27020 19852 27132 19908
rect 26796 19618 26852 19628
rect 26796 19346 26852 19358
rect 26796 19294 26798 19346
rect 26850 19294 26852 19346
rect 26684 19234 26740 19246
rect 26684 19182 26686 19234
rect 26738 19182 26740 19234
rect 26684 18900 26740 19182
rect 26684 18834 26740 18844
rect 26796 18564 26852 19294
rect 26236 14478 26238 14530
rect 26290 14478 26292 14530
rect 25788 13346 25844 13356
rect 26124 13636 26180 13646
rect 26236 13636 26292 14478
rect 26124 13634 26292 13636
rect 26124 13582 26126 13634
rect 26178 13582 26292 13634
rect 26124 13580 26292 13582
rect 26348 17836 26628 17892
rect 26684 18508 26852 18564
rect 27020 18900 27076 18910
rect 26684 18450 26740 18508
rect 26908 18452 26964 18462
rect 26684 18398 26686 18450
rect 26738 18398 26740 18450
rect 26124 13188 26180 13580
rect 25564 12962 25732 12964
rect 25564 12910 25678 12962
rect 25730 12910 25732 12962
rect 25564 12908 25732 12910
rect 25452 12852 25508 12862
rect 25452 12758 25508 12796
rect 25452 12404 25508 12414
rect 25564 12404 25620 12908
rect 25676 12898 25732 12908
rect 25788 13132 26180 13188
rect 25452 12402 25620 12404
rect 25452 12350 25454 12402
rect 25506 12350 25620 12402
rect 25452 12348 25620 12350
rect 25452 12338 25508 12348
rect 25788 9828 25844 13132
rect 26348 13076 26404 17836
rect 26460 17444 26516 17454
rect 26460 16098 26516 17388
rect 26684 17332 26740 18398
rect 26796 18450 26964 18452
rect 26796 18398 26910 18450
rect 26962 18398 26964 18450
rect 26796 18396 26964 18398
rect 26796 18116 26852 18396
rect 26908 18386 26964 18396
rect 26796 18050 26852 18060
rect 27020 17892 27076 18844
rect 27132 18676 27188 19852
rect 27356 19796 27412 19966
rect 27468 20020 27524 20132
rect 27804 20130 27972 20132
rect 27804 20078 27806 20130
rect 27858 20078 27972 20130
rect 27804 20076 27972 20078
rect 28028 20132 28084 20142
rect 27804 20066 27860 20076
rect 27468 19954 27524 19964
rect 27692 20020 27748 20030
rect 27580 19908 27636 19918
rect 27580 19796 27636 19852
rect 27356 19740 27636 19796
rect 27356 19124 27412 19740
rect 27692 19684 27748 19964
rect 27692 19618 27748 19628
rect 28028 19458 28084 20076
rect 28028 19406 28030 19458
rect 28082 19406 28084 19458
rect 28028 19394 28084 19406
rect 28140 19236 28196 20636
rect 28252 20020 28308 20030
rect 28252 19926 28308 19964
rect 27916 19180 28196 19236
rect 28364 19234 28420 19246
rect 28364 19182 28366 19234
rect 28418 19182 28420 19234
rect 27356 19030 27412 19068
rect 27692 19124 27748 19134
rect 27692 19030 27748 19068
rect 27132 18610 27188 18620
rect 27692 18676 27748 18686
rect 27692 18582 27748 18620
rect 27020 17826 27076 17836
rect 27468 17780 27524 17790
rect 27020 17666 27076 17678
rect 27020 17614 27022 17666
rect 27074 17614 27076 17666
rect 26684 17266 26740 17276
rect 26796 17556 26852 17566
rect 26460 16046 26462 16098
rect 26514 16046 26516 16098
rect 26460 16034 26516 16046
rect 26796 15316 26852 17500
rect 26908 17554 26964 17566
rect 26908 17502 26910 17554
rect 26962 17502 26964 17554
rect 26908 15538 26964 17502
rect 27020 17444 27076 17614
rect 27468 17666 27524 17724
rect 27468 17614 27470 17666
rect 27522 17614 27524 17666
rect 27468 17602 27524 17614
rect 27916 17668 27972 19180
rect 28252 18900 28308 18910
rect 28252 18340 28308 18844
rect 28364 18788 28420 19182
rect 28364 18722 28420 18732
rect 28476 18340 28532 25228
rect 28700 22148 28756 26126
rect 28812 24948 28868 24958
rect 28812 24854 28868 24892
rect 28700 22082 28756 22092
rect 28812 23268 28868 23278
rect 28700 21700 28756 21710
rect 28700 21586 28756 21644
rect 28700 21534 28702 21586
rect 28754 21534 28756 21586
rect 28700 21364 28756 21534
rect 28700 20242 28756 21308
rect 28700 20190 28702 20242
rect 28754 20190 28756 20242
rect 28700 20178 28756 20190
rect 28812 20020 28868 23212
rect 28812 19954 28868 19964
rect 28924 19460 28980 33068
rect 29148 33236 29204 33246
rect 29148 32786 29204 33180
rect 29148 32734 29150 32786
rect 29202 32734 29204 32786
rect 29148 32722 29204 32734
rect 29148 26964 29204 26974
rect 29260 26964 29316 33404
rect 29372 33394 29428 33404
rect 29372 33012 29428 33022
rect 29372 30100 29428 32956
rect 29484 30324 29540 34524
rect 29596 33236 29652 35420
rect 29820 35476 29876 35486
rect 29820 35308 29876 35420
rect 29708 35252 29876 35308
rect 29932 35364 29988 35532
rect 30044 35522 30100 35532
rect 30268 35476 30324 36092
rect 30380 35700 30436 36430
rect 31164 36258 31220 36270
rect 31164 36206 31166 36258
rect 31218 36206 31220 36258
rect 31052 36036 31108 36046
rect 31164 36036 31220 36206
rect 31500 36036 31556 37100
rect 31724 37156 31780 37166
rect 31724 37154 31892 37156
rect 31724 37102 31726 37154
rect 31778 37102 31892 37154
rect 31724 37100 31892 37102
rect 31724 37090 31780 37100
rect 31164 35980 31556 36036
rect 30940 35924 30996 35934
rect 30940 35830 30996 35868
rect 30380 35634 30436 35644
rect 30492 35700 30548 35710
rect 30492 35698 30660 35700
rect 30492 35646 30494 35698
rect 30546 35646 30660 35698
rect 30492 35644 30660 35646
rect 30492 35634 30548 35644
rect 30156 35420 30324 35476
rect 30492 35476 30548 35486
rect 30156 35364 30212 35420
rect 29932 35298 29988 35308
rect 30044 35308 30212 35364
rect 29708 35140 29764 35252
rect 29708 35084 29988 35140
rect 29708 34914 29764 34926
rect 29708 34862 29710 34914
rect 29762 34862 29764 34914
rect 29708 34580 29764 34862
rect 29820 34804 29876 34814
rect 29820 34710 29876 34748
rect 29708 34514 29764 34524
rect 29708 34356 29764 34366
rect 29708 34132 29764 34300
rect 29820 34132 29876 34142
rect 29708 34130 29876 34132
rect 29708 34078 29822 34130
rect 29874 34078 29876 34130
rect 29708 34076 29876 34078
rect 29708 33684 29764 34076
rect 29820 34066 29876 34076
rect 29932 33908 29988 35084
rect 29708 33618 29764 33628
rect 29820 33852 29988 33908
rect 29708 33236 29764 33246
rect 29596 33234 29764 33236
rect 29596 33182 29710 33234
rect 29762 33182 29764 33234
rect 29596 33180 29764 33182
rect 29708 33170 29764 33180
rect 29820 33012 29876 33852
rect 29708 32956 29876 33012
rect 29932 33348 29988 33358
rect 29932 33012 29988 33292
rect 29596 32452 29652 32462
rect 29596 32358 29652 32396
rect 29708 31668 29764 32956
rect 29932 32946 29988 32956
rect 29932 32676 29988 32686
rect 30044 32676 30100 35308
rect 30492 34914 30548 35420
rect 30492 34862 30494 34914
rect 30546 34862 30548 34914
rect 30492 34850 30548 34862
rect 30268 34468 30324 34478
rect 30268 34018 30324 34412
rect 30268 33966 30270 34018
rect 30322 33966 30324 34018
rect 30268 33954 30324 33966
rect 30380 34018 30436 34030
rect 30380 33966 30382 34018
rect 30434 33966 30436 34018
rect 30380 33460 30436 33966
rect 30604 33684 30660 35644
rect 30828 35474 30884 35486
rect 30828 35422 30830 35474
rect 30882 35422 30884 35474
rect 30828 34580 30884 35422
rect 31052 34914 31108 35980
rect 31388 35812 31444 35822
rect 31388 35588 31444 35756
rect 31052 34862 31054 34914
rect 31106 34862 31108 34914
rect 31052 34850 31108 34862
rect 31276 35586 31444 35588
rect 31276 35534 31390 35586
rect 31442 35534 31444 35586
rect 31276 35532 31444 35534
rect 31052 34692 31108 34702
rect 30828 34514 30884 34524
rect 30940 34690 31108 34692
rect 30940 34638 31054 34690
rect 31106 34638 31108 34690
rect 30940 34636 31108 34638
rect 30940 34242 30996 34636
rect 31052 34626 31108 34636
rect 30940 34190 30942 34242
rect 30994 34190 30996 34242
rect 30940 34178 30996 34190
rect 31052 34130 31108 34142
rect 31052 34078 31054 34130
rect 31106 34078 31108 34130
rect 30604 33618 30660 33628
rect 30716 34020 30772 34030
rect 30380 33394 30436 33404
rect 30716 33236 30772 33964
rect 31052 34020 31108 34078
rect 31052 33954 31108 33964
rect 30940 33348 30996 33358
rect 30940 33254 30996 33292
rect 30716 33142 30772 33180
rect 30604 32900 30660 32910
rect 30604 32786 30660 32844
rect 30604 32734 30606 32786
rect 30658 32734 30660 32786
rect 30604 32722 30660 32734
rect 29932 32674 30100 32676
rect 29932 32622 29934 32674
rect 29986 32622 30100 32674
rect 29932 32620 30100 32622
rect 29932 32610 29988 32620
rect 30156 32562 30212 32574
rect 30156 32510 30158 32562
rect 30210 32510 30212 32562
rect 29932 31668 29988 31678
rect 29708 31666 29988 31668
rect 29708 31614 29934 31666
rect 29986 31614 29988 31666
rect 29708 31612 29988 31614
rect 29932 31602 29988 31612
rect 30044 31220 30100 31230
rect 30156 31220 30212 32510
rect 30940 32562 30996 32574
rect 30940 32510 30942 32562
rect 30994 32510 30996 32562
rect 30268 31780 30324 31790
rect 30268 31778 30884 31780
rect 30268 31726 30270 31778
rect 30322 31726 30884 31778
rect 30268 31724 30884 31726
rect 30268 31714 30324 31724
rect 30604 31556 30660 31566
rect 30604 31220 30660 31500
rect 30828 31220 30884 31724
rect 30940 31556 30996 32510
rect 31164 31778 31220 31790
rect 31164 31726 31166 31778
rect 31218 31726 31220 31778
rect 31164 31668 31220 31726
rect 31164 31602 31220 31612
rect 30940 31490 30996 31500
rect 31276 31332 31332 35532
rect 31388 35522 31444 35532
rect 31500 34914 31556 35980
rect 31612 36258 31668 36270
rect 31612 36206 31614 36258
rect 31666 36206 31668 36258
rect 31612 35474 31668 36206
rect 31836 35812 31892 37100
rect 32060 37154 32116 37166
rect 32060 37102 32062 37154
rect 32114 37102 32116 37154
rect 32060 36372 32116 37102
rect 32284 36708 32340 38444
rect 32396 38612 32452 38622
rect 32396 36932 32452 38556
rect 32508 37156 32564 37166
rect 32508 37062 32564 37100
rect 32396 36876 32564 36932
rect 32396 36708 32452 36718
rect 32284 36706 32452 36708
rect 32284 36654 32398 36706
rect 32450 36654 32452 36706
rect 32284 36652 32452 36654
rect 32396 36642 32452 36652
rect 32172 36372 32228 36382
rect 32060 36370 32228 36372
rect 32060 36318 32174 36370
rect 32226 36318 32228 36370
rect 32060 36316 32228 36318
rect 32172 36148 32228 36316
rect 32172 36092 32452 36148
rect 32060 35980 32340 36036
rect 31948 35812 32004 35822
rect 31836 35756 31948 35812
rect 31948 35718 32004 35756
rect 31612 35422 31614 35474
rect 31666 35422 31668 35474
rect 31612 35410 31668 35422
rect 31724 35700 31780 35710
rect 31500 34862 31502 34914
rect 31554 34862 31556 34914
rect 31500 34244 31556 34862
rect 31612 34468 31668 34478
rect 31612 34354 31668 34412
rect 31612 34302 31614 34354
rect 31666 34302 31668 34354
rect 31612 34290 31668 34302
rect 31500 34178 31556 34188
rect 31724 33236 31780 35644
rect 31948 34244 32004 34254
rect 32060 34244 32116 35980
rect 32284 35922 32340 35980
rect 32284 35870 32286 35922
rect 32338 35870 32340 35922
rect 32284 35858 32340 35870
rect 32396 35812 32452 36092
rect 32284 35700 32340 35710
rect 32284 35606 32340 35644
rect 32396 35476 32452 35756
rect 32508 35810 32564 36876
rect 32508 35758 32510 35810
rect 32562 35758 32564 35810
rect 32508 35746 32564 35758
rect 31948 34242 32116 34244
rect 31948 34190 31950 34242
rect 32002 34190 32116 34242
rect 31948 34188 32116 34190
rect 32172 35420 32452 35476
rect 31948 34178 32004 34188
rect 32060 34020 32116 34030
rect 32060 33926 32116 33964
rect 31724 33170 31780 33180
rect 31500 33124 31556 33134
rect 31500 33030 31556 33068
rect 32172 32900 32228 35420
rect 32620 35026 32676 40348
rect 32956 37828 33012 41918
rect 33516 41970 33684 41972
rect 33516 41918 33630 41970
rect 33682 41918 33684 41970
rect 33516 41916 33684 41918
rect 33404 41188 33460 41198
rect 33292 41186 33460 41188
rect 33292 41134 33406 41186
rect 33458 41134 33460 41186
rect 33292 41132 33460 41134
rect 33068 40962 33124 40974
rect 33068 40910 33070 40962
rect 33122 40910 33124 40962
rect 33068 40514 33124 40910
rect 33068 40462 33070 40514
rect 33122 40462 33124 40514
rect 33068 40450 33124 40462
rect 33068 38724 33124 38734
rect 33124 38668 33236 38724
rect 33068 38658 33124 38668
rect 32956 37762 33012 37772
rect 33068 37266 33124 37278
rect 33068 37214 33070 37266
rect 33122 37214 33124 37266
rect 33068 37156 33124 37214
rect 33068 36708 33124 37100
rect 33068 36642 33124 36652
rect 33180 36594 33236 38668
rect 33292 38500 33348 41132
rect 33404 41122 33460 41132
rect 33404 40628 33460 40638
rect 33516 40628 33572 41916
rect 33628 41906 33684 41916
rect 33404 40626 33572 40628
rect 33404 40574 33406 40626
rect 33458 40574 33572 40626
rect 33404 40572 33572 40574
rect 33404 40562 33460 40572
rect 33292 38434 33348 38444
rect 33852 38500 33908 38510
rect 33852 38162 33908 38444
rect 33964 38388 34020 44044
rect 34076 44034 34132 44044
rect 34300 43650 34356 44156
rect 34300 43598 34302 43650
rect 34354 43598 34356 43650
rect 34300 43586 34356 43598
rect 34412 43652 34468 44270
rect 34636 43988 34692 46398
rect 34860 44324 34916 46732
rect 35196 46722 35252 46732
rect 35756 46786 35812 48188
rect 36204 48802 36260 48814
rect 36204 48750 36206 48802
rect 36258 48750 36260 48802
rect 35980 47236 36036 47246
rect 36204 47236 36260 48750
rect 36036 47180 36260 47236
rect 35980 47142 36036 47180
rect 35756 46734 35758 46786
rect 35810 46734 35812 46786
rect 35756 46722 35812 46734
rect 37100 47012 37156 48974
rect 37548 49026 37604 49038
rect 37548 48974 37550 49026
rect 37602 48974 37604 49026
rect 37548 48466 37604 48974
rect 37548 48414 37550 48466
rect 37602 48414 37604 48466
rect 37548 48402 37604 48414
rect 40012 48802 40068 48814
rect 40460 48804 40516 48814
rect 40012 48750 40014 48802
rect 40066 48750 40068 48802
rect 38892 48356 38948 48366
rect 38892 48262 38948 48300
rect 39900 48354 39956 48366
rect 39900 48302 39902 48354
rect 39954 48302 39956 48354
rect 37324 48244 37380 48254
rect 37996 48244 38052 48254
rect 37324 48242 38052 48244
rect 37324 48190 37326 48242
rect 37378 48190 37998 48242
rect 38050 48190 38052 48242
rect 37324 48188 38052 48190
rect 37324 48178 37380 48188
rect 37996 48178 38052 48188
rect 38780 48242 38836 48254
rect 39564 48244 39620 48254
rect 38780 48190 38782 48242
rect 38834 48190 38836 48242
rect 38332 48018 38388 48030
rect 38332 47966 38334 48018
rect 38386 47966 38388 48018
rect 37996 47346 38052 47358
rect 37996 47294 37998 47346
rect 38050 47294 38052 47346
rect 37996 47236 38052 47294
rect 38220 47348 38276 47358
rect 38220 47254 38276 47292
rect 37996 47170 38052 47180
rect 38332 47236 38388 47966
rect 38332 47170 38388 47180
rect 38556 47458 38612 47470
rect 38556 47406 38558 47458
rect 38610 47406 38612 47458
rect 34972 46564 35028 46574
rect 34972 46470 35028 46508
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 37100 45890 37156 46956
rect 38556 46788 38612 47406
rect 38780 47348 38836 48190
rect 39004 48242 39620 48244
rect 39004 48190 39566 48242
rect 39618 48190 39620 48242
rect 39004 48188 39620 48190
rect 38892 47684 38948 47694
rect 39004 47684 39060 48188
rect 39564 48178 39620 48188
rect 38892 47682 39060 47684
rect 38892 47630 38894 47682
rect 38946 47630 39060 47682
rect 38892 47628 39060 47630
rect 38892 47618 38948 47628
rect 39228 47458 39284 47470
rect 39228 47406 39230 47458
rect 39282 47406 39284 47458
rect 38892 47348 38948 47358
rect 38780 47292 38892 47348
rect 38668 46788 38724 46798
rect 38556 46732 38668 46788
rect 38668 46694 38724 46732
rect 38892 46674 38948 47292
rect 39228 47012 39284 47406
rect 39900 47458 39956 48302
rect 40012 48356 40068 48750
rect 40012 48020 40068 48300
rect 40236 48802 40516 48804
rect 40236 48750 40462 48802
rect 40514 48750 40516 48802
rect 40236 48748 40516 48750
rect 40124 48020 40180 48030
rect 40012 48018 40180 48020
rect 40012 47966 40126 48018
rect 40178 47966 40180 48018
rect 40012 47964 40180 47966
rect 40124 47954 40180 47964
rect 39900 47406 39902 47458
rect 39954 47406 39956 47458
rect 39900 47394 39956 47406
rect 40236 47012 40292 48748
rect 40460 48738 40516 48748
rect 39284 46956 39508 47012
rect 39228 46946 39284 46956
rect 39452 46898 39508 46956
rect 39452 46846 39454 46898
rect 39506 46846 39508 46898
rect 39452 46834 39508 46846
rect 40236 46898 40292 46956
rect 40236 46846 40238 46898
rect 40290 46846 40292 46898
rect 40236 46834 40292 46846
rect 40348 48130 40404 48142
rect 40348 48078 40350 48130
rect 40402 48078 40404 48130
rect 40348 48018 40404 48078
rect 40348 47966 40350 48018
rect 40402 47966 40404 48018
rect 38892 46622 38894 46674
rect 38946 46622 38948 46674
rect 37772 46452 37828 46462
rect 37772 46450 38052 46452
rect 37772 46398 37774 46450
rect 37826 46398 38052 46450
rect 37772 46396 38052 46398
rect 37772 46386 37828 46396
rect 37100 45838 37102 45890
rect 37154 45838 37156 45890
rect 37100 45826 37156 45838
rect 37660 45892 37716 45902
rect 37660 45890 37828 45892
rect 37660 45838 37662 45890
rect 37714 45838 37828 45890
rect 37660 45836 37828 45838
rect 37660 45826 37716 45836
rect 34636 43922 34692 43932
rect 34748 44322 34916 44324
rect 34748 44270 34862 44322
rect 34914 44270 34916 44322
rect 34748 44268 34916 44270
rect 34412 43586 34468 43596
rect 34076 43540 34132 43550
rect 34076 43446 34132 43484
rect 34188 41412 34244 41422
rect 34076 41186 34132 41198
rect 34076 41134 34078 41186
rect 34130 41134 34132 41186
rect 34076 41076 34132 41134
rect 34076 40292 34132 41020
rect 34188 41076 34244 41356
rect 34188 41074 34468 41076
rect 34188 41022 34190 41074
rect 34242 41022 34468 41074
rect 34188 41020 34468 41022
rect 34188 41010 34244 41020
rect 34076 40226 34132 40236
rect 34412 38836 34468 41020
rect 34524 39396 34580 39406
rect 34524 39302 34580 39340
rect 34748 38946 34804 44268
rect 34860 44258 34916 44268
rect 34972 45332 35028 45342
rect 34972 44212 35028 45276
rect 37436 45332 37492 45342
rect 37436 45238 37492 45276
rect 37772 45330 37828 45836
rect 37772 45278 37774 45330
rect 37826 45278 37828 45330
rect 37772 45266 37828 45278
rect 34972 44118 35028 44156
rect 35084 45106 35140 45118
rect 35084 45054 35086 45106
rect 35138 45054 35140 45106
rect 35084 44100 35140 45054
rect 37996 45106 38052 46396
rect 38108 46450 38164 46462
rect 38108 46398 38110 46450
rect 38162 46398 38164 46450
rect 38108 45332 38164 46398
rect 38108 45266 38164 45276
rect 37996 45054 37998 45106
rect 38050 45054 38052 45106
rect 37996 45042 38052 45054
rect 38892 44996 38948 46622
rect 40012 46788 40068 46798
rect 40012 46116 40068 46732
rect 40348 46676 40404 47966
rect 40012 46002 40068 46060
rect 40012 45950 40014 46002
rect 40066 45950 40068 46002
rect 40012 45938 40068 45950
rect 40236 46620 40404 46676
rect 41692 47236 41748 47246
rect 39788 45220 39844 45230
rect 39788 45106 39844 45164
rect 39788 45054 39790 45106
rect 39842 45054 39844 45106
rect 39788 45042 39844 45054
rect 39340 44996 39396 45006
rect 38892 44994 39396 44996
rect 38892 44942 39342 44994
rect 39394 44942 39396 44994
rect 38892 44940 39396 44942
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35868 44324 35924 44334
rect 35084 44034 35140 44044
rect 35196 44322 35924 44324
rect 35196 44270 35870 44322
rect 35922 44270 35924 44322
rect 35196 44268 35924 44270
rect 34860 43652 34916 43662
rect 34860 43538 34916 43596
rect 35196 43650 35252 44268
rect 35868 44258 35924 44268
rect 35644 44100 35700 44110
rect 35644 44006 35700 44044
rect 35196 43598 35198 43650
rect 35250 43598 35252 43650
rect 35196 43586 35252 43598
rect 36316 43764 36372 43774
rect 34860 43486 34862 43538
rect 34914 43486 34916 43538
rect 34860 43474 34916 43486
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 36316 42866 36372 43708
rect 36316 42814 36318 42866
rect 36370 42814 36372 42866
rect 36316 42802 36372 42814
rect 37996 43650 38052 43662
rect 37996 43598 37998 43650
rect 38050 43598 38052 43650
rect 37772 42754 37828 42766
rect 37772 42702 37774 42754
rect 37826 42702 37828 42754
rect 35308 42644 35364 42654
rect 34972 42642 35364 42644
rect 34972 42590 35310 42642
rect 35362 42590 35364 42642
rect 34972 42588 35364 42590
rect 34972 41410 35028 42588
rect 35308 42578 35364 42588
rect 35644 42530 35700 42542
rect 35644 42478 35646 42530
rect 35698 42478 35700 42530
rect 35644 41860 35700 42478
rect 37772 41972 37828 42702
rect 37996 42756 38052 43598
rect 39340 43650 39396 44940
rect 40236 44098 40292 46620
rect 41132 46116 41188 46126
rect 41132 46022 41188 46060
rect 41356 45778 41412 45790
rect 41356 45726 41358 45778
rect 41410 45726 41412 45778
rect 40236 44046 40238 44098
rect 40290 44046 40292 44098
rect 40236 43988 40292 44046
rect 39788 43932 40292 43988
rect 40796 45666 40852 45678
rect 40796 45614 40798 45666
rect 40850 45614 40852 45666
rect 39788 43708 39844 43932
rect 39340 43598 39342 43650
rect 39394 43598 39396 43650
rect 39340 43586 39396 43598
rect 39676 43652 39844 43708
rect 38332 43540 38388 43550
rect 38780 43540 38836 43550
rect 38332 43538 38836 43540
rect 38332 43486 38334 43538
rect 38386 43486 38782 43538
rect 38834 43486 38836 43538
rect 38332 43484 38836 43486
rect 38332 43474 38388 43484
rect 38780 43474 38836 43484
rect 39116 43316 39172 43326
rect 39676 43316 39732 43652
rect 39116 43314 39732 43316
rect 39116 43262 39118 43314
rect 39170 43262 39732 43314
rect 39116 43260 39732 43262
rect 39116 43250 39172 43260
rect 38220 42756 38276 42766
rect 37996 42754 38276 42756
rect 37996 42702 38222 42754
rect 38274 42702 38276 42754
rect 37996 42700 38276 42702
rect 38220 42690 38276 42700
rect 37772 41906 37828 41916
rect 38780 41970 38836 41982
rect 39340 41972 39396 41982
rect 38780 41918 38782 41970
rect 38834 41918 38836 41970
rect 35644 41794 35700 41804
rect 36092 41858 36148 41870
rect 36092 41806 36094 41858
rect 36146 41806 36148 41858
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 34972 41358 34974 41410
rect 35026 41358 35028 41410
rect 34972 41346 35028 41358
rect 35308 41412 35364 41422
rect 35308 41318 35364 41356
rect 36092 41412 36148 41806
rect 36092 41346 36148 41356
rect 36428 41858 36484 41870
rect 36428 41806 36430 41858
rect 36482 41806 36484 41858
rect 34972 41076 35028 41086
rect 34972 39730 35028 41020
rect 35532 41076 35588 41086
rect 35532 40982 35588 41020
rect 36092 41076 36148 41086
rect 36428 41076 36484 41806
rect 38780 41860 38836 41918
rect 38780 41794 38836 41804
rect 39228 41916 39340 41972
rect 38444 41188 38500 41198
rect 38892 41188 38948 41198
rect 39228 41188 39284 41916
rect 39340 41878 39396 41916
rect 39676 41748 39732 43260
rect 39900 43650 39956 43662
rect 39900 43598 39902 43650
rect 39954 43598 39956 43650
rect 39900 42196 39956 43598
rect 40684 42530 40740 42542
rect 40684 42478 40686 42530
rect 40738 42478 40740 42530
rect 39900 42140 40180 42196
rect 38444 41186 39284 41188
rect 38444 41134 38446 41186
rect 38498 41134 38894 41186
rect 38946 41134 39284 41186
rect 38444 41132 39284 41134
rect 39340 41692 39732 41748
rect 39788 42082 39844 42094
rect 39788 42030 39790 42082
rect 39842 42030 39844 42082
rect 38444 41122 38500 41132
rect 38892 41122 38948 41132
rect 36092 41074 36484 41076
rect 36092 41022 36094 41074
rect 36146 41022 36484 41074
rect 36092 41020 36484 41022
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34972 39678 34974 39730
rect 35026 39678 35028 39730
rect 34972 39666 35028 39678
rect 35532 39396 35588 39406
rect 34748 38894 34750 38946
rect 34802 38894 34804 38946
rect 34524 38836 34580 38846
rect 34412 38834 34580 38836
rect 34412 38782 34526 38834
rect 34578 38782 34580 38834
rect 34412 38780 34580 38782
rect 34524 38770 34580 38780
rect 34748 38668 34804 38894
rect 35084 38948 35140 38958
rect 35084 38854 35140 38892
rect 34188 38612 34244 38622
rect 34748 38612 35028 38668
rect 34188 38518 34244 38556
rect 33964 38322 34020 38332
rect 33852 38110 33854 38162
rect 33906 38110 33908 38162
rect 33852 38098 33908 38110
rect 33964 38164 34020 38174
rect 33180 36542 33182 36594
rect 33234 36542 33236 36594
rect 33180 36530 33236 36542
rect 33628 37156 33684 37166
rect 33516 36482 33572 36494
rect 33516 36430 33518 36482
rect 33570 36430 33572 36482
rect 32732 36372 32788 36382
rect 32732 36258 32788 36316
rect 32732 36206 32734 36258
rect 32786 36206 32788 36258
rect 32732 36194 32788 36206
rect 33292 35476 33348 35486
rect 33292 35474 33460 35476
rect 33292 35422 33294 35474
rect 33346 35422 33460 35474
rect 33292 35420 33460 35422
rect 33292 35410 33348 35420
rect 32620 34974 32622 35026
rect 32674 34974 32676 35026
rect 32284 34130 32340 34142
rect 32284 34078 32286 34130
rect 32338 34078 32340 34130
rect 32284 34020 32340 34078
rect 32508 34130 32564 34142
rect 32508 34078 32510 34130
rect 32562 34078 32564 34130
rect 32396 34020 32452 34030
rect 32284 33964 32396 34020
rect 32396 33954 32452 33964
rect 32508 33684 32564 34078
rect 32508 33618 32564 33628
rect 32396 33124 32452 33134
rect 32172 32834 32228 32844
rect 32284 33068 32396 33124
rect 32060 32788 32116 32798
rect 31612 32676 31668 32686
rect 31948 32676 32004 32686
rect 31612 32674 31948 32676
rect 31612 32622 31614 32674
rect 31666 32622 31948 32674
rect 31612 32620 31948 32622
rect 31612 32610 31668 32620
rect 31948 32582 32004 32620
rect 30044 31218 30660 31220
rect 30044 31166 30046 31218
rect 30098 31166 30660 31218
rect 30044 31164 30660 31166
rect 30716 31164 30828 31220
rect 30044 31154 30100 31164
rect 30268 30994 30324 31006
rect 30268 30942 30270 30994
rect 30322 30942 30324 30994
rect 29932 30324 29988 30334
rect 29484 30322 30100 30324
rect 29484 30270 29934 30322
rect 29986 30270 30100 30322
rect 29484 30268 30100 30270
rect 29932 30258 29988 30268
rect 29372 30044 29652 30100
rect 29372 29540 29428 29550
rect 29372 29446 29428 29484
rect 29484 29316 29540 29326
rect 29484 28644 29540 29260
rect 29596 28756 29652 30044
rect 29820 28756 29876 28766
rect 29596 28700 29820 28756
rect 29484 28550 29540 28588
rect 29820 28530 29876 28700
rect 29820 28478 29822 28530
rect 29874 28478 29876 28530
rect 29820 28466 29876 28478
rect 29932 28196 29988 28206
rect 29932 28082 29988 28140
rect 29932 28030 29934 28082
rect 29986 28030 29988 28082
rect 29932 28018 29988 28030
rect 30044 27524 30100 30268
rect 30268 29876 30324 30942
rect 30716 30660 30772 31164
rect 30828 31126 30884 31164
rect 31164 31276 31332 31332
rect 31388 32228 31444 32238
rect 30156 29820 30324 29876
rect 30380 30604 30772 30660
rect 30380 30210 30436 30604
rect 30380 30158 30382 30210
rect 30434 30158 30436 30210
rect 30156 29540 30212 29820
rect 30268 29652 30324 29662
rect 30380 29652 30436 30158
rect 30268 29650 30436 29652
rect 30268 29598 30270 29650
rect 30322 29598 30436 29650
rect 30268 29596 30436 29598
rect 30940 29986 30996 29998
rect 30940 29934 30942 29986
rect 30994 29934 30996 29986
rect 30268 29586 30324 29596
rect 30156 29474 30212 29484
rect 30604 29428 30660 29438
rect 30940 29428 30996 29934
rect 30604 29426 30996 29428
rect 30604 29374 30606 29426
rect 30658 29374 30996 29426
rect 30604 29372 30996 29374
rect 30492 29316 30548 29326
rect 30156 28644 30212 28654
rect 30212 28588 30324 28644
rect 30156 28550 30212 28588
rect 30268 28082 30324 28588
rect 30268 28030 30270 28082
rect 30322 28030 30324 28082
rect 30268 28018 30324 28030
rect 30380 28420 30436 28430
rect 30044 27458 30100 27468
rect 29148 26962 29316 26964
rect 29148 26910 29150 26962
rect 29202 26910 29316 26962
rect 29148 26908 29316 26910
rect 29148 26898 29204 26908
rect 29260 26068 29316 26908
rect 29148 26012 29316 26068
rect 29484 26962 29540 26974
rect 29484 26910 29486 26962
rect 29538 26910 29540 26962
rect 29148 24948 29204 26012
rect 29372 25844 29428 25854
rect 29372 25508 29428 25788
rect 29148 24882 29204 24892
rect 29260 25506 29428 25508
rect 29260 25454 29374 25506
rect 29426 25454 29428 25506
rect 29260 25452 29428 25454
rect 29148 24724 29204 24734
rect 29148 24630 29204 24668
rect 29148 23940 29204 23950
rect 29148 23846 29204 23884
rect 29148 22258 29204 22270
rect 29148 22206 29150 22258
rect 29202 22206 29204 22258
rect 29036 20020 29092 20030
rect 29036 19926 29092 19964
rect 29148 19572 29204 22206
rect 29260 21586 29316 25452
rect 29372 25442 29428 25452
rect 29484 24836 29540 26910
rect 30044 26850 30100 26862
rect 30044 26798 30046 26850
rect 30098 26798 30100 26850
rect 30044 26516 30100 26798
rect 30044 25844 30100 26460
rect 30044 25778 30100 25788
rect 29820 25618 29876 25630
rect 29820 25566 29822 25618
rect 29874 25566 29876 25618
rect 29820 25508 29876 25566
rect 30268 25508 30324 25518
rect 29820 25442 29876 25452
rect 30044 25452 30268 25508
rect 29708 24948 29764 24958
rect 30044 24948 30100 25452
rect 30268 25414 30324 25452
rect 30380 25060 30436 28364
rect 30492 27188 30548 29260
rect 30604 28868 30660 29372
rect 31164 29316 31220 31276
rect 31388 31220 31444 32172
rect 32060 31892 32116 32732
rect 32060 31798 32116 31836
rect 32284 32116 32340 33068
rect 32396 33030 32452 33068
rect 32620 32788 32676 34974
rect 33292 34244 33348 34254
rect 33292 33908 33348 34188
rect 33404 34130 33460 35420
rect 33516 34244 33572 36430
rect 33628 35698 33684 37100
rect 33628 35646 33630 35698
rect 33682 35646 33684 35698
rect 33628 35634 33684 35646
rect 33740 36370 33796 36382
rect 33740 36318 33742 36370
rect 33794 36318 33796 36370
rect 33740 35476 33796 36318
rect 33740 35410 33796 35420
rect 33852 35812 33908 35822
rect 33852 35364 33908 35756
rect 33852 35298 33908 35308
rect 33852 34356 33908 34366
rect 33964 34356 34020 38108
rect 34300 37828 34356 37838
rect 34300 37156 34356 37772
rect 34524 37156 34580 37166
rect 34300 37154 34580 37156
rect 34300 37102 34526 37154
rect 34578 37102 34580 37154
rect 34300 37100 34580 37102
rect 34412 36482 34468 36494
rect 34412 36430 34414 36482
rect 34466 36430 34468 36482
rect 34076 36372 34132 36382
rect 34076 36278 34132 36316
rect 34188 34692 34244 34702
rect 34188 34356 34244 34636
rect 33852 34354 34020 34356
rect 33852 34302 33854 34354
rect 33906 34302 34020 34354
rect 33852 34300 34020 34302
rect 34076 34354 34244 34356
rect 34076 34302 34190 34354
rect 34242 34302 34244 34354
rect 34076 34300 34244 34302
rect 33852 34290 33908 34300
rect 33628 34244 33684 34254
rect 33516 34242 33796 34244
rect 33516 34190 33630 34242
rect 33682 34190 33796 34242
rect 33516 34188 33796 34190
rect 33628 34178 33684 34188
rect 33404 34078 33406 34130
rect 33458 34078 33460 34130
rect 33404 34066 33460 34078
rect 33516 34020 33572 34030
rect 33516 33926 33572 33964
rect 33292 33852 33460 33908
rect 33180 33684 33236 33694
rect 32732 33346 32788 33358
rect 32732 33294 32734 33346
rect 32786 33294 32788 33346
rect 32732 33124 32788 33294
rect 32844 33236 32900 33246
rect 32844 33142 32900 33180
rect 32732 33058 32788 33068
rect 32956 33122 33012 33134
rect 32956 33070 32958 33122
rect 33010 33070 33012 33122
rect 32284 31668 32340 32060
rect 32060 31612 32340 31668
rect 32396 32732 32676 32788
rect 32396 32452 32452 32732
rect 32956 32676 33012 33070
rect 32620 32620 33012 32676
rect 31500 31556 31556 31566
rect 31500 31462 31556 31500
rect 31164 29250 31220 29260
rect 31276 31164 31444 31220
rect 31724 31220 31780 31230
rect 31276 30882 31332 31164
rect 31724 31126 31780 31164
rect 31276 30830 31278 30882
rect 31330 30830 31332 30882
rect 30604 28802 30660 28812
rect 30716 29092 30772 29102
rect 30716 28754 30772 29036
rect 30716 28702 30718 28754
rect 30770 28702 30772 28754
rect 30716 28690 30772 28702
rect 31164 28420 31220 28430
rect 31276 28420 31332 30830
rect 31948 30212 32004 30222
rect 31836 29764 31892 29774
rect 31836 29540 31892 29708
rect 31612 29538 31892 29540
rect 31612 29486 31838 29538
rect 31890 29486 31892 29538
rect 31612 29484 31892 29486
rect 31388 29428 31444 29438
rect 31388 29426 31556 29428
rect 31388 29374 31390 29426
rect 31442 29374 31556 29426
rect 31388 29372 31556 29374
rect 31388 29362 31444 29372
rect 31220 28364 31332 28420
rect 31500 28756 31556 29372
rect 31164 28354 31220 28364
rect 30604 27972 30660 27982
rect 30604 27878 30660 27916
rect 31388 27860 31444 27870
rect 31164 27858 31444 27860
rect 31164 27806 31390 27858
rect 31442 27806 31444 27858
rect 31164 27804 31444 27806
rect 30940 27746 30996 27758
rect 30940 27694 30942 27746
rect 30994 27694 30996 27746
rect 30940 27636 30996 27694
rect 30940 27570 30996 27580
rect 30940 27300 30996 27310
rect 30492 27186 30660 27188
rect 30492 27134 30494 27186
rect 30546 27134 30660 27186
rect 30492 27132 30660 27134
rect 30492 27122 30548 27132
rect 29708 24946 30100 24948
rect 29708 24894 29710 24946
rect 29762 24894 30100 24946
rect 29708 24892 30100 24894
rect 29708 24882 29764 24892
rect 29372 24780 29540 24836
rect 30044 24834 30100 24892
rect 30044 24782 30046 24834
rect 30098 24782 30100 24834
rect 29372 23044 29428 24780
rect 30044 24770 30100 24782
rect 30268 25004 30436 25060
rect 29708 24724 29764 24734
rect 29596 24276 29652 24286
rect 29596 23940 29652 24220
rect 29372 22978 29428 22988
rect 29484 23938 29652 23940
rect 29484 23886 29598 23938
rect 29650 23886 29652 23938
rect 29484 23884 29652 23886
rect 29260 21534 29262 21586
rect 29314 21534 29316 21586
rect 29260 20916 29316 21534
rect 29372 22484 29428 22494
rect 29372 21364 29428 22428
rect 29484 22370 29540 23884
rect 29596 23874 29652 23884
rect 29484 22318 29486 22370
rect 29538 22318 29540 22370
rect 29484 22306 29540 22318
rect 29708 22484 29764 24668
rect 30156 24610 30212 24622
rect 30156 24558 30158 24610
rect 30210 24558 30212 24610
rect 30044 24276 30100 24286
rect 30044 23826 30100 24220
rect 30044 23774 30046 23826
rect 30098 23774 30100 23826
rect 30044 23762 30100 23774
rect 30044 23380 30100 23390
rect 29708 22370 29764 22428
rect 29708 22318 29710 22370
rect 29762 22318 29764 22370
rect 29708 22306 29764 22318
rect 29932 23324 30044 23380
rect 29596 22260 29652 22270
rect 29596 22166 29652 22204
rect 29708 21700 29764 21710
rect 29708 21606 29764 21644
rect 29596 21588 29652 21598
rect 29596 21494 29652 21532
rect 29820 21476 29876 21486
rect 29708 21364 29764 21374
rect 29372 21308 29652 21364
rect 29260 20850 29316 20860
rect 29372 20132 29428 20142
rect 29260 20018 29316 20030
rect 29260 19966 29262 20018
rect 29314 19966 29316 20018
rect 29260 19908 29316 19966
rect 29260 19842 29316 19852
rect 29148 19516 29316 19572
rect 28924 19394 28980 19404
rect 28588 19348 28644 19358
rect 28588 19254 28644 19292
rect 29148 19234 29204 19246
rect 29148 19182 29150 19234
rect 29202 19182 29204 19234
rect 28700 18788 28756 18798
rect 29148 18788 29204 19182
rect 29260 18900 29316 19516
rect 29372 19348 29428 20076
rect 29372 19122 29428 19292
rect 29372 19070 29374 19122
rect 29426 19070 29428 19122
rect 29372 19058 29428 19070
rect 29484 20020 29540 20030
rect 29260 18844 29428 18900
rect 28756 18732 29204 18788
rect 28588 18564 28644 18574
rect 28700 18564 28756 18732
rect 29148 18676 29204 18732
rect 29260 18676 29316 18686
rect 29148 18674 29316 18676
rect 29148 18622 29262 18674
rect 29314 18622 29316 18674
rect 29148 18620 29316 18622
rect 29260 18610 29316 18620
rect 28588 18562 28756 18564
rect 28588 18510 28590 18562
rect 28642 18510 28756 18562
rect 28588 18508 28756 18510
rect 29036 18564 29092 18574
rect 28588 18498 28644 18508
rect 29036 18470 29092 18508
rect 28252 18274 28308 18284
rect 28364 18284 28532 18340
rect 28812 18450 28868 18462
rect 28812 18398 28814 18450
rect 28866 18398 28868 18450
rect 28252 17668 28308 17678
rect 27916 17666 28308 17668
rect 27916 17614 28254 17666
rect 28306 17614 28308 17666
rect 27916 17612 28308 17614
rect 28252 17602 28308 17612
rect 27692 17556 27748 17566
rect 27692 17462 27748 17500
rect 27020 17378 27076 17388
rect 27468 17444 27524 17454
rect 27468 17350 27524 17388
rect 27692 17276 28308 17332
rect 27692 17220 27748 17276
rect 27468 17164 27748 17220
rect 27356 17108 27412 17118
rect 27020 17106 27412 17108
rect 27020 17054 27358 17106
rect 27410 17054 27412 17106
rect 27020 17052 27412 17054
rect 27020 16100 27076 17052
rect 27356 17042 27412 17052
rect 27468 16994 27524 17164
rect 28252 17106 28308 17276
rect 28252 17054 28254 17106
rect 28306 17054 28308 17106
rect 28252 17042 28308 17054
rect 27468 16942 27470 16994
rect 27522 16942 27524 16994
rect 27468 16930 27524 16942
rect 27916 16994 27972 17006
rect 27916 16942 27918 16994
rect 27970 16942 27972 16994
rect 27356 16884 27412 16894
rect 27244 16772 27300 16782
rect 27132 16716 27244 16772
rect 27132 16322 27188 16716
rect 27244 16706 27300 16716
rect 27356 16658 27412 16828
rect 27356 16606 27358 16658
rect 27410 16606 27412 16658
rect 27356 16594 27412 16606
rect 27692 16882 27748 16894
rect 27692 16830 27694 16882
rect 27746 16830 27748 16882
rect 27132 16270 27134 16322
rect 27186 16270 27188 16322
rect 27132 16258 27188 16270
rect 27692 16100 27748 16830
rect 27916 16212 27972 16942
rect 28028 16884 28084 16894
rect 28364 16884 28420 18284
rect 28700 18228 28756 18238
rect 28476 18226 28756 18228
rect 28476 18174 28702 18226
rect 28754 18174 28756 18226
rect 28476 18172 28756 18174
rect 28476 17554 28532 18172
rect 28700 18162 28756 18172
rect 28812 17892 28868 18398
rect 29372 18228 29428 18844
rect 29484 18674 29540 19964
rect 29596 19908 29652 21308
rect 29708 21270 29764 21308
rect 29820 20802 29876 21420
rect 29820 20750 29822 20802
rect 29874 20750 29876 20802
rect 29820 20738 29876 20750
rect 29932 20580 29988 23324
rect 30044 23314 30100 23324
rect 30156 23266 30212 24558
rect 30156 23214 30158 23266
rect 30210 23214 30212 23266
rect 30156 23202 30212 23214
rect 30268 23154 30324 25004
rect 30380 24722 30436 24734
rect 30380 24670 30382 24722
rect 30434 24670 30436 24722
rect 30380 24388 30436 24670
rect 30380 24322 30436 24332
rect 30492 24722 30548 24734
rect 30492 24670 30494 24722
rect 30546 24670 30548 24722
rect 30492 24276 30548 24670
rect 30492 24210 30548 24220
rect 30268 23102 30270 23154
rect 30322 23102 30324 23154
rect 30268 23090 30324 23102
rect 30380 23826 30436 23838
rect 30380 23774 30382 23826
rect 30434 23774 30436 23826
rect 30044 22484 30100 22494
rect 30100 22428 30212 22484
rect 30044 22418 30100 22428
rect 30156 22370 30212 22428
rect 30156 22318 30158 22370
rect 30210 22318 30212 22370
rect 30156 22306 30212 22318
rect 30380 22372 30436 23774
rect 30492 23268 30548 23278
rect 30604 23268 30660 27132
rect 30828 27074 30884 27086
rect 30828 27022 30830 27074
rect 30882 27022 30884 27074
rect 30828 26852 30884 27022
rect 30828 26786 30884 26796
rect 30828 26516 30884 26526
rect 30940 26516 30996 27244
rect 30828 26514 30996 26516
rect 30828 26462 30830 26514
rect 30882 26462 30996 26514
rect 30828 26460 30996 26462
rect 31164 26852 31220 27804
rect 31388 27794 31444 27804
rect 31276 27076 31332 27114
rect 31276 27010 31332 27020
rect 31500 26908 31556 28700
rect 31612 28530 31668 29484
rect 31836 29474 31892 29484
rect 31612 28478 31614 28530
rect 31666 28478 31668 28530
rect 31612 28466 31668 28478
rect 31836 29092 31892 29102
rect 31724 28418 31780 28430
rect 31724 28366 31726 28418
rect 31778 28366 31780 28418
rect 30828 26450 30884 26460
rect 31164 26290 31220 26796
rect 31164 26238 31166 26290
rect 31218 26238 31220 26290
rect 30828 25844 30884 25854
rect 30828 25620 30884 25788
rect 30828 25618 31108 25620
rect 30828 25566 30830 25618
rect 30882 25566 31108 25618
rect 30828 25564 31108 25566
rect 30828 25554 30884 25564
rect 31052 24946 31108 25564
rect 31164 25284 31220 26238
rect 31276 26852 31556 26908
rect 31612 26962 31668 26974
rect 31612 26910 31614 26962
rect 31666 26910 31668 26962
rect 31276 25394 31332 26852
rect 31500 26402 31556 26414
rect 31500 26350 31502 26402
rect 31554 26350 31556 26402
rect 31500 25730 31556 26350
rect 31500 25678 31502 25730
rect 31554 25678 31556 25730
rect 31500 25508 31556 25678
rect 31500 25442 31556 25452
rect 31276 25342 31278 25394
rect 31330 25342 31332 25394
rect 31276 25330 31332 25342
rect 31612 25396 31668 26910
rect 31724 26740 31780 28366
rect 31836 27188 31892 29036
rect 31948 28084 32004 30156
rect 31948 27990 32004 28028
rect 32060 27636 32116 31612
rect 32172 30882 32228 30894
rect 32172 30830 32174 30882
rect 32226 30830 32228 30882
rect 32172 28644 32228 30830
rect 32284 30212 32340 30222
rect 32396 30212 32452 32396
rect 32508 32450 32564 32462
rect 32508 32398 32510 32450
rect 32562 32398 32564 32450
rect 32508 31780 32564 32398
rect 32508 30884 32564 31724
rect 32620 31778 32676 32620
rect 32620 31726 32622 31778
rect 32674 31726 32676 31778
rect 32620 31714 32676 31726
rect 32956 32452 33012 32462
rect 32956 31778 33012 32396
rect 32956 31726 32958 31778
rect 33010 31726 33012 31778
rect 32956 31714 33012 31726
rect 33180 31666 33236 33628
rect 33292 33572 33348 33582
rect 33292 33346 33348 33516
rect 33292 33294 33294 33346
rect 33346 33294 33348 33346
rect 33292 33282 33348 33294
rect 33404 32674 33460 33852
rect 33404 32622 33406 32674
rect 33458 32622 33460 32674
rect 33404 32610 33460 32622
rect 33740 32674 33796 34188
rect 33964 33460 34020 33470
rect 34076 33460 34132 34300
rect 34188 34290 34244 34300
rect 34412 34244 34468 36430
rect 34524 35700 34580 37100
rect 34524 35698 34692 35700
rect 34524 35646 34526 35698
rect 34578 35646 34692 35698
rect 34524 35644 34692 35646
rect 34524 35634 34580 35644
rect 34524 35364 34580 35374
rect 34524 35026 34580 35308
rect 34524 34974 34526 35026
rect 34578 34974 34580 35026
rect 34524 34962 34580 34974
rect 34636 34356 34692 35644
rect 34972 34580 35028 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35420 38052 35476 38062
rect 35532 38052 35588 39340
rect 36092 38948 36148 41020
rect 36092 38882 36148 38892
rect 37100 39618 37156 39630
rect 37100 39566 37102 39618
rect 37154 39566 37156 39618
rect 35868 38722 35924 38734
rect 35868 38670 35870 38722
rect 35922 38670 35924 38722
rect 35868 38164 35924 38670
rect 37100 38274 37156 39566
rect 37324 39394 37380 39406
rect 37324 39342 37326 39394
rect 37378 39342 37380 39394
rect 37212 38948 37268 38958
rect 37212 38668 37268 38892
rect 37324 38836 37380 39342
rect 38220 38836 38276 38846
rect 37324 38834 38276 38836
rect 37324 38782 38222 38834
rect 38274 38782 38276 38834
rect 37324 38780 38276 38782
rect 38220 38770 38276 38780
rect 39004 38836 39060 41132
rect 39228 40964 39284 40974
rect 39116 40908 39228 40964
rect 39116 40626 39172 40908
rect 39228 40898 39284 40908
rect 39116 40574 39118 40626
rect 39170 40574 39172 40626
rect 39116 40562 39172 40574
rect 39004 38742 39060 38780
rect 39228 38834 39284 38846
rect 39228 38782 39230 38834
rect 39282 38782 39284 38834
rect 39228 38668 39284 38782
rect 37212 38612 37492 38668
rect 37100 38222 37102 38274
rect 37154 38222 37156 38274
rect 37100 38210 37156 38222
rect 37436 38274 37492 38612
rect 37436 38222 37438 38274
rect 37490 38222 37492 38274
rect 37436 38210 37492 38222
rect 38780 38612 39284 38668
rect 38780 38274 38836 38612
rect 38780 38222 38782 38274
rect 38834 38222 38836 38274
rect 38780 38210 38836 38222
rect 35868 38098 35924 38108
rect 37996 38164 38052 38174
rect 35420 38050 35588 38052
rect 35420 37998 35422 38050
rect 35474 37998 35588 38050
rect 35420 37996 35588 37998
rect 35420 37986 35476 37996
rect 35868 37940 35924 37950
rect 35868 37846 35924 37884
rect 37660 37940 37716 37950
rect 37660 37846 37716 37884
rect 37996 37938 38052 38108
rect 39116 38052 39172 38062
rect 39116 37958 39172 37996
rect 37996 37886 37998 37938
rect 38050 37886 38052 37938
rect 37996 37874 38052 37886
rect 36988 37604 37044 37614
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35308 36482 35364 36494
rect 35308 36430 35310 36482
rect 35362 36430 35364 36482
rect 35084 36258 35140 36270
rect 35084 36206 35086 36258
rect 35138 36206 35140 36258
rect 35084 35698 35140 36206
rect 35084 35646 35086 35698
rect 35138 35646 35140 35698
rect 35084 35634 35140 35646
rect 35308 35476 35364 36430
rect 35084 35420 35364 35476
rect 36092 35588 36148 35598
rect 35084 35140 35140 35420
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 35140 35252 35150
rect 35084 35138 35252 35140
rect 35084 35086 35198 35138
rect 35250 35086 35252 35138
rect 35084 35084 35252 35086
rect 35196 35074 35252 35084
rect 35532 34916 35588 34926
rect 35532 34822 35588 34860
rect 36092 34804 36148 35532
rect 36092 34710 36148 34748
rect 36204 34914 36260 34926
rect 36204 34862 36206 34914
rect 36258 34862 36260 34914
rect 34972 34524 35252 34580
rect 35084 34356 35140 34366
rect 34636 34354 35140 34356
rect 34636 34302 35086 34354
rect 35138 34302 35140 34354
rect 34636 34300 35140 34302
rect 35084 34290 35140 34300
rect 34524 34244 34580 34254
rect 34412 34188 34524 34244
rect 34524 34020 34580 34188
rect 34524 33954 34580 33964
rect 34748 34132 34804 34142
rect 34748 33570 34804 34076
rect 35196 33908 35252 34524
rect 34748 33518 34750 33570
rect 34802 33518 34804 33570
rect 34748 33506 34804 33518
rect 35084 33852 35252 33908
rect 35868 34242 35924 34254
rect 35868 34190 35870 34242
rect 35922 34190 35924 34242
rect 35868 34132 35924 34190
rect 36204 34244 36260 34862
rect 36204 34150 36260 34188
rect 35084 33572 35140 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35084 33516 35364 33572
rect 33964 33458 34132 33460
rect 33964 33406 33966 33458
rect 34018 33406 34132 33458
rect 33964 33404 34132 33406
rect 33964 33394 34020 33404
rect 35084 33348 35140 33358
rect 35084 33254 35140 33292
rect 35196 33124 35252 33516
rect 35308 33234 35364 33516
rect 35868 33236 35924 34076
rect 36428 33908 36484 33918
rect 35308 33182 35310 33234
rect 35362 33182 35364 33234
rect 35308 33170 35364 33182
rect 35420 33234 35924 33236
rect 35420 33182 35870 33234
rect 35922 33182 35924 33234
rect 35420 33180 35924 33182
rect 33740 32622 33742 32674
rect 33794 32622 33796 32674
rect 33516 32562 33572 32574
rect 33516 32510 33518 32562
rect 33570 32510 33572 32562
rect 33516 32002 33572 32510
rect 33628 32452 33684 32462
rect 33628 32358 33684 32396
rect 33740 32228 33796 32622
rect 35084 33068 35252 33124
rect 33964 32564 34020 32574
rect 33964 32470 34020 32508
rect 33740 32162 33796 32172
rect 33516 31950 33518 32002
rect 33570 31950 33572 32002
rect 33516 31938 33572 31950
rect 33180 31614 33182 31666
rect 33234 31614 33236 31666
rect 32844 31556 32900 31566
rect 33180 31556 33236 31614
rect 33852 31778 33908 31790
rect 33852 31726 33854 31778
rect 33906 31726 33908 31778
rect 33628 31556 33684 31566
rect 33180 31500 33572 31556
rect 32844 31462 32900 31500
rect 33180 30884 33236 30894
rect 32508 30882 33348 30884
rect 32508 30830 33182 30882
rect 33234 30830 33348 30882
rect 32508 30828 33348 30830
rect 33180 30818 33236 30828
rect 32340 30156 32452 30212
rect 32284 30118 32340 30156
rect 32956 30098 33012 30110
rect 32956 30046 32958 30098
rect 33010 30046 33012 30098
rect 32508 29314 32564 29326
rect 32508 29262 32510 29314
rect 32562 29262 32564 29314
rect 32508 29092 32564 29262
rect 32956 29316 33012 30046
rect 33180 29538 33236 29550
rect 33180 29486 33182 29538
rect 33234 29486 33236 29538
rect 33068 29316 33124 29326
rect 32956 29314 33124 29316
rect 32956 29262 33070 29314
rect 33122 29262 33124 29314
rect 32956 29260 33124 29262
rect 33068 29250 33124 29260
rect 33180 29092 33236 29486
rect 33292 29428 33348 30828
rect 33292 29362 33348 29372
rect 33404 29316 33460 29326
rect 33404 29222 33460 29260
rect 33516 29092 33572 31500
rect 33684 31500 33796 31556
rect 33628 31490 33684 31500
rect 32508 29036 33236 29092
rect 32620 28644 32676 28654
rect 33180 28644 33236 29036
rect 32172 28588 32620 28644
rect 32620 28550 32676 28588
rect 33068 28588 33236 28644
rect 33292 29036 33572 29092
rect 33628 30884 33684 30894
rect 33628 29092 33684 30828
rect 32284 28084 32340 28094
rect 32172 27636 32228 27646
rect 32060 27580 32172 27636
rect 32172 27570 32228 27580
rect 31836 27122 31892 27132
rect 31836 26964 31892 27002
rect 31836 26898 31892 26908
rect 31724 26684 31892 26740
rect 31836 26516 31892 26684
rect 31836 26460 32004 26516
rect 31836 26290 31892 26302
rect 31836 26238 31838 26290
rect 31890 26238 31892 26290
rect 31836 25508 31892 26238
rect 31836 25414 31892 25452
rect 31612 25330 31668 25340
rect 31164 25218 31220 25228
rect 31388 25282 31444 25294
rect 31948 25284 32004 26460
rect 31388 25230 31390 25282
rect 31442 25230 31444 25282
rect 31052 24894 31054 24946
rect 31106 24894 31108 24946
rect 30940 24052 30996 24062
rect 31052 24052 31108 24894
rect 30940 24050 31108 24052
rect 30940 23998 30942 24050
rect 30994 23998 31108 24050
rect 30940 23996 31108 23998
rect 31164 24500 31220 24510
rect 30940 23986 30996 23996
rect 31164 23548 31220 24444
rect 31276 24388 31332 24398
rect 31276 24050 31332 24332
rect 31276 23998 31278 24050
rect 31330 23998 31332 24050
rect 31276 23986 31332 23998
rect 31164 23492 31332 23548
rect 30548 23212 30660 23268
rect 31052 23378 31108 23390
rect 31052 23326 31054 23378
rect 31106 23326 31108 23378
rect 30492 23202 30548 23212
rect 30716 22932 30772 22942
rect 30156 21028 30212 21038
rect 30044 20972 30156 21028
rect 30044 20802 30100 20972
rect 30156 20962 30212 20972
rect 30268 20804 30324 20814
rect 30044 20750 30046 20802
rect 30098 20750 30100 20802
rect 30044 20738 30100 20750
rect 30156 20802 30324 20804
rect 30156 20750 30270 20802
rect 30322 20750 30324 20802
rect 30156 20748 30324 20750
rect 29708 20524 29988 20580
rect 29708 20130 29764 20524
rect 30156 20356 30212 20748
rect 30268 20738 30324 20748
rect 29708 20078 29710 20130
rect 29762 20078 29764 20130
rect 29708 20066 29764 20078
rect 29820 20300 30212 20356
rect 29820 20130 29876 20300
rect 29820 20078 29822 20130
rect 29874 20078 29876 20130
rect 29820 20066 29876 20078
rect 29932 20132 29988 20142
rect 29932 20038 29988 20076
rect 30380 20130 30436 22316
rect 30380 20078 30382 20130
rect 30434 20078 30436 20130
rect 30380 20066 30436 20078
rect 30492 22930 30772 22932
rect 30492 22878 30718 22930
rect 30770 22878 30772 22930
rect 30492 22876 30772 22878
rect 30492 20802 30548 22876
rect 30716 22866 30772 22876
rect 30940 22930 30996 22942
rect 30940 22878 30942 22930
rect 30994 22878 30996 22930
rect 30604 22370 30660 22382
rect 30604 22318 30606 22370
rect 30658 22318 30660 22370
rect 30604 21812 30660 22318
rect 30716 22260 30772 22270
rect 30716 22166 30772 22204
rect 30660 21756 30772 21812
rect 30604 21746 30660 21756
rect 30492 20750 30494 20802
rect 30546 20750 30548 20802
rect 30268 20020 30324 20030
rect 30268 19926 30324 19964
rect 29596 19852 29764 19908
rect 29596 19460 29652 19470
rect 29596 19346 29652 19404
rect 29596 19294 29598 19346
rect 29650 19294 29652 19346
rect 29596 19282 29652 19294
rect 29484 18622 29486 18674
rect 29538 18622 29540 18674
rect 29484 18610 29540 18622
rect 29596 18788 29652 18798
rect 29596 18562 29652 18732
rect 29596 18510 29598 18562
rect 29650 18510 29652 18562
rect 29596 18498 29652 18510
rect 29372 18162 29428 18172
rect 29484 18452 29540 18462
rect 28812 17826 28868 17836
rect 29484 17668 29540 18396
rect 29484 17574 29540 17612
rect 28476 17502 28478 17554
rect 28530 17502 28532 17554
rect 28476 17220 28532 17502
rect 28588 17556 28644 17566
rect 29148 17556 29204 17566
rect 28588 17554 29204 17556
rect 28588 17502 28590 17554
rect 28642 17502 29150 17554
rect 29202 17502 29204 17554
rect 28588 17500 29204 17502
rect 28588 17490 28644 17500
rect 28476 17164 28756 17220
rect 28028 16790 28084 16828
rect 28140 16828 28420 16884
rect 28476 16994 28532 17006
rect 28476 16942 28478 16994
rect 28530 16942 28532 16994
rect 27916 16146 27972 16156
rect 27020 16098 27748 16100
rect 27020 16046 27022 16098
rect 27074 16046 27748 16098
rect 27020 16044 27748 16046
rect 27020 16034 27076 16044
rect 26908 15486 26910 15538
rect 26962 15486 26964 15538
rect 26908 15474 26964 15486
rect 27020 15876 27076 15886
rect 27020 15426 27076 15820
rect 27132 15874 27188 15886
rect 27804 15876 27860 15886
rect 27132 15822 27134 15874
rect 27186 15822 27188 15874
rect 27132 15652 27188 15822
rect 27132 15586 27188 15596
rect 27692 15874 27860 15876
rect 27692 15822 27806 15874
rect 27858 15822 27860 15874
rect 27692 15820 27860 15822
rect 27020 15374 27022 15426
rect 27074 15374 27076 15426
rect 27020 15362 27076 15374
rect 27244 15316 27300 15326
rect 26796 15260 26964 15316
rect 26460 14644 26516 14654
rect 26460 14642 26628 14644
rect 26460 14590 26462 14642
rect 26514 14590 26628 14642
rect 26460 14588 26628 14590
rect 26460 14578 26516 14588
rect 26460 13746 26516 13758
rect 26460 13694 26462 13746
rect 26514 13694 26516 13746
rect 26460 13524 26516 13694
rect 26460 13458 26516 13468
rect 26012 13020 26404 13076
rect 25900 12738 25956 12750
rect 25900 12686 25902 12738
rect 25954 12686 25956 12738
rect 25900 12404 25956 12686
rect 25900 12338 25956 12348
rect 25900 12180 25956 12190
rect 26012 12180 26068 13020
rect 26348 12964 26404 13020
rect 26460 12964 26516 12974
rect 26348 12962 26516 12964
rect 26348 12910 26462 12962
rect 26514 12910 26516 12962
rect 26348 12908 26516 12910
rect 26460 12898 26516 12908
rect 26124 12850 26180 12862
rect 26124 12798 26126 12850
rect 26178 12798 26180 12850
rect 26124 12740 26180 12798
rect 26572 12852 26628 14588
rect 26908 13972 26964 15260
rect 26684 13916 26964 13972
rect 26684 13858 26740 13916
rect 26684 13806 26686 13858
rect 26738 13806 26740 13858
rect 26684 13794 26740 13806
rect 26908 13076 26964 13916
rect 27132 14756 27188 14766
rect 27132 13524 27188 14700
rect 27244 13746 27300 15260
rect 27580 15204 27636 15214
rect 27468 14644 27524 14654
rect 27468 14550 27524 14588
rect 27580 14530 27636 15148
rect 27692 14756 27748 15820
rect 27804 15810 27860 15820
rect 27692 14690 27748 14700
rect 27804 15314 27860 15326
rect 27804 15262 27806 15314
rect 27858 15262 27860 15314
rect 27804 14532 27860 15262
rect 27580 14478 27582 14530
rect 27634 14478 27636 14530
rect 27580 14466 27636 14478
rect 27692 14476 27860 14532
rect 27916 14980 27972 14990
rect 27916 14530 27972 14924
rect 27916 14478 27918 14530
rect 27970 14478 27972 14530
rect 27244 13694 27246 13746
rect 27298 13694 27300 13746
rect 27244 13682 27300 13694
rect 27356 14306 27412 14318
rect 27356 14254 27358 14306
rect 27410 14254 27412 14306
rect 27132 13458 27188 13468
rect 27356 13188 27412 14254
rect 27692 13748 27748 14476
rect 27916 14466 27972 14478
rect 26908 13010 26964 13020
rect 27244 13132 27412 13188
rect 27468 13746 27748 13748
rect 27468 13694 27694 13746
rect 27746 13694 27748 13746
rect 27468 13692 27748 13694
rect 26572 12796 26740 12852
rect 26124 12404 26180 12684
rect 26236 12740 26292 12750
rect 26236 12738 26628 12740
rect 26236 12686 26238 12738
rect 26290 12686 26628 12738
rect 26236 12684 26628 12686
rect 26236 12674 26292 12684
rect 26236 12404 26292 12414
rect 26124 12402 26292 12404
rect 26124 12350 26238 12402
rect 26290 12350 26292 12402
rect 26124 12348 26292 12350
rect 25900 12178 26068 12180
rect 25900 12126 25902 12178
rect 25954 12126 26068 12178
rect 25900 12124 26068 12126
rect 25900 12114 25956 12124
rect 26236 10164 26292 12348
rect 26460 12292 26516 12302
rect 26460 11506 26516 12236
rect 26572 12178 26628 12684
rect 26572 12126 26574 12178
rect 26626 12126 26628 12178
rect 26572 12114 26628 12126
rect 26460 11454 26462 11506
rect 26514 11454 26516 11506
rect 26460 11442 26516 11454
rect 26236 10098 26292 10108
rect 26684 10052 26740 12796
rect 26796 12628 26852 12638
rect 26796 12292 26852 12572
rect 27020 12516 27076 12526
rect 27076 12460 27188 12516
rect 27020 12450 27076 12460
rect 26796 12226 26852 12236
rect 27020 12068 27076 12078
rect 26684 9986 26740 9996
rect 26908 12066 27076 12068
rect 26908 12014 27022 12066
rect 27074 12014 27076 12066
rect 26908 12012 27076 12014
rect 25788 9762 25844 9772
rect 26908 9716 26964 12012
rect 27020 12002 27076 12012
rect 27020 11508 27076 11518
rect 27132 11508 27188 12460
rect 27244 12404 27300 13132
rect 27356 12964 27412 12974
rect 27356 12870 27412 12908
rect 27356 12404 27412 12414
rect 27244 12348 27356 12404
rect 27356 12338 27412 12348
rect 27356 12180 27412 12190
rect 27020 11506 27188 11508
rect 27020 11454 27022 11506
rect 27074 11454 27188 11506
rect 27020 11452 27188 11454
rect 27244 12124 27356 12180
rect 27020 11442 27076 11452
rect 27244 11284 27300 12124
rect 27356 12114 27412 12124
rect 27468 11508 27524 13692
rect 27692 13682 27748 13692
rect 27580 13522 27636 13534
rect 27580 13470 27582 13522
rect 27634 13470 27636 13522
rect 27580 12290 27636 13470
rect 27916 13188 27972 13198
rect 27916 12962 27972 13132
rect 27916 12910 27918 12962
rect 27970 12910 27972 12962
rect 27916 12898 27972 12910
rect 28140 12964 28196 16828
rect 28476 16772 28532 16942
rect 28252 16716 28532 16772
rect 28588 16882 28644 16894
rect 28588 16830 28590 16882
rect 28642 16830 28644 16882
rect 28252 16100 28308 16716
rect 28588 16660 28644 16830
rect 28700 16884 28756 17164
rect 28700 16818 28756 16828
rect 28812 16660 28868 17500
rect 28588 16604 28868 16660
rect 28364 16212 28420 16222
rect 28364 16118 28420 16156
rect 28924 16212 28980 16222
rect 29148 16212 29204 17500
rect 29372 16212 29428 16222
rect 28980 16156 29092 16212
rect 29148 16210 29428 16212
rect 29148 16158 29374 16210
rect 29426 16158 29428 16210
rect 29148 16156 29428 16158
rect 28924 16146 28980 16156
rect 28252 15204 28308 16044
rect 28252 13970 28308 15148
rect 28588 15540 28644 15550
rect 28364 14418 28420 14430
rect 28364 14366 28366 14418
rect 28418 14366 28420 14418
rect 28364 14084 28420 14366
rect 28364 14018 28420 14028
rect 28476 14306 28532 14318
rect 28476 14254 28478 14306
rect 28530 14254 28532 14306
rect 28252 13918 28254 13970
rect 28306 13918 28308 13970
rect 28252 13906 28308 13918
rect 28476 13860 28532 14254
rect 28588 14308 28644 15484
rect 29036 14868 29092 16156
rect 29372 16146 29428 16156
rect 29484 16100 29540 16110
rect 29484 16006 29540 16044
rect 29036 14812 29316 14868
rect 28588 14242 28644 14252
rect 28700 14306 28756 14318
rect 28700 14254 28702 14306
rect 28754 14254 28756 14306
rect 28700 14084 28756 14254
rect 28700 14028 29092 14084
rect 28364 13636 28420 13646
rect 28364 13300 28420 13580
rect 28476 13524 28532 13804
rect 28588 13748 28644 13758
rect 29036 13748 29092 14028
rect 29260 13858 29316 14812
rect 29708 14196 29764 19852
rect 30492 19684 30548 20750
rect 30604 20580 30660 20590
rect 30604 20486 30660 20524
rect 30268 19628 30548 19684
rect 29708 14130 29764 14140
rect 29820 17892 29876 17902
rect 29820 14530 29876 17836
rect 29932 17778 29988 17790
rect 29932 17726 29934 17778
rect 29986 17726 29988 17778
rect 29932 17332 29988 17726
rect 29932 17266 29988 17276
rect 30044 17444 30100 17454
rect 29932 17108 29988 17118
rect 29932 17014 29988 17052
rect 30044 16994 30100 17388
rect 30044 16942 30046 16994
rect 30098 16942 30100 16994
rect 30044 16930 30100 16942
rect 29932 16660 29988 16670
rect 29932 16566 29988 16604
rect 30156 15986 30212 15998
rect 30156 15934 30158 15986
rect 30210 15934 30212 15986
rect 29820 14478 29822 14530
rect 29874 14478 29876 14530
rect 29260 13806 29262 13858
rect 29314 13806 29316 13858
rect 29148 13748 29204 13758
rect 29036 13746 29204 13748
rect 29036 13694 29150 13746
rect 29202 13694 29204 13746
rect 29036 13692 29204 13694
rect 28588 13654 28644 13692
rect 29148 13682 29204 13692
rect 28476 13468 28644 13524
rect 28364 13234 28420 13244
rect 28252 13188 28308 13198
rect 28252 13094 28308 13132
rect 28588 13186 28644 13468
rect 28588 13134 28590 13186
rect 28642 13134 28644 13186
rect 28588 13122 28644 13134
rect 29148 13300 29204 13310
rect 28140 12908 28308 12964
rect 27692 12850 27748 12862
rect 27692 12798 27694 12850
rect 27746 12798 27748 12850
rect 27692 12740 27748 12798
rect 27692 12674 27748 12684
rect 27804 12738 27860 12750
rect 27804 12686 27806 12738
rect 27858 12686 27860 12738
rect 27580 12238 27582 12290
rect 27634 12238 27636 12290
rect 27580 12226 27636 12238
rect 27692 12180 27748 12190
rect 27804 12180 27860 12686
rect 27692 12178 27860 12180
rect 27692 12126 27694 12178
rect 27746 12126 27860 12178
rect 27692 12124 27860 12126
rect 28140 12292 28196 12302
rect 27692 12114 27748 12124
rect 28140 11788 28196 12236
rect 27916 11732 27972 11742
rect 27804 11508 27860 11518
rect 27468 11506 27860 11508
rect 27468 11454 27806 11506
rect 27858 11454 27860 11506
rect 27468 11452 27860 11454
rect 27804 11396 27860 11452
rect 27804 11330 27860 11340
rect 27020 11228 27300 11284
rect 27020 10834 27076 11228
rect 27020 10782 27022 10834
rect 27074 10782 27076 10834
rect 27020 10770 27076 10782
rect 27356 10612 27412 10622
rect 27692 10612 27748 10622
rect 27132 10610 27748 10612
rect 27132 10558 27358 10610
rect 27410 10558 27694 10610
rect 27746 10558 27748 10610
rect 27132 10556 27748 10558
rect 27020 9940 27076 9950
rect 27132 9940 27188 10556
rect 27356 10546 27412 10556
rect 27692 10546 27748 10556
rect 27020 9938 27188 9940
rect 27020 9886 27022 9938
rect 27074 9886 27188 9938
rect 27020 9884 27188 9886
rect 27804 10500 27860 10510
rect 27020 9874 27076 9884
rect 26908 9650 26964 9660
rect 25676 9156 25732 9166
rect 25284 9100 25396 9156
rect 25564 9154 25732 9156
rect 25564 9102 25678 9154
rect 25730 9102 25732 9154
rect 25564 9100 25732 9102
rect 25228 9062 25284 9100
rect 25452 9042 25508 9054
rect 25452 8990 25454 9042
rect 25506 8990 25508 9042
rect 25228 8708 25284 8718
rect 25228 8148 25284 8652
rect 25228 8082 25284 8092
rect 25004 7410 25060 7420
rect 25004 6580 25060 6590
rect 25004 6486 25060 6524
rect 25228 6468 25284 6478
rect 24668 6244 24724 6254
rect 24220 6078 24222 6130
rect 24274 6078 24276 6130
rect 24220 6066 24276 6078
rect 24444 6132 24500 6142
rect 24444 6038 24500 6076
rect 24668 6130 24724 6188
rect 24668 6078 24670 6130
rect 24722 6078 24724 6130
rect 24668 6066 24724 6078
rect 23548 5966 23550 6018
rect 23602 5966 23604 6018
rect 23548 5954 23604 5966
rect 25228 6018 25284 6412
rect 25340 6356 25396 6366
rect 25340 6130 25396 6300
rect 25340 6078 25342 6130
rect 25394 6078 25396 6130
rect 25340 6066 25396 6078
rect 25452 6132 25508 8990
rect 25564 7588 25620 9100
rect 25676 9090 25732 9100
rect 27580 9044 27636 9054
rect 27580 8950 27636 8988
rect 27132 8930 27188 8942
rect 27132 8878 27134 8930
rect 27186 8878 27188 8930
rect 25788 8818 25844 8830
rect 25788 8766 25790 8818
rect 25842 8766 25844 8818
rect 25676 8372 25732 8382
rect 25676 8278 25732 8316
rect 25676 7588 25732 7598
rect 25564 7532 25676 7588
rect 25676 7474 25732 7532
rect 25676 7422 25678 7474
rect 25730 7422 25732 7474
rect 25676 7410 25732 7422
rect 25564 7252 25620 7262
rect 25564 7158 25620 7196
rect 25788 7028 25844 8766
rect 25900 8372 25956 8382
rect 25900 7362 25956 8316
rect 27132 8372 27188 8878
rect 27132 8306 27188 8316
rect 27804 8372 27860 10444
rect 27916 9826 27972 11676
rect 27916 9774 27918 9826
rect 27970 9774 27972 9826
rect 27916 9042 27972 9774
rect 27916 8990 27918 9042
rect 27970 8990 27972 9042
rect 27916 8978 27972 8990
rect 28028 11732 28196 11788
rect 28028 10610 28084 11732
rect 28028 10558 28030 10610
rect 28082 10558 28084 10610
rect 27804 8306 27860 8316
rect 27916 8372 27972 8382
rect 28028 8372 28084 10558
rect 28140 10500 28196 10510
rect 28252 10500 28308 12908
rect 28364 12738 28420 12750
rect 28364 12686 28366 12738
rect 28418 12686 28420 12738
rect 28364 12516 28420 12686
rect 28364 12450 28420 12460
rect 28196 10444 28308 10500
rect 28364 12292 28420 12302
rect 28140 10434 28196 10444
rect 28140 10052 28196 10062
rect 28196 9996 28308 10052
rect 28140 9986 28196 9996
rect 28140 9602 28196 9614
rect 28140 9550 28142 9602
rect 28194 9550 28196 9602
rect 28140 9492 28196 9550
rect 28140 9426 28196 9436
rect 28140 9156 28196 9166
rect 28140 8484 28196 9100
rect 28140 8418 28196 8428
rect 27916 8370 28084 8372
rect 27916 8318 27918 8370
rect 27970 8318 28084 8370
rect 27916 8316 28084 8318
rect 27916 8306 27972 8316
rect 28140 7588 28196 7598
rect 28252 7588 28308 9996
rect 28364 9492 28420 12236
rect 29148 12180 29204 13244
rect 29260 12962 29316 13806
rect 29820 13972 29876 14478
rect 29484 13748 29540 13758
rect 29260 12910 29262 12962
rect 29314 12910 29316 12962
rect 29260 12898 29316 12910
rect 29372 13188 29428 13198
rect 29372 12852 29428 13132
rect 29148 12086 29204 12124
rect 29260 12740 29316 12750
rect 29260 12516 29316 12684
rect 28588 11954 28644 11966
rect 28588 11902 28590 11954
rect 28642 11902 28644 11954
rect 28476 11396 28532 11406
rect 28588 11396 28644 11902
rect 28476 11394 29092 11396
rect 28476 11342 28478 11394
rect 28530 11342 29092 11394
rect 28476 11340 29092 11342
rect 28476 11330 28532 11340
rect 28476 10388 28532 10398
rect 28476 9604 28532 10332
rect 29036 10052 29092 11340
rect 29148 10052 29204 10062
rect 29036 10050 29204 10052
rect 29036 9998 29150 10050
rect 29202 9998 29204 10050
rect 29036 9996 29204 9998
rect 29148 9986 29204 9996
rect 29260 9828 29316 12460
rect 29372 11282 29428 12796
rect 29372 11230 29374 11282
rect 29426 11230 29428 11282
rect 29372 11218 29428 11230
rect 29484 10836 29540 13692
rect 29596 13074 29652 13086
rect 29596 13022 29598 13074
rect 29650 13022 29652 13074
rect 29596 12964 29652 13022
rect 29596 12898 29652 12908
rect 29820 12628 29876 13916
rect 29708 12572 29876 12628
rect 29932 15652 29988 15662
rect 29932 15314 29988 15596
rect 29932 15262 29934 15314
rect 29986 15262 29988 15314
rect 29596 12180 29652 12190
rect 29596 11394 29652 12124
rect 29596 11342 29598 11394
rect 29650 11342 29652 11394
rect 29596 11330 29652 11342
rect 29036 9772 29316 9828
rect 29372 10780 29540 10836
rect 29372 10052 29428 10780
rect 29484 10612 29540 10622
rect 29484 10518 29540 10556
rect 29484 10052 29540 10062
rect 29372 10050 29540 10052
rect 29372 9998 29486 10050
rect 29538 9998 29540 10050
rect 29372 9996 29540 9998
rect 28588 9604 28644 9614
rect 28476 9602 28644 9604
rect 28476 9550 28590 9602
rect 28642 9550 28644 9602
rect 28476 9548 28644 9550
rect 28364 9426 28420 9436
rect 28476 9042 28532 9054
rect 28476 8990 28478 9042
rect 28530 8990 28532 9042
rect 28476 8820 28532 8990
rect 28476 8754 28532 8764
rect 28476 8484 28532 8494
rect 28588 8484 28644 9548
rect 28532 8428 28644 8484
rect 28812 9042 28868 9054
rect 28812 8990 28814 9042
rect 28866 8990 28868 9042
rect 28476 8370 28532 8428
rect 28476 8318 28478 8370
rect 28530 8318 28532 8370
rect 28476 8306 28532 8318
rect 28812 8036 28868 8990
rect 28812 7970 28868 7980
rect 28140 7586 28308 7588
rect 28140 7534 28142 7586
rect 28194 7534 28308 7586
rect 28140 7532 28308 7534
rect 25900 7310 25902 7362
rect 25954 7310 25956 7362
rect 25900 7298 25956 7310
rect 26460 7476 26516 7486
rect 25788 6962 25844 6972
rect 26012 6692 26068 6702
rect 25452 6066 25508 6076
rect 25564 6690 26068 6692
rect 25564 6638 26014 6690
rect 26066 6638 26068 6690
rect 25564 6636 26068 6638
rect 25564 6130 25620 6636
rect 26012 6626 26068 6636
rect 26124 6692 26180 6702
rect 26124 6466 26180 6636
rect 26460 6692 26516 7420
rect 26908 7476 26964 7486
rect 26908 7382 26964 7420
rect 27468 7476 27524 7486
rect 27692 7476 27748 7486
rect 27468 7382 27524 7420
rect 27580 7474 27748 7476
rect 27580 7422 27694 7474
rect 27746 7422 27748 7474
rect 27580 7420 27748 7422
rect 26908 7028 26964 7038
rect 26460 6626 26516 6636
rect 26796 6692 26852 6702
rect 26124 6414 26126 6466
rect 26178 6414 26180 6466
rect 26124 6402 26180 6414
rect 26348 6580 26404 6590
rect 25564 6078 25566 6130
rect 25618 6078 25620 6130
rect 25564 6066 25620 6078
rect 26348 6130 26404 6524
rect 26348 6078 26350 6130
rect 26402 6078 26404 6130
rect 26348 6066 26404 6078
rect 26572 6578 26628 6590
rect 26572 6526 26574 6578
rect 26626 6526 26628 6578
rect 25228 5966 25230 6018
rect 25282 5966 25284 6018
rect 25228 5954 25284 5966
rect 23436 5854 23438 5906
rect 23490 5854 23492 5906
rect 23436 5842 23492 5854
rect 25788 5908 25844 5918
rect 25788 5814 25844 5852
rect 24556 5796 24612 5806
rect 24556 5702 24612 5740
rect 26012 5796 26068 5806
rect 26572 5796 26628 6526
rect 26796 6578 26852 6636
rect 26796 6526 26798 6578
rect 26850 6526 26852 6578
rect 26796 6514 26852 6526
rect 26908 5906 26964 6972
rect 27580 6580 27636 7420
rect 27692 7410 27748 7420
rect 27916 7362 27972 7374
rect 27916 7310 27918 7362
rect 27970 7310 27972 7362
rect 27244 6524 27636 6580
rect 27804 6580 27860 6590
rect 27244 6130 27300 6524
rect 27804 6486 27860 6524
rect 27244 6078 27246 6130
rect 27298 6078 27300 6130
rect 27244 6066 27300 6078
rect 27916 6020 27972 7310
rect 28140 6690 28196 7532
rect 28140 6638 28142 6690
rect 28194 6638 28196 6690
rect 28140 6626 28196 6638
rect 28364 7474 28420 7486
rect 28364 7422 28366 7474
rect 28418 7422 28420 7474
rect 28364 6692 28420 7422
rect 29036 7474 29092 9772
rect 29372 9380 29428 9996
rect 29484 9986 29540 9996
rect 29708 9938 29764 12572
rect 29932 12178 29988 15262
rect 30156 13748 30212 15934
rect 30156 13682 30212 13692
rect 30268 13074 30324 19628
rect 30716 18900 30772 21756
rect 30828 21364 30884 21374
rect 30828 20802 30884 21308
rect 30940 21028 30996 22878
rect 31052 22708 31108 23326
rect 31052 22642 31108 22652
rect 30940 20916 30996 20972
rect 31052 20916 31108 20926
rect 30940 20914 31108 20916
rect 30940 20862 31054 20914
rect 31106 20862 31108 20914
rect 30940 20860 31108 20862
rect 31276 20916 31332 23492
rect 31388 23380 31444 25230
rect 31836 25228 32004 25284
rect 32172 25284 32228 25294
rect 31388 23314 31444 23324
rect 31612 24610 31668 24622
rect 31612 24558 31614 24610
rect 31666 24558 31668 24610
rect 31500 22370 31556 22382
rect 31500 22318 31502 22370
rect 31554 22318 31556 22370
rect 31500 21588 31556 22318
rect 31500 21522 31556 21532
rect 31276 20860 31444 20916
rect 31052 20850 31108 20860
rect 30828 20750 30830 20802
rect 30882 20750 30884 20802
rect 30828 20738 30884 20750
rect 31164 20802 31220 20814
rect 31164 20750 31166 20802
rect 31218 20750 31220 20802
rect 30940 20692 30996 20702
rect 30996 20636 31108 20692
rect 30940 20626 30996 20636
rect 30828 19236 30884 19246
rect 30828 19142 30884 19180
rect 30380 18844 30772 18900
rect 30380 16994 30436 18844
rect 31052 18788 31108 20636
rect 31164 20244 31220 20750
rect 31164 20178 31220 20188
rect 31276 20692 31332 20702
rect 30492 18732 31108 18788
rect 31164 19796 31220 19806
rect 30492 18450 30548 18732
rect 30492 18398 30494 18450
rect 30546 18398 30548 18450
rect 30492 18386 30548 18398
rect 30604 17666 30660 17678
rect 30604 17614 30606 17666
rect 30658 17614 30660 17666
rect 30604 17108 30660 17614
rect 30828 17666 30884 18732
rect 30940 18564 30996 18574
rect 30940 18452 30996 18508
rect 31164 18452 31220 19740
rect 30940 18450 31220 18452
rect 30940 18398 30942 18450
rect 30994 18398 31220 18450
rect 30940 18396 31220 18398
rect 30940 18386 30996 18396
rect 31276 18340 31332 20636
rect 31164 18338 31332 18340
rect 31164 18286 31278 18338
rect 31330 18286 31332 18338
rect 31164 18284 31332 18286
rect 30828 17614 30830 17666
rect 30882 17614 30884 17666
rect 30828 17602 30884 17614
rect 31052 18228 31108 18238
rect 31052 17666 31108 18172
rect 31052 17614 31054 17666
rect 31106 17614 31108 17666
rect 31052 17602 31108 17614
rect 30940 17444 30996 17454
rect 30940 17350 30996 17388
rect 31164 17444 31220 18284
rect 31276 18274 31332 18284
rect 30604 17052 31108 17108
rect 30380 16942 30382 16994
rect 30434 16942 30436 16994
rect 30380 14756 30436 16942
rect 30940 16882 30996 16894
rect 30940 16830 30942 16882
rect 30994 16830 30996 16882
rect 30940 16772 30996 16830
rect 30492 16660 30548 16670
rect 30492 16210 30548 16604
rect 30492 16158 30494 16210
rect 30546 16158 30548 16210
rect 30492 16146 30548 16158
rect 30604 15874 30660 15886
rect 30604 15822 30606 15874
rect 30658 15822 30660 15874
rect 30492 15314 30548 15326
rect 30492 15262 30494 15314
rect 30546 15262 30548 15314
rect 30492 14980 30548 15262
rect 30604 15316 30660 15822
rect 30940 15764 30996 16716
rect 30940 15698 30996 15708
rect 30940 15316 30996 15326
rect 30604 15314 30996 15316
rect 30604 15262 30942 15314
rect 30994 15262 30996 15314
rect 30604 15260 30996 15262
rect 30940 15250 30996 15260
rect 31052 15148 31108 17052
rect 31164 16882 31220 17388
rect 31164 16830 31166 16882
rect 31218 16830 31220 16882
rect 31164 15988 31220 16830
rect 31276 17442 31332 17454
rect 31276 17390 31278 17442
rect 31330 17390 31332 17442
rect 31276 16772 31332 17390
rect 31276 16706 31332 16716
rect 31388 16996 31444 20860
rect 31500 20692 31556 20702
rect 31500 20598 31556 20636
rect 31612 17892 31668 24558
rect 31836 24612 31892 25228
rect 32172 25190 32228 25228
rect 32284 24724 32340 28028
rect 32620 27186 32676 27198
rect 32620 27134 32622 27186
rect 32674 27134 32676 27186
rect 32508 27076 32564 27086
rect 32396 26516 32452 26526
rect 32508 26516 32564 27020
rect 32396 26514 32564 26516
rect 32396 26462 32398 26514
rect 32450 26462 32564 26514
rect 32396 26460 32564 26462
rect 32396 26450 32452 26460
rect 32620 25508 32676 27134
rect 32956 27188 33012 27198
rect 32956 27074 33012 27132
rect 32956 27022 32958 27074
rect 33010 27022 33012 27074
rect 32956 27010 33012 27022
rect 33068 26908 33124 28588
rect 33180 27746 33236 27758
rect 33180 27694 33182 27746
rect 33234 27694 33236 27746
rect 33180 27076 33236 27694
rect 33180 27010 33236 27020
rect 33068 26852 33236 26908
rect 33180 26404 33236 26852
rect 33180 26338 33236 26348
rect 32508 25452 32676 25508
rect 33068 26066 33124 26078
rect 33068 26014 33070 26066
rect 33122 26014 33124 26066
rect 32284 24630 32340 24668
rect 32396 25282 32452 25294
rect 32396 25230 32398 25282
rect 32450 25230 32452 25282
rect 31836 24546 31892 24556
rect 31948 24498 32004 24510
rect 31948 24446 31950 24498
rect 32002 24446 32004 24498
rect 31948 24164 32004 24446
rect 31948 24098 32004 24108
rect 32396 24052 32452 25230
rect 32508 25060 32564 25452
rect 32732 25396 32788 25406
rect 33068 25396 33124 26014
rect 32788 25340 33124 25396
rect 32732 25302 32788 25340
rect 32620 25284 32676 25294
rect 32620 25190 32676 25228
rect 32508 25004 32676 25060
rect 32508 24610 32564 24622
rect 32508 24558 32510 24610
rect 32562 24558 32564 24610
rect 32508 24500 32564 24558
rect 32508 24434 32564 24444
rect 32620 24276 32676 25004
rect 32284 23996 32452 24052
rect 32508 24220 32676 24276
rect 32172 23716 32228 23726
rect 32172 23622 32228 23660
rect 31724 23266 31780 23278
rect 31724 23214 31726 23266
rect 31778 23214 31780 23266
rect 31724 23044 31780 23214
rect 31724 22978 31780 22988
rect 31836 23154 31892 23166
rect 31836 23102 31838 23154
rect 31890 23102 31892 23154
rect 31836 22932 31892 23102
rect 31836 22866 31892 22876
rect 31948 23042 32004 23054
rect 31948 22990 31950 23042
rect 32002 22990 32004 23042
rect 31836 22708 31892 22718
rect 31836 22370 31892 22652
rect 31836 22318 31838 22370
rect 31890 22318 31892 22370
rect 31836 22306 31892 22318
rect 31724 22036 31780 22046
rect 31724 21810 31780 21980
rect 31724 21758 31726 21810
rect 31778 21758 31780 21810
rect 31724 21746 31780 21758
rect 31836 21588 31892 21598
rect 31948 21588 32004 22990
rect 32172 22258 32228 22270
rect 32172 22206 32174 22258
rect 32226 22206 32228 22258
rect 32172 21812 32228 22206
rect 32284 22148 32340 23996
rect 32396 23826 32452 23838
rect 32396 23774 32398 23826
rect 32450 23774 32452 23826
rect 32396 23716 32452 23774
rect 32396 23650 32452 23660
rect 32508 23042 32564 24220
rect 32620 24052 32676 24062
rect 32620 23958 32676 23996
rect 33180 23940 33236 23950
rect 33180 23846 33236 23884
rect 32620 23714 32676 23726
rect 32620 23662 32622 23714
rect 32674 23662 32676 23714
rect 32620 23380 32676 23662
rect 33292 23604 33348 29036
rect 33628 29026 33684 29036
rect 33628 28532 33684 28542
rect 33628 28196 33684 28476
rect 33404 28140 33684 28196
rect 33404 26290 33460 28140
rect 33516 27970 33572 27982
rect 33516 27918 33518 27970
rect 33570 27918 33572 27970
rect 33516 27412 33572 27918
rect 33628 27858 33684 28140
rect 33628 27806 33630 27858
rect 33682 27806 33684 27858
rect 33628 27794 33684 27806
rect 33516 27346 33572 27356
rect 33740 27188 33796 31500
rect 33852 31444 33908 31726
rect 34076 31780 34132 31790
rect 34076 31686 34132 31724
rect 33852 31378 33908 31388
rect 34524 31554 34580 31566
rect 34524 31502 34526 31554
rect 34578 31502 34580 31554
rect 34524 31444 34580 31502
rect 34524 31378 34580 31388
rect 35084 31106 35140 33068
rect 35420 32786 35476 33180
rect 35868 33170 35924 33180
rect 36316 33906 36484 33908
rect 36316 33854 36430 33906
rect 36482 33854 36484 33906
rect 36316 33852 36484 33854
rect 36316 33348 36372 33852
rect 36428 33842 36484 33852
rect 36764 33908 36820 33918
rect 36764 33906 36932 33908
rect 36764 33854 36766 33906
rect 36818 33854 36932 33906
rect 36764 33852 36932 33854
rect 36764 33842 36820 33852
rect 36876 33348 36932 33852
rect 36988 33572 37044 37548
rect 37324 37156 37380 37166
rect 37324 37062 37380 37100
rect 37436 36708 37492 36718
rect 37436 36594 37492 36652
rect 37436 36542 37438 36594
rect 37490 36542 37492 36594
rect 37436 36530 37492 36542
rect 37436 35586 37492 35598
rect 37436 35534 37438 35586
rect 37490 35534 37492 35586
rect 37100 34804 37156 34814
rect 37436 34804 37492 35534
rect 39228 35588 39284 35598
rect 39228 35494 39284 35532
rect 38220 35140 38276 35150
rect 37660 34916 37716 34926
rect 38220 34916 38276 35084
rect 37660 34914 38052 34916
rect 37660 34862 37662 34914
rect 37714 34862 38052 34914
rect 37660 34860 38052 34862
rect 37660 34850 37716 34860
rect 37156 34748 37492 34804
rect 37100 34710 37156 34748
rect 37884 34692 37940 34702
rect 37884 34598 37940 34636
rect 37996 34354 38052 34860
rect 38220 34822 38276 34860
rect 38892 35140 38948 35150
rect 37996 34302 37998 34354
rect 38050 34302 38052 34354
rect 37996 34290 38052 34302
rect 38556 34244 38612 34254
rect 38668 34244 38724 34254
rect 38612 34242 38724 34244
rect 38612 34190 38670 34242
rect 38722 34190 38724 34242
rect 38612 34188 38724 34190
rect 38332 34132 38388 34142
rect 38332 34038 38388 34076
rect 36988 33516 37156 33572
rect 36988 33348 37044 33358
rect 36876 33346 37044 33348
rect 36876 33294 36990 33346
rect 37042 33294 37044 33346
rect 36876 33292 37044 33294
rect 35420 32734 35422 32786
rect 35474 32734 35476 32786
rect 35420 32722 35476 32734
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35980 31556 36036 31566
rect 35644 31554 36036 31556
rect 35644 31502 35982 31554
rect 36034 31502 36036 31554
rect 35644 31500 36036 31502
rect 35644 31218 35700 31500
rect 35644 31166 35646 31218
rect 35698 31166 35700 31218
rect 35644 31154 35700 31166
rect 35084 31054 35086 31106
rect 35138 31054 35140 31106
rect 35084 31042 35140 31054
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35084 30322 35140 30334
rect 35084 30270 35086 30322
rect 35138 30270 35140 30322
rect 34076 29540 34132 29550
rect 33964 29316 34020 29326
rect 33964 29222 34020 29260
rect 33964 28532 34020 28542
rect 33516 27132 33796 27188
rect 33852 27412 33908 27422
rect 33852 27188 33908 27356
rect 33516 26740 33572 27132
rect 33852 26908 33908 27132
rect 33964 27074 34020 28476
rect 33964 27022 33966 27074
rect 34018 27022 34020 27074
rect 33964 27010 34020 27022
rect 33516 26674 33572 26684
rect 33628 26852 33908 26908
rect 34076 26908 34132 29484
rect 34524 29540 34580 29550
rect 34524 29446 34580 29484
rect 34300 29426 34356 29438
rect 34300 29374 34302 29426
rect 34354 29374 34356 29426
rect 34300 29316 34356 29374
rect 34972 29428 35028 29438
rect 35084 29428 35140 30270
rect 35532 30212 35588 30222
rect 35532 30118 35588 30156
rect 35980 29652 36036 31500
rect 36316 30882 36372 33292
rect 36988 33282 37044 33292
rect 36316 30830 36318 30882
rect 36370 30830 36372 30882
rect 36316 30100 36372 30830
rect 36316 30034 36372 30044
rect 36428 32676 36484 32686
rect 35980 29586 36036 29596
rect 34972 29426 35140 29428
rect 34972 29374 34974 29426
rect 35026 29374 35140 29426
rect 34972 29372 35140 29374
rect 35980 29426 36036 29438
rect 35980 29374 35982 29426
rect 36034 29374 36036 29426
rect 34972 29316 35028 29372
rect 34300 29260 35028 29316
rect 34188 28980 34244 28990
rect 34188 28754 34244 28924
rect 34188 28702 34190 28754
rect 34242 28702 34244 28754
rect 34188 28690 34244 28702
rect 34860 28642 34916 28654
rect 34860 28590 34862 28642
rect 34914 28590 34916 28642
rect 34524 28532 34580 28542
rect 34524 28438 34580 28476
rect 34860 28084 34916 28590
rect 34860 28018 34916 28028
rect 34636 27860 34692 27870
rect 34972 27860 35028 29260
rect 35532 29316 35588 29326
rect 35980 29316 36036 29374
rect 35532 29314 36036 29316
rect 35532 29262 35534 29314
rect 35586 29262 36036 29314
rect 35532 29260 36036 29262
rect 35532 29250 35588 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35980 28756 36036 29260
rect 36428 29314 36484 32620
rect 37100 30548 37156 33516
rect 38556 33460 38612 34188
rect 38668 34178 38724 34188
rect 38892 34242 38948 35084
rect 38892 34190 38894 34242
rect 38946 34190 38948 34242
rect 38892 34178 38948 34190
rect 39004 34468 39060 34478
rect 38444 33458 38612 33460
rect 38444 33406 38558 33458
rect 38610 33406 38612 33458
rect 38444 33404 38612 33406
rect 38220 33346 38276 33358
rect 38220 33294 38222 33346
rect 38274 33294 38276 33346
rect 37324 33122 37380 33134
rect 37324 33070 37326 33122
rect 37378 33070 37380 33122
rect 37324 32564 37380 33070
rect 37772 33124 37828 33134
rect 38220 33124 38276 33294
rect 37772 33122 38276 33124
rect 37772 33070 37774 33122
rect 37826 33070 38276 33122
rect 37772 33068 38276 33070
rect 37772 33058 37828 33068
rect 37772 32564 37828 32574
rect 37324 32562 37828 32564
rect 37324 32510 37774 32562
rect 37826 32510 37828 32562
rect 37324 32508 37828 32510
rect 37772 32498 37828 32508
rect 37212 31780 37268 31790
rect 37212 31778 37828 31780
rect 37212 31726 37214 31778
rect 37266 31726 37828 31778
rect 37212 31724 37828 31726
rect 37212 31714 37268 31724
rect 37436 31554 37492 31566
rect 37436 31502 37438 31554
rect 37490 31502 37492 31554
rect 37436 30996 37492 31502
rect 37436 30930 37492 30940
rect 37100 30492 37492 30548
rect 36428 29262 36430 29314
rect 36482 29262 36484 29314
rect 36428 29092 36484 29262
rect 36428 29026 36484 29036
rect 36764 29652 36820 29662
rect 36204 28868 36260 28878
rect 36092 28756 36148 28766
rect 35980 28700 36092 28756
rect 36092 28662 36148 28700
rect 34636 27858 35028 27860
rect 34636 27806 34638 27858
rect 34690 27806 35028 27858
rect 34636 27804 35028 27806
rect 35196 28532 35252 28542
rect 35196 27858 35252 28476
rect 35196 27806 35198 27858
rect 35250 27806 35252 27858
rect 34188 27746 34244 27758
rect 34188 27694 34190 27746
rect 34242 27694 34244 27746
rect 34188 27412 34244 27694
rect 34188 27346 34244 27356
rect 34636 27076 34692 27804
rect 35196 27794 35252 27806
rect 35420 28418 35476 28430
rect 35420 28366 35422 28418
rect 35474 28366 35476 28418
rect 35420 27860 35476 28366
rect 35980 28420 36036 28430
rect 36204 28420 36260 28812
rect 35980 28418 36260 28420
rect 35980 28366 35982 28418
rect 36034 28366 36260 28418
rect 35980 28364 36260 28366
rect 35980 28354 36036 28364
rect 35644 27860 35700 27870
rect 35420 27858 35700 27860
rect 35420 27806 35646 27858
rect 35698 27806 35700 27858
rect 35420 27804 35700 27806
rect 35644 27748 35700 27804
rect 36092 27748 36148 27758
rect 35644 27746 36148 27748
rect 35644 27694 36094 27746
rect 36146 27694 36148 27746
rect 35644 27692 36148 27694
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35644 27300 35700 27692
rect 36092 27682 36148 27692
rect 35084 27244 35700 27300
rect 34860 27076 34916 27086
rect 34636 27074 34916 27076
rect 34636 27022 34862 27074
rect 34914 27022 34916 27074
rect 34636 27020 34916 27022
rect 34860 27010 34916 27020
rect 35084 27074 35140 27244
rect 35084 27022 35086 27074
rect 35138 27022 35140 27074
rect 35084 27010 35140 27022
rect 35196 26962 35252 26974
rect 35196 26910 35198 26962
rect 35250 26910 35252 26962
rect 34076 26852 34244 26908
rect 33404 26238 33406 26290
rect 33458 26238 33460 26290
rect 33404 26226 33460 26238
rect 33516 26404 33572 26414
rect 33516 25284 33572 26348
rect 33628 26404 33684 26852
rect 33964 26404 34020 26414
rect 33628 26402 34020 26404
rect 33628 26350 33630 26402
rect 33682 26350 33966 26402
rect 34018 26350 34020 26402
rect 33628 26348 34020 26350
rect 33628 26338 33684 26348
rect 33964 26338 34020 26348
rect 33516 25228 33684 25284
rect 32620 23314 32676 23324
rect 33068 23548 33348 23604
rect 33628 23548 33684 25228
rect 34188 24500 34244 26852
rect 35196 26516 35252 26910
rect 35644 26850 35700 26862
rect 35644 26798 35646 26850
rect 35698 26798 35700 26850
rect 35308 26516 35364 26526
rect 35196 26514 35364 26516
rect 35196 26462 35310 26514
rect 35362 26462 35364 26514
rect 35196 26460 35364 26462
rect 35308 26404 35364 26460
rect 35308 26338 35364 26348
rect 34188 24434 34244 24444
rect 34412 26180 34468 26190
rect 33852 24052 33908 24062
rect 33852 23958 33908 23996
rect 32508 22990 32510 23042
rect 32562 22990 32564 23042
rect 32508 22932 32564 22990
rect 32508 22484 32564 22876
rect 32508 22428 32900 22484
rect 32732 22260 32788 22270
rect 32284 22092 32452 22148
rect 32172 21746 32228 21756
rect 32284 21700 32340 21710
rect 32284 21606 32340 21644
rect 31836 21586 32004 21588
rect 31836 21534 31838 21586
rect 31890 21534 32004 21586
rect 31836 21532 32004 21534
rect 32172 21586 32228 21598
rect 32172 21534 32174 21586
rect 32226 21534 32228 21586
rect 31724 21364 31780 21374
rect 31724 21270 31780 21308
rect 31836 20692 31892 21532
rect 32172 21364 32228 21534
rect 32172 21298 32228 21308
rect 32284 21362 32340 21374
rect 32284 21310 32286 21362
rect 32338 21310 32340 21362
rect 32284 21028 32340 21310
rect 32284 20962 32340 20972
rect 31948 20916 32004 20926
rect 31948 20822 32004 20860
rect 32396 20804 32452 22092
rect 32732 22146 32788 22204
rect 32732 22094 32734 22146
rect 32786 22094 32788 22146
rect 31836 20626 31892 20636
rect 32284 20692 32340 20702
rect 31724 20356 31780 20366
rect 31780 20300 31892 20356
rect 31724 20290 31780 20300
rect 31836 18452 31892 20300
rect 32172 20132 32228 20142
rect 32172 20038 32228 20076
rect 31948 19124 32004 19134
rect 31948 19030 32004 19068
rect 31948 18452 32004 18462
rect 31836 18396 31948 18452
rect 31948 18358 32004 18396
rect 31500 16996 31556 17006
rect 31388 16994 31556 16996
rect 31388 16942 31502 16994
rect 31554 16942 31556 16994
rect 31388 16940 31556 16942
rect 31388 16548 31444 16940
rect 31500 16930 31556 16940
rect 31612 16884 31668 17836
rect 32172 17778 32228 17790
rect 32172 17726 32174 17778
rect 32226 17726 32228 17778
rect 31724 17444 31780 17454
rect 31724 17350 31780 17388
rect 32172 17108 32228 17726
rect 32172 17042 32228 17052
rect 31724 16884 31780 16894
rect 31612 16882 32116 16884
rect 31612 16830 31726 16882
rect 31778 16830 32116 16882
rect 31612 16828 32116 16830
rect 31724 16818 31780 16828
rect 31276 16492 31444 16548
rect 31948 16658 32004 16670
rect 31948 16606 31950 16658
rect 32002 16606 32004 16658
rect 31276 16210 31332 16492
rect 31276 16158 31278 16210
rect 31330 16158 31332 16210
rect 31276 16146 31332 16158
rect 31164 15922 31220 15932
rect 31836 15988 31892 15998
rect 31948 15988 32004 16606
rect 31836 15986 32004 15988
rect 31836 15934 31838 15986
rect 31890 15934 32004 15986
rect 31836 15932 32004 15934
rect 31836 15764 31892 15932
rect 31500 15708 31892 15764
rect 30492 14914 30548 14924
rect 30940 15092 31108 15148
rect 31276 15652 31332 15662
rect 30380 14700 30548 14756
rect 30380 14530 30436 14542
rect 30380 14478 30382 14530
rect 30434 14478 30436 14530
rect 30380 14084 30436 14478
rect 30492 14084 30548 14700
rect 30940 14644 30996 15092
rect 30940 14578 30996 14588
rect 31052 14420 31108 14430
rect 31052 14326 31108 14364
rect 30940 14084 30996 14094
rect 30492 14028 30772 14084
rect 30380 14018 30436 14028
rect 30268 13022 30270 13074
rect 30322 13022 30324 13074
rect 30268 13010 30324 13022
rect 30492 13748 30548 13758
rect 30380 12740 30436 12750
rect 29932 12126 29934 12178
rect 29986 12126 29988 12178
rect 29820 12068 29876 12078
rect 29820 11954 29876 12012
rect 29820 11902 29822 11954
rect 29874 11902 29876 11954
rect 29820 11890 29876 11902
rect 29932 11732 29988 12126
rect 29932 11666 29988 11676
rect 30268 12178 30324 12190
rect 30268 12126 30270 12178
rect 30322 12126 30324 12178
rect 29708 9886 29710 9938
rect 29762 9886 29764 9938
rect 29708 9874 29764 9886
rect 29932 11506 29988 11518
rect 29932 11454 29934 11506
rect 29986 11454 29988 11506
rect 29372 9314 29428 9324
rect 29484 9604 29540 9614
rect 29148 9044 29204 9054
rect 29148 8950 29204 8988
rect 29260 8820 29316 8830
rect 29260 8258 29316 8764
rect 29484 8372 29540 9548
rect 29932 9268 29988 11454
rect 30268 11508 30324 12126
rect 30268 11442 30324 11452
rect 30380 11282 30436 12684
rect 30492 12402 30548 13692
rect 30492 12350 30494 12402
rect 30546 12350 30548 12402
rect 30492 12338 30548 12350
rect 30604 13412 30660 13422
rect 30492 12068 30548 12078
rect 30604 12068 30660 13356
rect 30716 13188 30772 14028
rect 30716 13122 30772 13132
rect 30828 13746 30884 13758
rect 30828 13694 30830 13746
rect 30882 13694 30884 13746
rect 30716 12964 30772 12974
rect 30716 12870 30772 12908
rect 30492 12066 30660 12068
rect 30492 12014 30494 12066
rect 30546 12014 30660 12066
rect 30492 12012 30660 12014
rect 30716 12178 30772 12190
rect 30716 12126 30718 12178
rect 30770 12126 30772 12178
rect 30492 12002 30548 12012
rect 30604 11396 30660 11406
rect 30604 11302 30660 11340
rect 30380 11230 30382 11282
rect 30434 11230 30436 11282
rect 30380 11218 30436 11230
rect 30716 10610 30772 12126
rect 30828 11396 30884 13694
rect 30828 11330 30884 11340
rect 30940 13748 30996 14028
rect 31052 13748 31108 13758
rect 30940 13746 31108 13748
rect 30940 13694 31054 13746
rect 31106 13694 31108 13746
rect 30940 13692 31108 13694
rect 30716 10558 30718 10610
rect 30770 10558 30772 10610
rect 30380 9716 30436 9726
rect 30268 9714 30436 9716
rect 30268 9662 30382 9714
rect 30434 9662 30436 9714
rect 30268 9660 30436 9662
rect 30044 9268 30100 9278
rect 29932 9212 30044 9268
rect 30044 9202 30100 9212
rect 29260 8206 29262 8258
rect 29314 8206 29316 8258
rect 29260 8194 29316 8206
rect 29372 8370 29540 8372
rect 29372 8318 29486 8370
rect 29538 8318 29540 8370
rect 29372 8316 29540 8318
rect 29260 7588 29316 7598
rect 29372 7588 29428 8316
rect 29484 8306 29540 8316
rect 29708 8372 29764 8382
rect 30268 8372 30324 9660
rect 30380 9650 30436 9660
rect 30716 9604 30772 10558
rect 30940 10612 30996 13692
rect 31052 13682 31108 13692
rect 31164 13636 31220 13646
rect 31164 13074 31220 13580
rect 31164 13022 31166 13074
rect 31218 13022 31220 13074
rect 31164 13010 31220 13022
rect 31052 12292 31108 12302
rect 31052 12178 31108 12236
rect 31052 12126 31054 12178
rect 31106 12126 31108 12178
rect 31052 12114 31108 12126
rect 31276 11060 31332 15596
rect 31500 15314 31556 15708
rect 31500 15262 31502 15314
rect 31554 15262 31556 15314
rect 31388 14532 31444 14542
rect 31388 14438 31444 14476
rect 31500 14420 31556 15262
rect 31948 15316 32004 15326
rect 31500 14326 31556 14364
rect 31724 15090 31780 15102
rect 31724 15038 31726 15090
rect 31778 15038 31780 15090
rect 31612 13636 31668 13646
rect 31612 13076 31668 13580
rect 31724 13188 31780 15038
rect 31948 14532 32004 15260
rect 31836 13860 31892 13870
rect 31948 13860 32004 14476
rect 31836 13858 32004 13860
rect 31836 13806 31838 13858
rect 31890 13806 32004 13858
rect 31836 13804 32004 13806
rect 31836 13794 31892 13804
rect 31724 13132 31892 13188
rect 31612 13020 31780 13076
rect 31724 12850 31780 13020
rect 31724 12798 31726 12850
rect 31778 12798 31780 12850
rect 31500 12292 31556 12302
rect 31500 12198 31556 12236
rect 31612 12068 31668 12078
rect 31612 11394 31668 12012
rect 31724 11732 31780 12798
rect 31724 11666 31780 11676
rect 31612 11342 31614 11394
rect 31666 11342 31668 11394
rect 31612 11330 31668 11342
rect 31836 11282 31892 13132
rect 31948 12962 32004 12974
rect 31948 12910 31950 12962
rect 32002 12910 32004 12962
rect 31948 12068 32004 12910
rect 31948 12002 32004 12012
rect 31836 11230 31838 11282
rect 31890 11230 31892 11282
rect 31836 11218 31892 11230
rect 31948 11732 32004 11742
rect 31276 11004 31780 11060
rect 31052 10612 31108 10622
rect 30940 10556 31052 10612
rect 31052 10518 31108 10556
rect 30716 9538 30772 9548
rect 30828 10276 30884 10286
rect 29260 7586 29428 7588
rect 29260 7534 29262 7586
rect 29314 7534 29428 7586
rect 29260 7532 29428 7534
rect 29708 7588 29764 8316
rect 29820 8316 30324 8372
rect 30380 9268 30436 9278
rect 29820 8258 29876 8316
rect 29820 8206 29822 8258
rect 29874 8206 29876 8258
rect 29820 7698 29876 8206
rect 30380 8146 30436 9212
rect 30380 8094 30382 8146
rect 30434 8094 30436 8146
rect 30380 8082 30436 8094
rect 30716 9044 30772 9054
rect 29932 8036 29988 8046
rect 29932 7942 29988 7980
rect 29820 7646 29822 7698
rect 29874 7646 29876 7698
rect 29820 7634 29876 7646
rect 29260 7522 29316 7532
rect 29708 7494 29764 7532
rect 29036 7422 29038 7474
rect 29090 7422 29092 7474
rect 29036 7410 29092 7422
rect 30716 7474 30772 8988
rect 30828 7698 30884 10220
rect 31052 9940 31108 9950
rect 31052 9826 31108 9884
rect 31052 9774 31054 9826
rect 31106 9774 31108 9826
rect 31052 9762 31108 9774
rect 31388 9828 31444 9838
rect 31388 9734 31444 9772
rect 31724 9716 31780 11004
rect 31836 10722 31892 10734
rect 31836 10670 31838 10722
rect 31890 10670 31892 10722
rect 31836 9940 31892 10670
rect 31948 10498 32004 11676
rect 31948 10446 31950 10498
rect 32002 10446 32004 10498
rect 31948 10434 32004 10446
rect 31836 9874 31892 9884
rect 31948 9716 32004 9726
rect 31724 9714 32004 9716
rect 31724 9662 31950 9714
rect 32002 9662 32004 9714
rect 31724 9660 32004 9662
rect 31500 9602 31556 9614
rect 31500 9550 31502 9602
rect 31554 9550 31556 9602
rect 31052 8930 31108 8942
rect 31052 8878 31054 8930
rect 31106 8878 31108 8930
rect 31052 8596 31108 8878
rect 31052 8530 31108 8540
rect 30828 7646 30830 7698
rect 30882 7646 30884 7698
rect 30828 7634 30884 7646
rect 30940 7700 30996 7710
rect 30716 7422 30718 7474
rect 30770 7422 30772 7474
rect 30716 7410 30772 7422
rect 30940 7476 30996 7644
rect 30940 7474 31332 7476
rect 30940 7422 30942 7474
rect 30994 7422 31332 7474
rect 30940 7420 31332 7422
rect 30940 7410 30996 7420
rect 29820 6802 29876 6814
rect 29820 6750 29822 6802
rect 29874 6750 29876 6802
rect 28364 6598 28420 6636
rect 29148 6692 29204 6702
rect 29148 6598 29204 6636
rect 29260 6690 29316 6702
rect 29260 6638 29262 6690
rect 29314 6638 29316 6690
rect 29260 6580 29316 6638
rect 29596 6692 29652 6702
rect 29596 6690 29764 6692
rect 29596 6638 29598 6690
rect 29650 6638 29764 6690
rect 29596 6636 29764 6638
rect 29596 6626 29652 6636
rect 29260 6514 29316 6524
rect 28028 6468 28084 6478
rect 28028 6374 28084 6412
rect 28252 6020 28308 6030
rect 27916 5964 28252 6020
rect 28252 5926 28308 5964
rect 26908 5854 26910 5906
rect 26962 5854 26964 5906
rect 26908 5842 26964 5854
rect 28364 5906 28420 5918
rect 28364 5854 28366 5906
rect 28418 5854 28420 5906
rect 26684 5796 26740 5806
rect 26572 5740 26684 5796
rect 26012 5702 26068 5740
rect 26684 5702 26740 5740
rect 25228 5684 25284 5694
rect 24892 5236 24948 5246
rect 23212 4946 23268 4956
rect 24444 5234 24948 5236
rect 24444 5182 24894 5234
rect 24946 5182 24948 5234
rect 24444 5180 24948 5182
rect 22540 4398 22542 4450
rect 22594 4398 22596 4450
rect 22540 4386 22596 4398
rect 22764 4898 22820 4910
rect 22764 4846 22766 4898
rect 22818 4846 22820 4898
rect 22092 3780 22148 3790
rect 21980 3724 22092 3780
rect 21084 3686 21140 3724
rect 22092 3714 22148 3724
rect 21420 3556 21476 3566
rect 21420 3462 21476 3500
rect 20972 3390 20974 3442
rect 21026 3390 21028 3442
rect 20972 3378 21028 3390
rect 22764 3388 22820 4846
rect 22652 3332 22820 3388
rect 23212 3442 23268 3454
rect 23212 3390 23214 3442
rect 23266 3390 23268 3442
rect 23212 3388 23268 3390
rect 23212 3332 23380 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 19628 2940 20020 2996
rect 19964 800 20020 2940
rect 22652 980 22708 3332
rect 22204 924 22708 980
rect 22204 800 22260 924
rect 23324 800 23380 3332
rect 24444 800 24500 5180
rect 24892 5170 24948 5180
rect 24780 5012 24836 5022
rect 24668 4228 24724 4238
rect 24668 4134 24724 4172
rect 24556 3780 24612 3790
rect 24556 3686 24612 3724
rect 24780 3442 24836 4956
rect 25228 4788 25284 5628
rect 27244 5292 28308 5348
rect 27244 5122 27300 5292
rect 27244 5070 27246 5122
rect 27298 5070 27300 5122
rect 27244 5058 27300 5070
rect 27580 5124 27636 5134
rect 27580 5030 27636 5068
rect 28252 5010 28308 5292
rect 28252 4958 28254 5010
rect 28306 4958 28308 5010
rect 28252 4946 28308 4958
rect 28364 5236 28420 5854
rect 29596 5794 29652 5806
rect 29596 5742 29598 5794
rect 29650 5742 29652 5794
rect 28812 5684 28868 5694
rect 28812 5590 28868 5628
rect 29148 5682 29204 5694
rect 29148 5630 29150 5682
rect 29202 5630 29204 5682
rect 27916 4900 27972 4910
rect 27916 4898 28084 4900
rect 27916 4846 27918 4898
rect 27970 4846 28084 4898
rect 27916 4844 28084 4846
rect 27916 4834 27972 4844
rect 25228 4722 25284 4732
rect 24892 4452 24948 4462
rect 24892 3778 24948 4396
rect 25900 4450 25956 4462
rect 25900 4398 25902 4450
rect 25954 4398 25956 4450
rect 25900 4340 25956 4398
rect 26236 4452 26292 4462
rect 26236 4358 26292 4396
rect 25900 4274 25956 4284
rect 26908 4340 26964 4350
rect 26908 4246 26964 4284
rect 25676 4228 25732 4238
rect 25676 4134 25732 4172
rect 25340 4116 25396 4126
rect 25340 4022 25396 4060
rect 26684 4116 26740 4126
rect 24892 3726 24894 3778
rect 24946 3726 24948 3778
rect 24892 3714 24948 3726
rect 24780 3390 24782 3442
rect 24834 3390 24836 3442
rect 24780 3378 24836 3390
rect 25228 3554 25284 3566
rect 25228 3502 25230 3554
rect 25282 3502 25284 3554
rect 25228 3444 25284 3502
rect 25228 3378 25284 3388
rect 26236 3330 26292 3342
rect 26236 3278 26238 3330
rect 26290 3278 26292 3330
rect 25564 924 25956 980
rect 25564 800 25620 924
rect 2492 700 2884 756
rect 3136 0 3248 800
rect 4256 0 4368 800
rect 5376 0 5488 800
rect 6496 0 6608 800
rect 7616 0 7728 800
rect 8736 0 8848 800
rect 9856 0 9968 800
rect 10976 0 11088 800
rect 12096 0 12208 800
rect 13216 0 13328 800
rect 14336 0 14448 800
rect 15456 0 15568 800
rect 16576 0 16688 800
rect 17696 0 17808 800
rect 18816 0 18928 800
rect 19936 0 20048 800
rect 21056 0 21168 800
rect 22176 0 22288 800
rect 23296 0 23408 800
rect 24416 0 24528 800
rect 25536 0 25648 800
rect 25900 756 25956 924
rect 26236 756 26292 3278
rect 26684 800 26740 4060
rect 27916 4116 27972 4126
rect 27916 4022 27972 4060
rect 27804 3668 27860 3678
rect 27804 800 27860 3612
rect 28028 3556 28084 4844
rect 28364 4228 28420 5180
rect 28588 5124 28644 5134
rect 28588 5030 28644 5068
rect 28364 4162 28420 4172
rect 28924 4116 28980 4126
rect 28364 3556 28420 3566
rect 28028 3554 28420 3556
rect 28028 3502 28366 3554
rect 28418 3502 28420 3554
rect 28028 3500 28420 3502
rect 28364 3490 28420 3500
rect 28924 800 28980 4060
rect 29148 3556 29204 5630
rect 29596 5346 29652 5742
rect 29596 5294 29598 5346
rect 29650 5294 29652 5346
rect 29596 5282 29652 5294
rect 29260 5124 29316 5134
rect 29260 5030 29316 5068
rect 29596 5012 29652 5022
rect 29708 5012 29764 6636
rect 29820 6468 29876 6750
rect 31276 6802 31332 7420
rect 31500 7474 31556 9550
rect 31836 8258 31892 9660
rect 31948 9650 32004 9660
rect 32060 9716 32116 16828
rect 32172 16660 32228 16670
rect 32172 16566 32228 16604
rect 32284 15652 32340 20636
rect 32396 20690 32452 20748
rect 32396 20638 32398 20690
rect 32450 20638 32452 20690
rect 32396 20626 32452 20638
rect 32508 21700 32564 21710
rect 32508 20468 32564 21644
rect 32620 20692 32676 20702
rect 32620 20598 32676 20636
rect 32508 20412 32676 20468
rect 32396 20132 32452 20142
rect 32396 20038 32452 20076
rect 32508 20018 32564 20030
rect 32508 19966 32510 20018
rect 32562 19966 32564 20018
rect 32508 18676 32564 19966
rect 32508 18582 32564 18620
rect 32620 18452 32676 20412
rect 32732 20132 32788 22094
rect 32844 21028 32900 22428
rect 33068 22258 33124 23548
rect 33628 23492 33908 23548
rect 33068 22206 33070 22258
rect 33122 22206 33124 22258
rect 33068 22036 33124 22206
rect 33068 21970 33124 21980
rect 33292 23380 33348 23390
rect 33180 21700 33236 21710
rect 32844 20962 32900 20972
rect 33068 21698 33236 21700
rect 33068 21646 33182 21698
rect 33234 21646 33236 21698
rect 33068 21644 33236 21646
rect 32844 20690 32900 20702
rect 32844 20638 32846 20690
rect 32898 20638 32900 20690
rect 32844 20580 32900 20638
rect 32844 20514 32900 20524
rect 32956 20578 33012 20590
rect 32956 20526 32958 20578
rect 33010 20526 33012 20578
rect 32844 20132 32900 20142
rect 32732 20076 32844 20132
rect 32844 20066 32900 20076
rect 32284 15586 32340 15596
rect 32508 18396 32676 18452
rect 32844 19684 32900 19694
rect 32284 15316 32340 15326
rect 32284 15222 32340 15260
rect 32508 15148 32564 18396
rect 32732 17892 32788 17902
rect 32732 17778 32788 17836
rect 32732 17726 32734 17778
rect 32786 17726 32788 17778
rect 32732 17714 32788 17726
rect 32620 16658 32676 16670
rect 32620 16606 32622 16658
rect 32674 16606 32676 16658
rect 32620 15652 32676 16606
rect 32620 15586 32676 15596
rect 32396 15092 32564 15148
rect 32844 15148 32900 19628
rect 32956 15876 33012 20526
rect 33068 19908 33124 21644
rect 33180 21634 33236 21644
rect 33292 21586 33348 23324
rect 33740 22260 33796 22270
rect 33740 22166 33796 22204
rect 33292 21534 33294 21586
rect 33346 21534 33348 21586
rect 33292 21522 33348 21534
rect 33628 21474 33684 21486
rect 33628 21422 33630 21474
rect 33682 21422 33684 21474
rect 33292 21028 33348 21038
rect 33068 19842 33124 19852
rect 33180 20578 33236 20590
rect 33180 20526 33182 20578
rect 33234 20526 33236 20578
rect 33068 19124 33124 19134
rect 33068 18676 33124 19068
rect 33068 17780 33124 18620
rect 33180 18450 33236 20526
rect 33180 18398 33182 18450
rect 33234 18398 33236 18450
rect 33180 18386 33236 18398
rect 33292 18452 33348 20972
rect 33516 20916 33572 20926
rect 33404 20804 33460 20814
rect 33404 20710 33460 20748
rect 33516 20690 33572 20860
rect 33516 20638 33518 20690
rect 33570 20638 33572 20690
rect 33516 20626 33572 20638
rect 33516 20132 33572 20142
rect 33404 20018 33460 20030
rect 33404 19966 33406 20018
rect 33458 19966 33460 20018
rect 33404 19346 33460 19966
rect 33404 19294 33406 19346
rect 33458 19294 33460 19346
rect 33404 19282 33460 19294
rect 33404 18452 33460 18462
rect 33292 18450 33460 18452
rect 33292 18398 33406 18450
rect 33458 18398 33460 18450
rect 33292 18396 33460 18398
rect 33404 18386 33460 18396
rect 33068 17724 33236 17780
rect 33180 17666 33236 17724
rect 33180 17614 33182 17666
rect 33234 17614 33236 17666
rect 33180 17602 33236 17614
rect 33516 17666 33572 20076
rect 33628 19906 33684 21422
rect 33740 20804 33796 20814
rect 33740 20710 33796 20748
rect 33852 20244 33908 23492
rect 34076 23380 34132 23390
rect 34076 23286 34132 23324
rect 34188 23042 34244 23054
rect 34188 22990 34190 23042
rect 34242 22990 34244 23042
rect 33964 22372 34020 22382
rect 33964 22278 34020 22316
rect 34188 22260 34244 22990
rect 34412 22820 34468 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34524 24724 34580 24734
rect 34524 23266 34580 24668
rect 34524 23214 34526 23266
rect 34578 23214 34580 23266
rect 34524 23202 34580 23214
rect 34748 24500 34804 24510
rect 34748 23154 34804 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34748 23102 34750 23154
rect 34802 23102 34804 23154
rect 34748 23090 34804 23102
rect 34412 22754 34468 22764
rect 34972 22930 35028 22942
rect 34972 22878 34974 22930
rect 35026 22878 35028 22930
rect 34860 22370 34916 22382
rect 34860 22318 34862 22370
rect 34914 22318 34916 22370
rect 34412 22260 34468 22270
rect 34188 22258 34468 22260
rect 34188 22206 34414 22258
rect 34466 22206 34468 22258
rect 34188 22204 34468 22206
rect 34076 21812 34132 21822
rect 34076 21586 34132 21756
rect 34412 21812 34468 22204
rect 34860 22260 34916 22318
rect 34860 22194 34916 22204
rect 34412 21746 34468 21756
rect 34076 21534 34078 21586
rect 34130 21534 34132 21586
rect 34076 21522 34132 21534
rect 34524 21588 34580 21598
rect 34524 21494 34580 21532
rect 34188 21028 34244 21038
rect 34188 20934 34244 20972
rect 34636 20804 34692 20814
rect 34860 20804 34916 20814
rect 34692 20802 34916 20804
rect 34692 20750 34862 20802
rect 34914 20750 34916 20802
rect 34692 20748 34916 20750
rect 34636 20738 34692 20748
rect 34860 20738 34916 20748
rect 34972 20804 35028 22878
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35644 22596 35700 26798
rect 35756 26178 35812 26190
rect 35756 26126 35758 26178
rect 35810 26126 35812 26178
rect 35756 25508 35812 26126
rect 35756 24834 35812 25452
rect 35756 24782 35758 24834
rect 35810 24782 35812 24834
rect 35756 23154 35812 24782
rect 35756 23102 35758 23154
rect 35810 23102 35812 23154
rect 35756 23090 35812 23102
rect 35980 24722 36036 24734
rect 35980 24670 35982 24722
rect 36034 24670 36036 24722
rect 35980 24050 36036 24670
rect 35980 23998 35982 24050
rect 36034 23998 36036 24050
rect 35980 23268 36036 23998
rect 36092 23268 36148 23278
rect 35980 23266 36148 23268
rect 35980 23214 36094 23266
rect 36146 23214 36148 23266
rect 35980 23212 36148 23214
rect 35196 22540 35700 22596
rect 35196 22482 35252 22540
rect 35196 22430 35198 22482
rect 35250 22430 35252 22482
rect 35196 22418 35252 22430
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34524 20690 34580 20702
rect 34524 20638 34526 20690
rect 34578 20638 34580 20690
rect 33852 20178 33908 20188
rect 34300 20578 34356 20590
rect 34300 20526 34302 20578
rect 34354 20526 34356 20578
rect 34300 20356 34356 20526
rect 34524 20580 34580 20638
rect 34972 20690 35028 20748
rect 34972 20638 34974 20690
rect 35026 20638 35028 20690
rect 34972 20626 35028 20638
rect 34524 20514 34580 20524
rect 35196 20578 35252 20590
rect 35196 20526 35198 20578
rect 35250 20526 35252 20578
rect 35196 20356 35252 20526
rect 34300 20300 35252 20356
rect 33740 20020 33796 20029
rect 33852 20020 33908 20030
rect 33740 20017 33852 20020
rect 33740 19965 33742 20017
rect 33794 19965 33852 20017
rect 33740 19964 33852 19965
rect 33740 19953 33796 19964
rect 33852 19954 33908 19964
rect 34076 20020 34132 20030
rect 33628 19854 33630 19906
rect 33682 19854 33684 19906
rect 33628 19842 33684 19854
rect 33516 17614 33518 17666
rect 33570 17614 33572 17666
rect 33516 17602 33572 17614
rect 33964 19122 34020 19134
rect 33964 19070 33966 19122
rect 34018 19070 34020 19122
rect 33964 18452 34020 19070
rect 34076 18674 34132 19964
rect 34076 18622 34078 18674
rect 34130 18622 34132 18674
rect 34076 18610 34132 18622
rect 34188 19908 34244 19918
rect 33068 17554 33124 17566
rect 33068 17502 33070 17554
rect 33122 17502 33124 17554
rect 33068 17332 33124 17502
rect 33068 16884 33124 17276
rect 33516 17332 33572 17342
rect 33516 16996 33572 17276
rect 33516 16930 33572 16940
rect 33740 16996 33796 17006
rect 33740 16902 33796 16940
rect 33180 16884 33236 16894
rect 33068 16882 33236 16884
rect 33068 16830 33182 16882
rect 33234 16830 33236 16882
rect 33068 16828 33236 16830
rect 33964 16884 34020 18396
rect 34188 18450 34244 19852
rect 34300 18562 34356 20300
rect 34860 20132 34916 20142
rect 34412 20020 34468 20030
rect 34412 19926 34468 19964
rect 34300 18510 34302 18562
rect 34354 18510 34356 18562
rect 34300 18498 34356 18510
rect 34524 19234 34580 19246
rect 34524 19182 34526 19234
rect 34578 19182 34580 19234
rect 34188 18398 34190 18450
rect 34242 18398 34244 18450
rect 34188 18386 34244 18398
rect 34524 17780 34580 19182
rect 34188 17444 34244 17454
rect 34076 17442 34244 17444
rect 34076 17390 34190 17442
rect 34242 17390 34244 17442
rect 34076 17388 34244 17390
rect 34076 17108 34132 17388
rect 34188 17378 34244 17388
rect 34524 17332 34580 17724
rect 34748 17780 34804 17790
rect 34748 17686 34804 17724
rect 34076 17042 34132 17052
rect 34300 17276 34580 17332
rect 34188 16994 34244 17006
rect 34188 16942 34190 16994
rect 34242 16942 34244 16994
rect 34188 16884 34244 16942
rect 34300 16996 34356 17276
rect 34300 16902 34356 16940
rect 34636 17220 34692 17230
rect 34860 17220 34916 20076
rect 35532 20130 35588 22540
rect 35868 22372 35924 22382
rect 35980 22372 36036 23212
rect 36092 23202 36148 23212
rect 36204 22708 36260 28364
rect 36764 26908 36820 29596
rect 37100 29426 37156 29438
rect 37100 29374 37102 29426
rect 37154 29374 37156 29426
rect 36988 29316 37044 29326
rect 36988 27298 37044 29260
rect 36988 27246 36990 27298
rect 37042 27246 37044 27298
rect 36988 27188 37044 27246
rect 36988 27122 37044 27132
rect 37100 28756 37156 29374
rect 36652 26852 36820 26908
rect 36540 24724 36596 24734
rect 36540 24630 36596 24668
rect 35868 22370 36036 22372
rect 35868 22318 35870 22370
rect 35922 22318 36036 22370
rect 35868 22316 36036 22318
rect 36092 22652 36260 22708
rect 36316 24498 36372 24510
rect 36316 24446 36318 24498
rect 36370 24446 36372 24498
rect 35868 22306 35924 22316
rect 36092 22148 36148 22652
rect 36204 22482 36260 22494
rect 36204 22430 36206 22482
rect 36258 22430 36260 22482
rect 36204 22372 36260 22430
rect 36316 22484 36372 24446
rect 36428 24052 36484 24090
rect 36428 23986 36484 23996
rect 36652 24052 36708 26852
rect 36988 26404 37044 26414
rect 36988 25618 37044 26348
rect 36988 25566 36990 25618
rect 37042 25566 37044 25618
rect 36988 25554 37044 25566
rect 36764 24836 36820 24846
rect 37100 24836 37156 28700
rect 37436 28868 37492 30492
rect 37772 30434 37828 31724
rect 37772 30382 37774 30434
rect 37826 30382 37828 30434
rect 37772 30370 37828 30382
rect 38108 30212 38164 30222
rect 38108 30118 38164 30156
rect 37436 28754 37492 28812
rect 38220 28868 38276 33068
rect 38444 30098 38500 33404
rect 38556 33394 38612 33404
rect 38556 32564 38612 32574
rect 38556 32470 38612 32508
rect 38668 30996 38724 31006
rect 38668 30902 38724 30940
rect 38444 30046 38446 30098
rect 38498 30046 38500 30098
rect 38444 30034 38500 30046
rect 38668 30100 38724 30110
rect 38668 30006 38724 30044
rect 39004 29876 39060 34412
rect 39340 34356 39396 41692
rect 39452 41188 39508 41198
rect 39788 41188 39844 42030
rect 40124 42084 40180 42140
rect 40684 42084 40740 42478
rect 40124 42028 40740 42084
rect 39452 41186 39844 41188
rect 39452 41134 39454 41186
rect 39506 41134 39844 41186
rect 39452 41132 39844 41134
rect 40012 41970 40068 41982
rect 40012 41918 40014 41970
rect 40066 41918 40068 41970
rect 39452 41122 39508 41132
rect 40012 40964 40068 41918
rect 40012 40898 40068 40908
rect 40124 41076 40180 41086
rect 40012 40516 40068 40526
rect 40012 40422 40068 40460
rect 40124 40402 40180 41020
rect 40124 40350 40126 40402
rect 40178 40350 40180 40402
rect 40124 40338 40180 40350
rect 39340 34290 39396 34300
rect 39452 40180 39508 40190
rect 40236 40180 40292 42028
rect 39452 40178 40292 40180
rect 39452 40126 39454 40178
rect 39506 40126 40292 40178
rect 39452 40124 40292 40126
rect 40684 40964 40740 40974
rect 40684 40516 40740 40908
rect 39452 33124 39508 40124
rect 40348 39394 40404 39406
rect 40348 39342 40350 39394
rect 40402 39342 40404 39394
rect 39564 38946 39620 38958
rect 39564 38894 39566 38946
rect 39618 38894 39620 38946
rect 39564 37268 39620 38894
rect 40012 38836 40068 38846
rect 40012 38724 40068 38780
rect 40348 38724 40404 39342
rect 40012 38722 40404 38724
rect 40012 38670 40014 38722
rect 40066 38670 40404 38722
rect 40012 38668 40404 38670
rect 40012 38658 40068 38668
rect 39788 38050 39844 38062
rect 39788 37998 39790 38050
rect 39842 37998 39844 38050
rect 39788 37828 39844 37998
rect 40348 38052 40404 38668
rect 40572 38052 40628 38062
rect 40348 38050 40628 38052
rect 40348 37998 40574 38050
rect 40626 37998 40628 38050
rect 40348 37996 40628 37998
rect 39676 37268 39732 37278
rect 39564 37266 39732 37268
rect 39564 37214 39678 37266
rect 39730 37214 39732 37266
rect 39564 37212 39732 37214
rect 39676 37202 39732 37212
rect 39788 37268 39844 37772
rect 39788 37202 39844 37212
rect 39900 37940 39956 37950
rect 39900 37156 39956 37884
rect 39900 37090 39956 37100
rect 40460 37268 40516 37996
rect 40572 37986 40628 37996
rect 39788 36708 39844 36718
rect 39788 35698 39844 36652
rect 40460 36260 40516 37212
rect 40572 36260 40628 36270
rect 40460 36258 40628 36260
rect 40460 36206 40574 36258
rect 40626 36206 40628 36258
rect 40460 36204 40628 36206
rect 39788 35646 39790 35698
rect 39842 35646 39844 35698
rect 39676 34356 39732 34366
rect 39788 34356 39844 35646
rect 40572 35588 40628 36204
rect 40572 35522 40628 35532
rect 40572 34916 40628 34926
rect 40572 34822 40628 34860
rect 39564 34354 39844 34356
rect 39564 34302 39678 34354
rect 39730 34302 39844 34354
rect 39564 34300 39844 34302
rect 39564 33346 39620 34300
rect 39676 34290 39732 34300
rect 39564 33294 39566 33346
rect 39618 33294 39620 33346
rect 39564 33282 39620 33294
rect 40012 33460 40068 33470
rect 39452 33068 39844 33124
rect 39340 32788 39396 32798
rect 39340 32786 39620 32788
rect 39340 32734 39342 32786
rect 39394 32734 39620 32786
rect 39340 32732 39620 32734
rect 39340 32722 39396 32732
rect 39452 32564 39508 32574
rect 39452 32004 39508 32508
rect 39452 30994 39508 31948
rect 39452 30942 39454 30994
rect 39506 30942 39508 30994
rect 39452 30930 39508 30942
rect 39564 32450 39620 32732
rect 39788 32562 39844 33068
rect 39788 32510 39790 32562
rect 39842 32510 39844 32562
rect 39788 32498 39844 32510
rect 39564 32398 39566 32450
rect 39618 32398 39620 32450
rect 39564 31668 39620 32398
rect 40012 31892 40068 33404
rect 40124 32564 40180 32574
rect 40124 32450 40180 32508
rect 40124 32398 40126 32450
rect 40178 32398 40180 32450
rect 40124 32386 40180 32398
rect 40684 32228 40740 40460
rect 40348 32172 40740 32228
rect 40124 31892 40180 31902
rect 40012 31890 40180 31892
rect 40012 31838 40126 31890
rect 40178 31838 40180 31890
rect 40012 31836 40180 31838
rect 40124 31826 40180 31836
rect 39228 30212 39284 30222
rect 39004 29810 39060 29820
rect 39116 30156 39228 30212
rect 38668 29426 38724 29438
rect 38668 29374 38670 29426
rect 38722 29374 38724 29426
rect 38332 29316 38388 29326
rect 38668 29316 38724 29374
rect 38332 29314 38724 29316
rect 38332 29262 38334 29314
rect 38386 29262 38724 29314
rect 38332 29260 38724 29262
rect 38332 29204 38388 29260
rect 38332 29138 38388 29148
rect 38220 28802 38276 28812
rect 38780 28868 38836 28878
rect 37436 28702 37438 28754
rect 37490 28702 37492 28754
rect 37436 28690 37492 28702
rect 38556 28644 38612 28654
rect 38668 28644 38724 28654
rect 38556 28642 38668 28644
rect 38556 28590 38558 28642
rect 38610 28590 38668 28642
rect 38556 28588 38668 28590
rect 37996 28418 38052 28430
rect 37996 28366 37998 28418
rect 38050 28366 38052 28418
rect 37996 27972 38052 28366
rect 38556 28196 38612 28588
rect 38668 28578 38724 28588
rect 38556 28130 38612 28140
rect 37996 27906 38052 27916
rect 38220 27748 38276 27758
rect 37324 27746 38276 27748
rect 37324 27694 38222 27746
rect 38274 27694 38276 27746
rect 37324 27692 38276 27694
rect 37324 27298 37380 27692
rect 38220 27682 38276 27692
rect 37324 27246 37326 27298
rect 37378 27246 37380 27298
rect 37324 27234 37380 27246
rect 37660 27524 37716 27534
rect 36764 24834 37156 24836
rect 36764 24782 36766 24834
rect 36818 24782 37156 24834
rect 36764 24780 37156 24782
rect 37212 26964 37268 27002
rect 36764 24770 36820 24780
rect 36652 23986 36708 23996
rect 36988 24164 37044 24174
rect 37044 24108 37156 24164
rect 36428 23548 36484 23558
rect 36988 23548 37044 24108
rect 37100 23938 37156 24108
rect 37100 23886 37102 23938
rect 37154 23886 37156 23938
rect 37100 23874 37156 23886
rect 36428 22596 36484 23492
rect 36540 23492 37044 23548
rect 36540 23266 36596 23492
rect 36540 23214 36542 23266
rect 36594 23214 36596 23266
rect 36540 23202 36596 23214
rect 36764 23266 36820 23278
rect 36764 23214 36766 23266
rect 36818 23214 36820 23266
rect 36764 22932 36820 23214
rect 36764 22866 36820 22876
rect 36876 22930 36932 22942
rect 36876 22878 36878 22930
rect 36930 22878 36932 22930
rect 36428 22540 36820 22596
rect 36316 22428 36596 22484
rect 36260 22316 36484 22372
rect 36204 22306 36260 22316
rect 35868 22092 36148 22148
rect 35756 21588 35812 21598
rect 35756 21494 35812 21532
rect 35532 20078 35534 20130
rect 35586 20078 35588 20130
rect 35532 20066 35588 20078
rect 35644 21364 35700 21374
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34972 19010 35028 19022
rect 34972 18958 34974 19010
rect 35026 18958 35028 19010
rect 34972 18900 35028 18958
rect 35308 19012 35364 19022
rect 35308 18918 35364 18956
rect 34972 18834 35028 18844
rect 35420 18900 35476 18910
rect 35476 18844 35588 18900
rect 35420 18834 35476 18844
rect 35532 18450 35588 18844
rect 35532 18398 35534 18450
rect 35586 18398 35588 18450
rect 35532 18386 35588 18398
rect 35084 18338 35140 18350
rect 35084 18286 35086 18338
rect 35138 18286 35140 18338
rect 35084 17892 35140 18286
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35084 17826 35140 17836
rect 35420 17892 35476 17902
rect 35420 17666 35476 17836
rect 35532 17780 35588 17790
rect 35644 17780 35700 21308
rect 35532 17778 35700 17780
rect 35532 17726 35534 17778
rect 35586 17726 35700 17778
rect 35532 17724 35700 17726
rect 35756 19012 35812 19022
rect 35532 17714 35588 17724
rect 35420 17614 35422 17666
rect 35474 17614 35476 17666
rect 35420 17602 35476 17614
rect 35644 17556 35700 17566
rect 35756 17556 35812 18956
rect 35868 18900 35924 22092
rect 36092 21924 36148 21934
rect 36092 21586 36148 21868
rect 36092 21534 36094 21586
rect 36146 21534 36148 21586
rect 36092 21522 36148 21534
rect 36316 21812 36372 21822
rect 36316 21586 36372 21756
rect 36316 21534 36318 21586
rect 36370 21534 36372 21586
rect 36316 21522 36372 21534
rect 36428 20130 36484 22316
rect 36428 20078 36430 20130
rect 36482 20078 36484 20130
rect 36428 20066 36484 20078
rect 36204 20018 36260 20030
rect 36204 19966 36206 20018
rect 36258 19966 36260 20018
rect 36204 19796 36260 19966
rect 36204 19730 36260 19740
rect 36428 19906 36484 19918
rect 36428 19854 36430 19906
rect 36482 19854 36484 19906
rect 35868 18834 35924 18844
rect 35980 19346 36036 19358
rect 35980 19294 35982 19346
rect 36034 19294 36036 19346
rect 35980 18564 36036 19294
rect 36428 19236 36484 19854
rect 36540 19684 36596 22428
rect 36540 19618 36596 19628
rect 36428 19142 36484 19180
rect 35980 18498 36036 18508
rect 36652 18562 36708 18574
rect 36652 18510 36654 18562
rect 36706 18510 36708 18562
rect 36428 18450 36484 18462
rect 36428 18398 36430 18450
rect 36482 18398 36484 18450
rect 35980 18338 36036 18350
rect 35980 18286 35982 18338
rect 36034 18286 36036 18338
rect 35980 18004 36036 18286
rect 36428 18340 36484 18398
rect 36652 18452 36708 18510
rect 36652 18386 36708 18396
rect 36428 18274 36484 18284
rect 36428 18004 36484 18014
rect 35980 17948 36428 18004
rect 35644 17554 35756 17556
rect 35644 17502 35646 17554
rect 35698 17502 35756 17554
rect 35644 17500 35756 17502
rect 35812 17500 35924 17556
rect 35644 17490 35700 17500
rect 35756 17462 35812 17500
rect 35196 17442 35252 17454
rect 35196 17390 35198 17442
rect 35250 17390 35252 17442
rect 34860 17164 35028 17220
rect 33964 16828 34244 16884
rect 33180 16818 33236 16828
rect 33516 16770 33572 16782
rect 33516 16718 33518 16770
rect 33570 16718 33572 16770
rect 33516 16660 33572 16718
rect 34636 16770 34692 17164
rect 34636 16718 34638 16770
rect 34690 16718 34692 16770
rect 34636 16706 34692 16718
rect 34748 16996 34804 17006
rect 33516 16594 33572 16604
rect 34188 16658 34244 16670
rect 34188 16606 34190 16658
rect 34242 16606 34244 16658
rect 33404 16098 33460 16110
rect 33404 16046 33406 16098
rect 33458 16046 33460 16098
rect 33180 15876 33236 15886
rect 32956 15820 33180 15876
rect 33180 15782 33236 15820
rect 33180 15652 33236 15662
rect 33180 15314 33236 15596
rect 33180 15262 33182 15314
rect 33234 15262 33236 15314
rect 33180 15250 33236 15262
rect 33404 15316 33460 16046
rect 33404 15222 33460 15260
rect 33740 16098 33796 16110
rect 33740 16046 33742 16098
rect 33794 16046 33796 16098
rect 33740 15314 33796 16046
rect 33740 15262 33742 15314
rect 33794 15262 33796 15314
rect 33740 15148 33796 15262
rect 32844 15092 33124 15148
rect 32284 14532 32340 14542
rect 32284 13074 32340 14476
rect 32396 14306 32452 15092
rect 32396 14254 32398 14306
rect 32450 14254 32452 14306
rect 32396 14242 32452 14254
rect 32284 13022 32286 13074
rect 32338 13022 32340 13074
rect 32284 13010 32340 13022
rect 32732 13748 32788 13758
rect 32732 13074 32788 13692
rect 32732 13022 32734 13074
rect 32786 13022 32788 13074
rect 32732 13010 32788 13022
rect 33068 13076 33124 15092
rect 33404 15092 33796 15148
rect 34076 15204 34132 15214
rect 33404 14532 33460 15092
rect 33964 14980 34020 14990
rect 33404 14438 33460 14476
rect 33740 14868 33796 14878
rect 33628 13746 33684 13758
rect 33628 13694 33630 13746
rect 33682 13694 33684 13746
rect 33180 13636 33236 13646
rect 33180 13542 33236 13580
rect 33628 13636 33684 13694
rect 33292 13524 33348 13534
rect 33180 13076 33236 13086
rect 33068 13020 33180 13076
rect 33180 12982 33236 13020
rect 32620 12740 32676 12750
rect 32620 12646 32676 12684
rect 33292 12404 33348 13468
rect 33292 12338 33348 12348
rect 33516 12964 33572 12974
rect 32284 12290 32340 12302
rect 32284 12238 32286 12290
rect 32338 12238 32340 12290
rect 32060 9650 32116 9660
rect 32172 11506 32228 11518
rect 32172 11454 32174 11506
rect 32226 11454 32228 11506
rect 32172 9380 32228 11454
rect 32284 9492 32340 12238
rect 32396 12292 32452 12302
rect 32396 11284 32452 12236
rect 33068 12292 33124 12302
rect 32508 12180 32564 12190
rect 32508 12086 32564 12124
rect 33068 12178 33124 12236
rect 33068 12126 33070 12178
rect 33122 12126 33124 12178
rect 33068 12114 33124 12126
rect 33516 12178 33572 12908
rect 33628 12516 33684 13580
rect 33740 13074 33796 14812
rect 33964 14420 34020 14924
rect 33964 14326 34020 14364
rect 34076 13858 34132 15148
rect 34076 13806 34078 13858
rect 34130 13806 34132 13858
rect 34076 13794 34132 13806
rect 34188 13748 34244 16606
rect 34748 16548 34804 16940
rect 34860 16772 34916 16782
rect 34860 16678 34916 16716
rect 34748 16492 34916 16548
rect 34300 15988 34356 15998
rect 34300 15894 34356 15932
rect 34412 15314 34468 15326
rect 34412 15262 34414 15314
rect 34466 15262 34468 15314
rect 34412 15204 34468 15262
rect 34636 15316 34692 15326
rect 34636 15204 34692 15260
rect 34412 15148 34692 15204
rect 34860 14756 34916 16492
rect 34972 15426 35028 17164
rect 35196 17106 35252 17390
rect 35196 17054 35198 17106
rect 35250 17054 35252 17106
rect 35196 17042 35252 17054
rect 35532 16884 35588 16894
rect 35308 16882 35588 16884
rect 35308 16830 35534 16882
rect 35586 16830 35588 16882
rect 35308 16828 35588 16830
rect 35308 16660 35364 16828
rect 35532 16818 35588 16828
rect 35756 16772 35812 16782
rect 35756 16678 35812 16716
rect 34972 15374 34974 15426
rect 35026 15374 35028 15426
rect 34972 14868 35028 15374
rect 34972 14802 35028 14812
rect 35084 16604 35364 16660
rect 35532 16660 35588 16670
rect 35084 14756 35140 16604
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35420 15652 35476 15662
rect 35308 15204 35364 15214
rect 35420 15204 35476 15596
rect 35308 15202 35476 15204
rect 35308 15150 35310 15202
rect 35362 15150 35476 15202
rect 35308 15148 35476 15150
rect 35532 15148 35588 16604
rect 35868 16098 35924 17500
rect 36092 17444 36148 17454
rect 35980 17442 36148 17444
rect 35980 17390 36094 17442
rect 36146 17390 36148 17442
rect 35980 17388 36148 17390
rect 35980 17220 36036 17388
rect 36092 17378 36148 17388
rect 35980 17154 36036 17164
rect 36092 17106 36148 17118
rect 36092 17054 36094 17106
rect 36146 17054 36148 17106
rect 35980 16996 36036 17006
rect 35980 16210 36036 16940
rect 36092 16884 36148 17054
rect 36316 16884 36372 16894
rect 36092 16882 36372 16884
rect 36092 16830 36318 16882
rect 36370 16830 36372 16882
rect 36092 16828 36372 16830
rect 36316 16818 36372 16828
rect 35980 16158 35982 16210
rect 36034 16158 36036 16210
rect 35980 16146 36036 16158
rect 35868 16046 35870 16098
rect 35922 16046 35924 16098
rect 35868 16034 35924 16046
rect 36316 16100 36372 16110
rect 36428 16100 36484 17948
rect 36764 17668 36820 22540
rect 36876 21700 36932 22878
rect 37212 22372 37268 26908
rect 37660 26962 37716 27468
rect 38444 27188 38500 27198
rect 38332 27132 38444 27188
rect 37660 26910 37662 26962
rect 37714 26910 37716 26962
rect 37660 26898 37716 26910
rect 37884 27074 37940 27086
rect 37884 27022 37886 27074
rect 37938 27022 37940 27074
rect 37324 26404 37380 26414
rect 37324 26310 37380 26348
rect 37436 26066 37492 26078
rect 37436 26014 37438 26066
rect 37490 26014 37492 26066
rect 37436 24724 37492 26014
rect 37436 23938 37492 24668
rect 37436 23886 37438 23938
rect 37490 23886 37492 23938
rect 37436 23874 37492 23886
rect 37884 24836 37940 27022
rect 37548 23828 37604 23838
rect 37324 23042 37380 23054
rect 37324 22990 37326 23042
rect 37378 22990 37380 23042
rect 37324 22932 37380 22990
rect 37324 22866 37380 22876
rect 37548 22596 37604 23772
rect 37884 23044 37940 24780
rect 38332 24276 38388 27132
rect 38444 27094 38500 27132
rect 38780 26908 38836 28812
rect 39116 28756 39172 30156
rect 39228 30146 39284 30156
rect 39452 29988 39508 29998
rect 39564 29988 39620 31612
rect 40236 31668 40292 31678
rect 39900 31556 39956 31566
rect 40236 31556 40292 31612
rect 39900 31554 40292 31556
rect 39900 31502 39902 31554
rect 39954 31502 40292 31554
rect 39900 31500 40292 31502
rect 39900 31490 39956 31500
rect 40236 30660 40292 31500
rect 40348 31220 40404 32172
rect 40796 31892 40852 45614
rect 40908 45220 40964 45230
rect 40908 45126 40964 45164
rect 41132 44100 41188 44110
rect 41132 42530 41188 44044
rect 41132 42478 41134 42530
rect 41186 42478 41188 42530
rect 41020 41972 41076 41982
rect 41132 41972 41188 42478
rect 41076 41916 41188 41972
rect 41356 43538 41412 45726
rect 41692 45778 41748 47180
rect 42364 47236 42420 47246
rect 42364 47142 42420 47180
rect 41804 47012 41860 47022
rect 41860 46956 41972 47012
rect 41804 46946 41860 46956
rect 41692 45726 41694 45778
rect 41746 45726 41748 45778
rect 41692 45714 41748 45726
rect 41916 45108 41972 46956
rect 43036 45892 43092 45902
rect 42476 45890 43092 45892
rect 42476 45838 43038 45890
rect 43090 45838 43092 45890
rect 42476 45836 43092 45838
rect 42028 45108 42084 45118
rect 41916 45106 42084 45108
rect 41916 45054 42030 45106
rect 42082 45054 42084 45106
rect 41916 45052 42084 45054
rect 41468 44996 41524 45006
rect 41468 44902 41524 44940
rect 41804 44436 41860 44446
rect 41916 44436 41972 45052
rect 42028 45042 42084 45052
rect 42476 44546 42532 45836
rect 43036 45826 43092 45836
rect 42812 45666 42868 45678
rect 42812 45614 42814 45666
rect 42866 45614 42868 45666
rect 42812 45106 42868 45614
rect 42812 45054 42814 45106
rect 42866 45054 42868 45106
rect 42812 45042 42868 45054
rect 42476 44494 42478 44546
rect 42530 44494 42532 44546
rect 42476 44482 42532 44494
rect 43036 44996 43092 45006
rect 41804 44434 41972 44436
rect 41804 44382 41806 44434
rect 41858 44382 41972 44434
rect 41804 44380 41972 44382
rect 41468 44212 41524 44222
rect 41468 43650 41524 44156
rect 41804 44100 41860 44380
rect 41804 44034 41860 44044
rect 42812 44322 42868 44334
rect 42812 44270 42814 44322
rect 42866 44270 42868 44322
rect 42812 43708 42868 44270
rect 43036 44212 43092 44940
rect 45164 44994 45220 45006
rect 45164 44942 45166 44994
rect 45218 44942 45220 44994
rect 43372 44212 43428 44222
rect 43036 44210 43316 44212
rect 43036 44158 43038 44210
rect 43090 44158 43316 44210
rect 43036 44156 43316 44158
rect 43036 44146 43092 44156
rect 43260 43708 43316 44156
rect 43372 44118 43428 44156
rect 45164 44212 45220 44942
rect 45164 44146 45220 44156
rect 42812 43652 42980 43708
rect 41468 43598 41470 43650
rect 41522 43598 41524 43650
rect 41468 43586 41524 43598
rect 41356 43486 41358 43538
rect 41410 43486 41412 43538
rect 41020 41878 41076 41916
rect 41356 40404 41412 43486
rect 42812 43538 42868 43550
rect 42812 43486 42814 43538
rect 42866 43486 42868 43538
rect 42028 43316 42084 43326
rect 42364 43316 42420 43326
rect 42028 43222 42084 43260
rect 42252 43314 42420 43316
rect 42252 43262 42366 43314
rect 42418 43262 42420 43314
rect 42252 43260 42420 43262
rect 41692 41972 41748 41982
rect 41692 40628 41748 41916
rect 42252 41188 42308 43260
rect 42364 43250 42420 43260
rect 42700 42980 42756 42990
rect 42812 42980 42868 43486
rect 42700 42978 42868 42980
rect 42700 42926 42702 42978
rect 42754 42926 42868 42978
rect 42700 42924 42868 42926
rect 42924 43316 42980 43652
rect 42700 42914 42756 42924
rect 42924 42196 42980 43260
rect 43148 43650 43204 43662
rect 43260 43652 43540 43708
rect 43148 43598 43150 43650
rect 43202 43598 43204 43650
rect 42924 42130 42980 42140
rect 43036 42754 43092 42766
rect 43036 42702 43038 42754
rect 43090 42702 43092 42754
rect 42364 41972 42420 41982
rect 42588 41972 42644 41982
rect 42420 41970 42644 41972
rect 42420 41918 42590 41970
rect 42642 41918 42644 41970
rect 42420 41916 42644 41918
rect 42364 41878 42420 41916
rect 42588 41906 42644 41916
rect 42252 41132 42532 41188
rect 41804 40964 41860 40974
rect 41804 40870 41860 40908
rect 42252 40962 42308 40974
rect 42252 40910 42254 40962
rect 42306 40910 42308 40962
rect 41692 40626 41972 40628
rect 41692 40574 41694 40626
rect 41746 40574 41972 40626
rect 41692 40572 41972 40574
rect 41692 40562 41748 40572
rect 41356 40338 41412 40348
rect 41916 40402 41972 40572
rect 41916 40350 41918 40402
rect 41970 40350 41972 40402
rect 41916 40338 41972 40350
rect 42252 39618 42308 40910
rect 42252 39566 42254 39618
rect 42306 39566 42308 39618
rect 42252 39554 42308 39566
rect 42364 40404 42420 40414
rect 41244 38946 41300 38958
rect 41244 38894 41246 38946
rect 41298 38894 41300 38946
rect 41020 38834 41076 38846
rect 41020 38782 41022 38834
rect 41074 38782 41076 38834
rect 41020 37492 41076 38782
rect 41244 38050 41300 38894
rect 41244 37998 41246 38050
rect 41298 37998 41300 38050
rect 41244 37986 41300 37998
rect 41468 37940 41524 37950
rect 41132 37492 41188 37502
rect 41020 37490 41188 37492
rect 41020 37438 41134 37490
rect 41186 37438 41188 37490
rect 41020 37436 41188 37438
rect 41132 37426 41188 37436
rect 41468 37266 41524 37884
rect 42252 37492 42308 37502
rect 42252 37380 42308 37436
rect 42028 37378 42308 37380
rect 42028 37326 42254 37378
rect 42306 37326 42308 37378
rect 42028 37324 42308 37326
rect 41468 37214 41470 37266
rect 41522 37214 41524 37266
rect 41468 37202 41524 37214
rect 41916 37266 41972 37278
rect 41916 37214 41918 37266
rect 41970 37214 41972 37266
rect 41916 37156 41972 37214
rect 41916 37090 41972 37100
rect 41916 35700 41972 35710
rect 42028 35700 42084 37324
rect 42252 37314 42308 37324
rect 42364 35700 42420 40348
rect 42476 38668 42532 41132
rect 42588 41186 42644 41198
rect 42588 41134 42590 41186
rect 42642 41134 42644 41186
rect 42588 40964 42644 41134
rect 42812 41076 42868 41086
rect 43036 41076 43092 42702
rect 43148 41972 43204 43598
rect 43484 42754 43540 43652
rect 43484 42702 43486 42754
rect 43538 42702 43540 42754
rect 43260 41972 43316 41982
rect 43148 41970 43316 41972
rect 43148 41918 43262 41970
rect 43314 41918 43316 41970
rect 43148 41916 43316 41918
rect 43260 41906 43316 41916
rect 43148 41076 43204 41086
rect 43036 41074 43204 41076
rect 43036 41022 43150 41074
rect 43202 41022 43204 41074
rect 43036 41020 43204 41022
rect 42812 40982 42868 41020
rect 42588 40898 42644 40908
rect 42588 40402 42644 40414
rect 42588 40350 42590 40402
rect 42642 40350 42644 40402
rect 42588 39506 42644 40350
rect 42588 39454 42590 39506
rect 42642 39454 42644 39506
rect 42588 39442 42644 39454
rect 42812 40404 42868 40414
rect 42476 38612 42644 38668
rect 41916 35698 42084 35700
rect 41916 35646 41918 35698
rect 41970 35646 42084 35698
rect 41916 35644 42084 35646
rect 42140 35698 42420 35700
rect 42140 35646 42366 35698
rect 42418 35646 42420 35698
rect 42140 35644 42420 35646
rect 41916 35634 41972 35644
rect 41244 35588 41300 35598
rect 41244 35586 41412 35588
rect 41244 35534 41246 35586
rect 41298 35534 41412 35586
rect 41244 35532 41412 35534
rect 41244 35522 41300 35532
rect 41356 35308 41412 35532
rect 41580 35476 41636 35486
rect 41580 35474 41748 35476
rect 41580 35422 41582 35474
rect 41634 35422 41748 35474
rect 41580 35420 41748 35422
rect 41580 35410 41636 35420
rect 41356 35252 41524 35308
rect 41244 34914 41300 34926
rect 41244 34862 41246 34914
rect 41298 34862 41300 34914
rect 41020 34356 41076 34366
rect 41020 34262 41076 34300
rect 41244 33572 41300 34862
rect 41244 33458 41300 33516
rect 41244 33406 41246 33458
rect 41298 33406 41300 33458
rect 41244 33394 41300 33406
rect 41468 34692 41524 35252
rect 41580 34692 41636 34702
rect 41468 34690 41636 34692
rect 41468 34638 41582 34690
rect 41634 34638 41636 34690
rect 41468 34636 41636 34638
rect 41356 32676 41412 32686
rect 41468 32676 41524 34636
rect 41580 34626 41636 34636
rect 41580 33908 41636 33918
rect 41580 33814 41636 33852
rect 41412 32620 41524 32676
rect 41580 32788 41636 32798
rect 41356 32610 41412 32620
rect 40908 32564 40964 32574
rect 40908 32470 40964 32508
rect 41244 32562 41300 32574
rect 41244 32510 41246 32562
rect 41298 32510 41300 32562
rect 40684 31836 40852 31892
rect 41132 32450 41188 32462
rect 41132 32398 41134 32450
rect 41186 32398 41188 32450
rect 40572 31780 40628 31818
rect 40572 31714 40628 31724
rect 40348 31154 40404 31164
rect 40460 31666 40516 31678
rect 40460 31614 40462 31666
rect 40514 31614 40516 31666
rect 40348 30884 40404 30894
rect 40348 30790 40404 30828
rect 40236 30604 40404 30660
rect 39452 29986 39620 29988
rect 39452 29934 39454 29986
rect 39506 29934 39620 29986
rect 39452 29932 39620 29934
rect 39452 29922 39508 29932
rect 39564 29538 39620 29932
rect 39564 29486 39566 29538
rect 39618 29486 39620 29538
rect 39564 29474 39620 29486
rect 39788 29428 39844 29438
rect 39788 29334 39844 29372
rect 39228 29316 39284 29326
rect 39228 29314 39396 29316
rect 39228 29262 39230 29314
rect 39282 29262 39396 29314
rect 39228 29260 39396 29262
rect 39228 29250 39284 29260
rect 38892 28644 38948 28654
rect 38892 28550 38948 28588
rect 39116 28642 39172 28700
rect 39116 28590 39118 28642
rect 39170 28590 39172 28642
rect 39116 28578 39172 28590
rect 39228 28530 39284 28542
rect 39228 28478 39230 28530
rect 39282 28478 39284 28530
rect 39228 28084 39284 28478
rect 39340 28532 39396 29260
rect 40124 29204 40180 29214
rect 40012 29202 40180 29204
rect 40012 29150 40126 29202
rect 40178 29150 40180 29202
rect 40012 29148 40180 29150
rect 39900 28644 39956 28654
rect 40012 28644 40068 29148
rect 40124 29138 40180 29148
rect 39900 28642 40068 28644
rect 39900 28590 39902 28642
rect 39954 28590 40068 28642
rect 39900 28588 40068 28590
rect 40236 28642 40292 28654
rect 40236 28590 40238 28642
rect 40290 28590 40292 28642
rect 39900 28578 39956 28588
rect 40236 28532 40292 28590
rect 39340 28466 39396 28476
rect 40124 28476 40236 28532
rect 39228 28018 39284 28028
rect 38892 27858 38948 27870
rect 38892 27806 38894 27858
rect 38946 27806 38948 27858
rect 38892 27636 38948 27806
rect 38892 27570 38948 27580
rect 39564 27746 39620 27758
rect 39564 27694 39566 27746
rect 39618 27694 39620 27746
rect 39564 27636 39620 27694
rect 38892 27300 38948 27310
rect 38892 27188 38948 27244
rect 38892 27186 39284 27188
rect 38892 27134 38894 27186
rect 38946 27134 39284 27186
rect 38892 27132 39284 27134
rect 38892 27122 38948 27132
rect 39228 27074 39284 27132
rect 39228 27022 39230 27074
rect 39282 27022 39284 27074
rect 39228 27010 39284 27022
rect 39452 27076 39508 27086
rect 39452 26982 39508 27020
rect 38780 26852 39284 26908
rect 39116 25396 39172 25406
rect 38668 25394 39172 25396
rect 38668 25342 39118 25394
rect 39170 25342 39172 25394
rect 38668 25340 39172 25342
rect 38556 24836 38612 24846
rect 38556 24742 38612 24780
rect 38332 24162 38388 24220
rect 38332 24110 38334 24162
rect 38386 24110 38388 24162
rect 37996 23828 38052 23838
rect 37996 23734 38052 23772
rect 37884 22978 37940 22988
rect 37996 23044 38052 23054
rect 38332 23044 38388 24110
rect 38444 24388 38500 24398
rect 38444 23716 38500 24332
rect 38668 24162 38724 25340
rect 39116 25330 39172 25340
rect 38780 24724 38836 24734
rect 38780 24630 38836 24668
rect 38668 24110 38670 24162
rect 38722 24110 38724 24162
rect 38668 24098 38724 24110
rect 39228 23940 39284 26852
rect 39564 26068 39620 27580
rect 39788 27412 39844 27422
rect 40012 27412 40068 27422
rect 39788 26964 39844 27356
rect 39900 27356 40012 27412
rect 39900 27074 39956 27356
rect 40012 27346 40068 27356
rect 39900 27022 39902 27074
rect 39954 27022 39956 27074
rect 39900 27010 39956 27022
rect 40124 27076 40180 28476
rect 40236 28466 40292 28476
rect 39676 26852 39732 26862
rect 39676 26758 39732 26796
rect 39788 26516 39844 26908
rect 40124 26962 40180 27020
rect 40124 26910 40126 26962
rect 40178 26910 40180 26962
rect 40124 26898 40180 26910
rect 40348 27748 40404 30604
rect 40460 30324 40516 31614
rect 40460 30258 40516 30268
rect 40572 31556 40628 31566
rect 40348 26908 40404 27692
rect 40572 26908 40628 31500
rect 40684 30210 40740 31836
rect 41020 31778 41076 31790
rect 41020 31726 41022 31778
rect 41074 31726 41076 31778
rect 40908 31668 40964 31678
rect 40908 31574 40964 31612
rect 40796 31220 40852 31230
rect 40852 31164 40964 31220
rect 40796 31154 40852 31164
rect 40908 31106 40964 31164
rect 41020 31218 41076 31726
rect 41132 31780 41188 32398
rect 41132 31714 41188 31724
rect 41020 31166 41022 31218
rect 41074 31166 41076 31218
rect 41020 31154 41076 31166
rect 41132 31220 41188 31230
rect 40908 31054 40910 31106
rect 40962 31054 40964 31106
rect 40908 31042 40964 31054
rect 41132 30436 41188 31164
rect 41020 30380 41188 30436
rect 40796 30324 40852 30334
rect 40796 30230 40852 30268
rect 40684 30158 40686 30210
rect 40738 30158 40740 30210
rect 40684 30146 40740 30158
rect 40908 30210 40964 30222
rect 40908 30158 40910 30210
rect 40962 30158 40964 30210
rect 40796 30100 40852 30110
rect 40796 28644 40852 30044
rect 40908 29764 40964 30158
rect 41020 30212 41076 30380
rect 41244 30324 41300 32510
rect 41356 31556 41412 31566
rect 41356 30994 41412 31500
rect 41356 30942 41358 30994
rect 41410 30942 41412 30994
rect 41356 30930 41412 30942
rect 41468 31106 41524 31118
rect 41468 31054 41470 31106
rect 41522 31054 41524 31106
rect 41468 30884 41524 31054
rect 41468 30818 41524 30828
rect 41580 30324 41636 32732
rect 41020 30146 41076 30156
rect 41132 30268 41300 30324
rect 41356 30268 41636 30324
rect 40908 29698 40964 29708
rect 40908 28644 40964 28654
rect 40796 28642 40964 28644
rect 40796 28590 40910 28642
rect 40962 28590 40964 28642
rect 40796 28588 40964 28590
rect 40908 27972 40964 28588
rect 41132 28532 41188 30268
rect 41244 30100 41300 30110
rect 41244 30006 41300 30044
rect 41244 29540 41300 29550
rect 41244 29446 41300 29484
rect 41132 28466 41188 28476
rect 40908 27906 40964 27916
rect 41020 28418 41076 28430
rect 41020 28366 41022 28418
rect 41074 28366 41076 28418
rect 41020 27860 41076 28366
rect 41020 27794 41076 27804
rect 41132 27858 41188 27870
rect 41132 27806 41134 27858
rect 41186 27806 41188 27858
rect 40684 27300 40740 27310
rect 40684 27074 40740 27244
rect 40684 27022 40686 27074
rect 40738 27022 40740 27074
rect 40684 27010 40740 27022
rect 40236 26852 40404 26908
rect 40460 26852 40628 26908
rect 40908 26852 40964 26862
rect 39900 26516 39956 26526
rect 39788 26514 39956 26516
rect 39788 26462 39902 26514
rect 39954 26462 39956 26514
rect 39788 26460 39956 26462
rect 39900 26450 39956 26460
rect 40236 26292 40292 26852
rect 40348 26740 40404 26750
rect 40348 26514 40404 26684
rect 40348 26462 40350 26514
rect 40402 26462 40404 26514
rect 40348 26450 40404 26462
rect 40236 26226 40292 26236
rect 39564 26012 39956 26068
rect 39900 25506 39956 26012
rect 39900 25454 39902 25506
rect 39954 25454 39956 25506
rect 39900 25284 39956 25454
rect 40348 25284 40404 25294
rect 39900 25282 40404 25284
rect 39900 25230 40350 25282
rect 40402 25230 40404 25282
rect 39900 25228 40404 25230
rect 38780 23938 39284 23940
rect 38780 23886 39230 23938
rect 39282 23886 39284 23938
rect 38780 23884 39284 23886
rect 38556 23828 38612 23838
rect 38556 23734 38612 23772
rect 38444 23650 38500 23660
rect 38780 23380 38836 23884
rect 39228 23874 39284 23884
rect 39340 24612 39396 24622
rect 38780 23286 38836 23324
rect 37996 23042 38388 23044
rect 37996 22990 37998 23042
rect 38050 22990 38388 23042
rect 37996 22988 38388 22990
rect 37996 22708 38052 22988
rect 37996 22642 38052 22652
rect 37548 22540 37940 22596
rect 37548 22482 37604 22540
rect 37548 22430 37550 22482
rect 37602 22430 37604 22482
rect 37548 22418 37604 22430
rect 37772 22372 37828 22382
rect 36876 21634 36932 21644
rect 36988 22316 37268 22372
rect 37660 22370 37828 22372
rect 37660 22318 37774 22370
rect 37826 22318 37828 22370
rect 37660 22316 37828 22318
rect 36988 21588 37044 22316
rect 37100 22146 37156 22158
rect 37100 22094 37102 22146
rect 37154 22094 37156 22146
rect 37100 21810 37156 22094
rect 37212 22146 37268 22158
rect 37212 22094 37214 22146
rect 37266 22094 37268 22146
rect 37212 21924 37268 22094
rect 37212 21858 37268 21868
rect 37324 22146 37380 22158
rect 37324 22094 37326 22146
rect 37378 22094 37380 22146
rect 37100 21758 37102 21810
rect 37154 21758 37156 21810
rect 37100 21746 37156 21758
rect 36988 21532 37156 21588
rect 36876 21476 36932 21486
rect 36932 21420 37044 21476
rect 36876 21410 36932 21420
rect 36988 20914 37044 21420
rect 36988 20862 36990 20914
rect 37042 20862 37044 20914
rect 36988 20850 37044 20862
rect 37100 20804 37156 21532
rect 37212 21364 37268 21374
rect 37212 21270 37268 21308
rect 37324 21028 37380 22094
rect 37436 21588 37492 21598
rect 37436 21494 37492 21532
rect 37324 20972 37492 21028
rect 37324 20804 37380 20814
rect 37100 20802 37380 20804
rect 37100 20750 37326 20802
rect 37378 20750 37380 20802
rect 37100 20748 37380 20750
rect 37100 19684 37156 20748
rect 37324 20738 37380 20748
rect 37100 19628 37380 19684
rect 37100 19234 37156 19628
rect 37100 19182 37102 19234
rect 37154 19182 37156 19234
rect 37100 19170 37156 19182
rect 37212 19458 37268 19470
rect 37212 19406 37214 19458
rect 37266 19406 37268 19458
rect 37212 18788 37268 19406
rect 37100 18732 37268 18788
rect 36988 18562 37044 18574
rect 36988 18510 36990 18562
rect 37042 18510 37044 18562
rect 36988 18452 37044 18510
rect 36988 18386 37044 18396
rect 37100 18228 37156 18732
rect 36652 17612 36820 17668
rect 36876 18172 37156 18228
rect 36652 17220 36708 17612
rect 36652 16660 36708 17164
rect 36764 17444 36820 17454
rect 36764 16884 36820 17388
rect 36876 16996 36932 18172
rect 37100 18116 37156 18172
rect 37100 18050 37156 18060
rect 37212 18564 37268 18574
rect 37212 18450 37268 18508
rect 37212 18398 37214 18450
rect 37266 18398 37268 18450
rect 37212 18004 37268 18398
rect 37324 18452 37380 19628
rect 37436 18674 37492 20972
rect 37660 19346 37716 22316
rect 37772 22306 37828 22316
rect 37772 21700 37828 21710
rect 37884 21700 37940 22540
rect 37996 22372 38052 22382
rect 37996 22370 38388 22372
rect 37996 22318 37998 22370
rect 38050 22318 38388 22370
rect 37996 22316 38388 22318
rect 37996 22306 38052 22316
rect 37996 21700 38052 21710
rect 37884 21698 38052 21700
rect 37884 21646 37998 21698
rect 38050 21646 38052 21698
rect 37884 21644 38052 21646
rect 37772 21606 37828 21644
rect 37996 21634 38052 21644
rect 38332 21698 38388 22316
rect 39004 22148 39060 22158
rect 38332 21646 38334 21698
rect 38386 21646 38388 21698
rect 38332 21634 38388 21646
rect 38444 21700 38500 21710
rect 38444 21586 38500 21644
rect 38444 21534 38446 21586
rect 38498 21534 38500 21586
rect 38444 21522 38500 21534
rect 38668 21588 38724 21598
rect 38668 21494 38724 21532
rect 38780 21362 38836 21374
rect 38780 21310 38782 21362
rect 38834 21310 38836 21362
rect 38780 21252 38836 21310
rect 37884 20804 37940 20814
rect 37884 20802 38276 20804
rect 37884 20750 37886 20802
rect 37938 20750 38276 20802
rect 37884 20748 38276 20750
rect 37884 20738 37940 20748
rect 37996 20580 38052 20590
rect 37996 20486 38052 20524
rect 38108 20020 38164 20030
rect 38108 19926 38164 19964
rect 37996 19684 38052 19694
rect 38052 19628 38164 19684
rect 37996 19618 38052 19628
rect 37660 19294 37662 19346
rect 37714 19294 37716 19346
rect 37660 19282 37716 19294
rect 37548 19236 37604 19246
rect 37548 19142 37604 19180
rect 37772 19122 37828 19134
rect 37772 19070 37774 19122
rect 37826 19070 37828 19122
rect 37436 18622 37438 18674
rect 37490 18622 37492 18674
rect 37436 18610 37492 18622
rect 37660 18788 37716 18798
rect 37548 18452 37604 18462
rect 37324 18450 37604 18452
rect 37324 18398 37550 18450
rect 37602 18398 37604 18450
rect 37324 18396 37604 18398
rect 37548 18386 37604 18396
rect 37436 18226 37492 18238
rect 37436 18174 37438 18226
rect 37490 18174 37492 18226
rect 37436 18004 37492 18174
rect 37212 17948 37380 18004
rect 37212 17780 37268 17790
rect 37212 17686 37268 17724
rect 36988 17556 37044 17566
rect 36988 17106 37044 17500
rect 36988 17054 36990 17106
rect 37042 17054 37044 17106
rect 36988 17042 37044 17054
rect 36876 16930 36932 16940
rect 37100 16996 37156 17006
rect 36764 16790 36820 16828
rect 36876 16772 36932 16782
rect 36876 16678 36932 16716
rect 36652 16594 36708 16604
rect 37100 16436 37156 16940
rect 37324 16884 37380 17948
rect 37436 17938 37492 17948
rect 37436 17668 37492 17678
rect 37436 17220 37492 17612
rect 37436 17106 37492 17164
rect 37436 17054 37438 17106
rect 37490 17054 37492 17106
rect 37436 17042 37492 17054
rect 37660 17108 37716 18732
rect 37772 18452 37828 19070
rect 37772 18386 37828 18396
rect 37996 18450 38052 18462
rect 37996 18398 37998 18450
rect 38050 18398 38052 18450
rect 37996 18340 38052 18398
rect 37884 18284 37996 18340
rect 37660 17014 37716 17052
rect 37772 17108 37828 17118
rect 37884 17108 37940 18284
rect 37996 18274 38052 18284
rect 38108 17892 38164 19628
rect 38220 18450 38276 20748
rect 38444 20692 38500 20702
rect 38444 20598 38500 20636
rect 38556 20132 38724 20188
rect 38556 19906 38612 20132
rect 38668 20066 38724 20076
rect 38556 19854 38558 19906
rect 38610 19854 38612 19906
rect 38220 18398 38222 18450
rect 38274 18398 38276 18450
rect 38220 18386 38276 18398
rect 38332 19236 38388 19246
rect 38332 18450 38388 19180
rect 38556 19236 38612 19854
rect 38444 19124 38500 19134
rect 38444 18676 38500 19068
rect 38444 18610 38500 18620
rect 38332 18398 38334 18450
rect 38386 18398 38388 18450
rect 38332 18228 38388 18398
rect 38332 18162 38388 18172
rect 37772 17106 37940 17108
rect 37772 17054 37774 17106
rect 37826 17054 37940 17106
rect 37772 17052 37940 17054
rect 37996 17836 38164 17892
rect 37772 17042 37828 17052
rect 37100 16370 37156 16380
rect 37212 16828 37380 16884
rect 37884 16884 37940 16894
rect 37996 16884 38052 17836
rect 37884 16882 38052 16884
rect 37884 16830 37886 16882
rect 37938 16830 38052 16882
rect 37884 16828 38052 16830
rect 36988 16212 37044 16222
rect 36372 16044 36484 16100
rect 36540 16210 37044 16212
rect 36540 16158 36990 16210
rect 37042 16158 37044 16210
rect 36540 16156 37044 16158
rect 36540 16098 36596 16156
rect 36988 16146 37044 16156
rect 36540 16046 36542 16098
rect 36594 16046 36596 16098
rect 36316 16034 36372 16044
rect 36540 16034 36596 16046
rect 36092 15988 36148 15998
rect 36092 15894 36148 15932
rect 36988 15988 37044 15998
rect 36540 15876 36596 15886
rect 35756 15596 36260 15652
rect 35756 15314 35812 15596
rect 36204 15538 36260 15596
rect 36204 15486 36206 15538
rect 36258 15486 36260 15538
rect 36204 15474 36260 15486
rect 36316 15540 36372 15550
rect 36540 15540 36596 15820
rect 36988 15540 37044 15932
rect 36316 15538 36596 15540
rect 36316 15486 36318 15538
rect 36370 15486 36596 15538
rect 36316 15484 36596 15486
rect 36876 15484 37044 15540
rect 37100 15764 37156 15774
rect 36316 15474 36372 15484
rect 35756 15262 35758 15314
rect 35810 15262 35812 15314
rect 35756 15250 35812 15262
rect 36092 15314 36148 15326
rect 36092 15262 36094 15314
rect 36146 15262 36148 15314
rect 35308 15138 35364 15148
rect 35532 15092 35812 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35084 14700 35364 14756
rect 34860 14690 34916 14700
rect 35196 14420 35252 14430
rect 34524 13972 34580 13982
rect 34524 13878 34580 13916
rect 34972 13972 35028 13982
rect 35028 13916 35140 13972
rect 34972 13906 35028 13916
rect 34860 13860 34916 13870
rect 34860 13766 34916 13804
rect 34188 13682 34244 13692
rect 33740 13022 33742 13074
rect 33794 13022 33796 13074
rect 33740 13010 33796 13022
rect 33852 13076 33908 13086
rect 34076 13076 34132 13086
rect 33852 12962 33908 13020
rect 33852 12910 33854 12962
rect 33906 12910 33908 12962
rect 33852 12898 33908 12910
rect 33964 13074 34132 13076
rect 33964 13022 34078 13074
rect 34130 13022 34132 13074
rect 33964 13020 34132 13022
rect 33628 12450 33684 12460
rect 33516 12126 33518 12178
rect 33570 12126 33572 12178
rect 33516 12114 33572 12126
rect 32620 12068 32676 12078
rect 32620 12066 33012 12068
rect 32620 12014 32622 12066
rect 32674 12014 33012 12066
rect 32620 12012 33012 12014
rect 32620 12002 32676 12012
rect 32508 11732 32564 11742
rect 32564 11676 32676 11732
rect 32508 11666 32564 11676
rect 32620 11394 32676 11676
rect 32620 11342 32622 11394
rect 32674 11342 32676 11394
rect 32620 11330 32676 11342
rect 32956 11396 33012 12012
rect 32956 11340 33236 11396
rect 32508 11284 32564 11294
rect 32396 11282 32564 11284
rect 32396 11230 32510 11282
rect 32562 11230 32564 11282
rect 32396 11228 32564 11230
rect 32396 9826 32452 11228
rect 32508 11218 32564 11228
rect 33180 10722 33236 11340
rect 33964 11284 34020 13020
rect 34076 13010 34132 13020
rect 34972 13074 35028 13086
rect 34972 13022 34974 13074
rect 35026 13022 35028 13074
rect 34972 12964 35028 13022
rect 34972 12898 35028 12908
rect 34188 12852 34244 12862
rect 34188 12758 34244 12796
rect 34412 12852 34468 12862
rect 34412 12758 34468 12796
rect 34860 12852 34916 12862
rect 35084 12852 35140 13916
rect 35196 13858 35252 14364
rect 35196 13806 35198 13858
rect 35250 13806 35252 13858
rect 35196 13794 35252 13806
rect 35308 13524 35364 14700
rect 35644 14644 35700 14654
rect 35644 14550 35700 14588
rect 35308 13458 35364 13468
rect 35532 14418 35588 14430
rect 35532 14366 35534 14418
rect 35586 14366 35588 14418
rect 35532 13860 35588 14366
rect 35756 14084 35812 15092
rect 36092 14980 36148 15262
rect 36652 15316 36708 15354
rect 36652 15250 36708 15260
rect 36876 15148 36932 15484
rect 36988 15316 37044 15326
rect 37100 15316 37156 15708
rect 37212 15428 37268 16828
rect 37884 16818 37940 16828
rect 37324 16660 37380 16670
rect 37324 16324 37380 16604
rect 37324 16322 37716 16324
rect 37324 16270 37326 16322
rect 37378 16270 37716 16322
rect 37324 16268 37716 16270
rect 37324 16258 37380 16268
rect 37548 15986 37604 15998
rect 37548 15934 37550 15986
rect 37602 15934 37604 15986
rect 37548 15540 37604 15934
rect 37548 15474 37604 15484
rect 37436 15428 37492 15438
rect 37212 15362 37268 15372
rect 37324 15372 37436 15428
rect 36988 15314 37156 15316
rect 36988 15262 36990 15314
rect 37042 15262 37156 15314
rect 36988 15260 37156 15262
rect 36988 15250 37044 15260
rect 37324 15148 37380 15372
rect 37436 15362 37492 15372
rect 37548 15316 37604 15326
rect 37548 15222 37604 15260
rect 36876 15092 37156 15148
rect 36092 14914 36148 14924
rect 36204 14868 36260 14878
rect 36204 14642 36260 14812
rect 36204 14590 36206 14642
rect 36258 14590 36260 14642
rect 36204 14578 36260 14590
rect 36988 14756 37044 14766
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 13076 35252 13086
rect 35196 12982 35252 13020
rect 35532 12962 35588 13804
rect 35532 12910 35534 12962
rect 35586 12910 35588 12962
rect 35532 12898 35588 12910
rect 35644 14028 35812 14084
rect 35980 14532 36036 14542
rect 35084 12796 35476 12852
rect 34524 12740 34580 12750
rect 33628 11228 34020 11284
rect 34076 12516 34132 12526
rect 33292 10836 33348 10846
rect 33292 10834 33572 10836
rect 33292 10782 33294 10834
rect 33346 10782 33572 10834
rect 33292 10780 33572 10782
rect 33292 10770 33348 10780
rect 33180 10670 33182 10722
rect 33234 10670 33236 10722
rect 33180 10658 33236 10670
rect 32396 9774 32398 9826
rect 32450 9774 32452 9826
rect 32396 9762 32452 9774
rect 33068 10052 33124 10062
rect 33068 9826 33124 9996
rect 33068 9774 33070 9826
rect 33122 9774 33124 9826
rect 33068 9762 33124 9774
rect 33180 9828 33236 9838
rect 33404 9828 33460 9838
rect 33180 9826 33460 9828
rect 33180 9774 33182 9826
rect 33234 9774 33406 9826
rect 33458 9774 33460 9826
rect 33180 9772 33460 9774
rect 33180 9762 33236 9772
rect 33404 9762 33460 9772
rect 32844 9716 32900 9726
rect 32844 9622 32900 9660
rect 32620 9604 32676 9614
rect 33516 9604 33572 10780
rect 33628 10050 33684 11228
rect 34076 11172 34132 12460
rect 34412 12516 34468 12526
rect 34300 12180 34356 12190
rect 34300 12086 34356 12124
rect 34412 11788 34468 12460
rect 34524 12180 34580 12684
rect 34524 12086 34580 12124
rect 34860 12178 34916 12796
rect 35420 12402 35476 12796
rect 35420 12350 35422 12402
rect 35474 12350 35476 12402
rect 35420 12338 35476 12350
rect 34860 12126 34862 12178
rect 34914 12126 34916 12178
rect 34860 12114 34916 12126
rect 34860 11956 34916 11966
rect 35196 11956 35252 11966
rect 34412 11732 34692 11788
rect 34636 11620 34692 11732
rect 34636 11554 34692 11564
rect 34524 11284 34580 11294
rect 33628 9998 33630 10050
rect 33682 9998 33684 10050
rect 33628 9986 33684 9998
rect 33852 11116 34132 11172
rect 34412 11282 34580 11284
rect 34412 11230 34526 11282
rect 34578 11230 34580 11282
rect 34412 11228 34580 11230
rect 33852 10050 33908 11116
rect 33852 9998 33854 10050
rect 33906 9998 33908 10050
rect 33852 9828 33908 9998
rect 33852 9762 33908 9772
rect 32620 9510 32676 9548
rect 33404 9548 33572 9604
rect 33964 9714 34020 9726
rect 33964 9662 33966 9714
rect 34018 9662 34020 9714
rect 32284 9426 32340 9436
rect 31836 8206 31838 8258
rect 31890 8206 31892 8258
rect 31836 8194 31892 8206
rect 32060 9324 32228 9380
rect 31500 7422 31502 7474
rect 31554 7422 31556 7474
rect 31500 7410 31556 7422
rect 31276 6750 31278 6802
rect 31330 6750 31332 6802
rect 31276 6738 31332 6750
rect 31948 6690 32004 6702
rect 31948 6638 31950 6690
rect 32002 6638 32004 6690
rect 30156 6580 30212 6590
rect 30492 6580 30548 6590
rect 30156 6578 30548 6580
rect 30156 6526 30158 6578
rect 30210 6526 30494 6578
rect 30546 6526 30548 6578
rect 30156 6524 30548 6526
rect 30156 6514 30212 6524
rect 30492 6514 30548 6524
rect 29820 6020 29876 6412
rect 30828 6468 30884 6478
rect 30828 6466 31220 6468
rect 30828 6414 30830 6466
rect 30882 6414 31220 6466
rect 30828 6412 31220 6414
rect 30828 6402 30884 6412
rect 31164 6132 31220 6412
rect 31164 6076 31780 6132
rect 31052 6020 31108 6030
rect 29820 5964 30324 6020
rect 30044 5236 30100 5246
rect 30044 5122 30100 5180
rect 30044 5070 30046 5122
rect 30098 5070 30100 5122
rect 30044 5058 30100 5070
rect 29652 4956 29764 5012
rect 30268 5010 30324 5964
rect 31052 5346 31108 5964
rect 31724 6018 31780 6076
rect 31724 5966 31726 6018
rect 31778 5966 31780 6018
rect 31724 5954 31780 5966
rect 31948 5908 32004 6638
rect 32060 6356 32116 9324
rect 32172 9154 32228 9166
rect 32172 9102 32174 9154
rect 32226 9102 32228 9154
rect 32172 8372 32228 9102
rect 32284 9042 32340 9054
rect 32284 8990 32286 9042
rect 32338 8990 32340 9042
rect 32284 8932 32340 8990
rect 33404 9044 33460 9548
rect 33964 9268 34020 9662
rect 33628 9212 34020 9268
rect 34076 9716 34132 9726
rect 33628 9154 33684 9212
rect 33628 9102 33630 9154
rect 33682 9102 33684 9154
rect 33628 9090 33684 9102
rect 33404 8950 33460 8988
rect 34076 9042 34132 9660
rect 34300 9602 34356 9614
rect 34300 9550 34302 9602
rect 34354 9550 34356 9602
rect 34300 9492 34356 9550
rect 34300 9426 34356 9436
rect 34300 9268 34356 9278
rect 34412 9268 34468 11228
rect 34524 11218 34580 11228
rect 34300 9266 34468 9268
rect 34300 9214 34302 9266
rect 34354 9214 34468 9266
rect 34300 9212 34468 9214
rect 34524 11060 34580 11070
rect 34300 9202 34356 9212
rect 34076 8990 34078 9042
rect 34130 8990 34132 9042
rect 32284 8866 32340 8876
rect 33068 8932 33124 8942
rect 33068 8838 33124 8876
rect 32172 8148 32228 8316
rect 33292 8484 33348 8494
rect 32396 8148 32452 8158
rect 32172 8146 32452 8148
rect 32172 8094 32398 8146
rect 32450 8094 32452 8146
rect 32172 8092 32452 8094
rect 32396 8082 32452 8092
rect 32508 7700 32564 7710
rect 32060 6290 32116 6300
rect 32172 7586 32228 7598
rect 32172 7534 32174 7586
rect 32226 7534 32228 7586
rect 32172 6132 32228 7534
rect 32508 7476 32564 7644
rect 33292 7698 33348 8428
rect 34076 8484 34132 8990
rect 34076 8372 34132 8428
rect 34412 8818 34468 8830
rect 34412 8766 34414 8818
rect 34466 8766 34468 8818
rect 34412 8484 34468 8766
rect 34412 8418 34468 8428
rect 34524 8372 34580 11004
rect 34636 10948 34692 10958
rect 34636 10610 34692 10892
rect 34636 10558 34638 10610
rect 34690 10558 34692 10610
rect 34636 10546 34692 10558
rect 34860 10276 34916 11900
rect 35084 11900 35196 11956
rect 34748 10220 34916 10276
rect 34972 11620 35028 11630
rect 34636 9604 34692 9614
rect 34636 9510 34692 9548
rect 34748 8484 34804 10220
rect 34860 10052 34916 10062
rect 34860 9266 34916 9996
rect 34860 9214 34862 9266
rect 34914 9214 34916 9266
rect 34860 9202 34916 9214
rect 34748 8428 34916 8484
rect 34076 8370 34356 8372
rect 34076 8318 34078 8370
rect 34130 8318 34356 8370
rect 34076 8316 34356 8318
rect 34524 8316 34804 8372
rect 34076 8306 34132 8316
rect 34300 8260 34356 8316
rect 34748 8260 34804 8316
rect 34300 8204 34692 8260
rect 33292 7646 33294 7698
rect 33346 7646 33348 7698
rect 33292 7634 33348 7646
rect 34636 7698 34692 8204
rect 34748 8166 34804 8204
rect 34636 7646 34638 7698
rect 34690 7646 34692 7698
rect 34636 7634 34692 7646
rect 34076 7588 34132 7598
rect 34076 7494 34132 7532
rect 32508 7410 32564 7420
rect 33628 7362 33684 7374
rect 33628 7310 33630 7362
rect 33682 7310 33684 7362
rect 32620 6692 32676 6702
rect 32620 6598 32676 6636
rect 32172 6066 32228 6076
rect 33516 6468 33572 6478
rect 31948 5842 32004 5852
rect 32508 5908 32564 5918
rect 32508 5814 32564 5852
rect 33516 5906 33572 6412
rect 33516 5854 33518 5906
rect 33570 5854 33572 5906
rect 33516 5842 33572 5854
rect 31052 5294 31054 5346
rect 31106 5294 31108 5346
rect 31052 5282 31108 5294
rect 31724 5684 31780 5694
rect 31724 5234 31780 5628
rect 31724 5182 31726 5234
rect 31778 5182 31780 5234
rect 31724 5170 31780 5182
rect 30828 5124 30884 5134
rect 30828 5030 30884 5068
rect 33628 5124 33684 7310
rect 34748 6804 34804 6814
rect 34860 6804 34916 8428
rect 34972 7700 35028 11564
rect 35084 11394 35140 11900
rect 35196 11890 35252 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35420 11508 35476 11518
rect 35420 11414 35476 11452
rect 35084 11342 35086 11394
rect 35138 11342 35140 11394
rect 35084 11330 35140 11342
rect 35532 11396 35588 11406
rect 35644 11396 35700 14028
rect 35756 13746 35812 13758
rect 35756 13694 35758 13746
rect 35810 13694 35812 13746
rect 35756 13076 35812 13694
rect 35756 13010 35812 13020
rect 35868 12852 35924 12862
rect 35868 12758 35924 12796
rect 35532 11394 35700 11396
rect 35532 11342 35534 11394
rect 35586 11342 35700 11394
rect 35532 11340 35700 11342
rect 35756 12178 35812 12190
rect 35756 12126 35758 12178
rect 35810 12126 35812 12178
rect 35532 11284 35588 11340
rect 35308 11228 35588 11284
rect 35084 10948 35140 10958
rect 35084 9938 35140 10892
rect 35196 10612 35252 10622
rect 35308 10612 35364 11228
rect 35196 10610 35364 10612
rect 35196 10558 35198 10610
rect 35250 10558 35364 10610
rect 35196 10556 35364 10558
rect 35532 10836 35588 10846
rect 35196 10546 35252 10556
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35532 10052 35588 10780
rect 35084 9886 35086 9938
rect 35138 9886 35140 9938
rect 35084 9874 35140 9886
rect 35420 9996 35588 10052
rect 35644 10722 35700 10734
rect 35644 10670 35646 10722
rect 35698 10670 35700 10722
rect 35420 9156 35476 9996
rect 35532 9828 35588 9838
rect 35532 9380 35588 9772
rect 35644 9716 35700 10670
rect 35756 9940 35812 12126
rect 35756 9874 35812 9884
rect 35868 10052 35924 10062
rect 35868 9938 35924 9996
rect 35868 9886 35870 9938
rect 35922 9886 35924 9938
rect 35868 9874 35924 9886
rect 35644 9650 35700 9660
rect 35532 9314 35588 9324
rect 35420 9100 35588 9156
rect 35420 8930 35476 8942
rect 35420 8878 35422 8930
rect 35474 8878 35476 8930
rect 35420 8820 35476 8878
rect 35420 8754 35476 8764
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 8370 35252 8382
rect 35196 8318 35198 8370
rect 35250 8318 35252 8370
rect 35196 8148 35252 8318
rect 35196 8082 35252 8092
rect 34972 7606 35028 7644
rect 35532 7700 35588 9100
rect 35756 8260 35812 8270
rect 35756 8166 35812 8204
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35532 6914 35588 7644
rect 35868 7700 35924 7710
rect 35980 7700 36036 14476
rect 36092 14420 36148 14430
rect 36092 13970 36148 14364
rect 36988 14418 37044 14700
rect 36988 14366 36990 14418
rect 37042 14366 37044 14418
rect 36988 14354 37044 14366
rect 36092 13918 36094 13970
rect 36146 13918 36148 13970
rect 36092 13906 36148 13918
rect 36876 14306 36932 14318
rect 36876 14254 36878 14306
rect 36930 14254 36932 14306
rect 36316 13748 36372 13758
rect 36876 13748 36932 14254
rect 36988 13972 37044 13982
rect 37100 13972 37156 15092
rect 37212 15092 37380 15148
rect 37436 15204 37492 15214
rect 37212 15090 37268 15092
rect 37212 15038 37214 15090
rect 37266 15038 37268 15090
rect 37212 15026 37268 15038
rect 37436 14530 37492 15148
rect 37436 14478 37438 14530
rect 37490 14478 37492 14530
rect 37436 14466 37492 14478
rect 37212 14308 37268 14318
rect 37212 14306 37492 14308
rect 37212 14254 37214 14306
rect 37266 14254 37492 14306
rect 37212 14252 37492 14254
rect 37212 14242 37268 14252
rect 36988 13970 37156 13972
rect 36988 13918 36990 13970
rect 37042 13918 37156 13970
rect 36988 13916 37156 13918
rect 37212 14084 37268 14094
rect 36988 13906 37044 13916
rect 36876 13692 37156 13748
rect 36316 13074 36372 13692
rect 36540 13636 36596 13646
rect 36540 13542 36596 13580
rect 36316 13022 36318 13074
rect 36370 13022 36372 13074
rect 36316 12628 36372 13022
rect 36316 12562 36372 12572
rect 36428 12852 36484 12862
rect 36092 12404 36148 12414
rect 36092 12178 36148 12348
rect 36428 12180 36484 12796
rect 36092 12126 36094 12178
rect 36146 12126 36148 12178
rect 36092 12114 36148 12126
rect 36316 12124 36484 12180
rect 36092 11956 36148 11966
rect 36092 11862 36148 11900
rect 36204 11284 36260 11294
rect 36316 11284 36372 12124
rect 36204 11282 36372 11284
rect 36204 11230 36206 11282
rect 36258 11230 36372 11282
rect 36204 11228 36372 11230
rect 36428 11954 36484 11966
rect 36428 11902 36430 11954
rect 36482 11902 36484 11954
rect 36204 11218 36260 11228
rect 36092 9940 36148 9950
rect 36092 9714 36148 9884
rect 36092 9662 36094 9714
rect 36146 9662 36148 9714
rect 36092 9650 36148 9662
rect 36428 8708 36484 11902
rect 36988 11394 37044 11406
rect 36988 11342 36990 11394
rect 37042 11342 37044 11394
rect 36988 10052 37044 11342
rect 37100 10724 37156 13692
rect 37212 11396 37268 14028
rect 37212 11302 37268 11340
rect 37324 13748 37380 13758
rect 37324 12850 37380 13692
rect 37324 12798 37326 12850
rect 37378 12798 37380 12850
rect 37324 11172 37380 12798
rect 37436 12852 37492 14252
rect 37660 13972 37716 16268
rect 37996 15540 38052 16828
rect 38108 17668 38164 17678
rect 38108 16210 38164 17612
rect 38556 17668 38612 19180
rect 38668 18450 38724 18462
rect 38668 18398 38670 18450
rect 38722 18398 38724 18450
rect 38668 18004 38724 18398
rect 38668 17938 38724 17948
rect 38556 17602 38612 17612
rect 38220 17108 38276 17118
rect 38220 17014 38276 17052
rect 38556 16994 38612 17006
rect 38556 16942 38558 16994
rect 38610 16942 38612 16994
rect 38444 16772 38500 16782
rect 38108 16158 38110 16210
rect 38162 16158 38164 16210
rect 38108 16146 38164 16158
rect 38220 16660 38276 16670
rect 37996 15474 38052 15484
rect 37884 15316 37940 15354
rect 37884 15250 37940 15260
rect 38108 15202 38164 15214
rect 38108 15150 38110 15202
rect 38162 15150 38164 15202
rect 38108 15148 38164 15150
rect 38220 15148 38276 16604
rect 38444 16098 38500 16716
rect 38444 16046 38446 16098
rect 38498 16046 38500 16098
rect 38444 16034 38500 16046
rect 38556 16436 38612 16942
rect 38780 16548 38836 21196
rect 39004 20132 39060 22092
rect 39340 21924 39396 24556
rect 39788 24164 39844 24174
rect 39452 23940 39508 23950
rect 39452 23548 39508 23884
rect 39676 23826 39732 23838
rect 39676 23774 39678 23826
rect 39730 23774 39732 23826
rect 39676 23604 39732 23774
rect 39452 23492 39620 23548
rect 39676 23538 39732 23548
rect 39564 22372 39620 23492
rect 39676 23044 39732 23054
rect 39788 23044 39844 24108
rect 39900 23940 39956 25228
rect 40348 25218 40404 25228
rect 40348 24948 40404 24958
rect 40460 24948 40516 26852
rect 40796 26514 40852 26526
rect 40796 26462 40798 26514
rect 40850 26462 40852 26514
rect 40796 25956 40852 26462
rect 40908 26290 40964 26796
rect 41132 26850 41188 27806
rect 41244 27076 41300 27086
rect 41356 27076 41412 30268
rect 41580 30098 41636 30110
rect 41580 30046 41582 30098
rect 41634 30046 41636 30098
rect 41580 29540 41636 30046
rect 41580 29474 41636 29484
rect 41692 28642 41748 35420
rect 42140 35026 42196 35644
rect 42364 35634 42420 35644
rect 42140 34974 42142 35026
rect 42194 34974 42196 35026
rect 42140 34242 42196 34974
rect 42476 34692 42532 34702
rect 42476 34598 42532 34636
rect 42140 34190 42142 34242
rect 42194 34190 42196 34242
rect 42140 34178 42196 34190
rect 42476 34356 42532 34366
rect 42140 34020 42196 34030
rect 41916 33906 41972 33918
rect 41916 33854 41918 33906
rect 41970 33854 41972 33906
rect 41916 33796 41972 33854
rect 41916 33740 42084 33796
rect 41916 33572 41972 33582
rect 41804 33516 41916 33572
rect 41804 32004 41860 33516
rect 41916 33506 41972 33516
rect 42028 33348 42084 33740
rect 42028 33282 42084 33292
rect 42140 33346 42196 33964
rect 42140 33294 42142 33346
rect 42194 33294 42196 33346
rect 42140 33282 42196 33294
rect 42364 33348 42420 33358
rect 41916 33234 41972 33246
rect 41916 33182 41918 33234
rect 41970 33182 41972 33234
rect 41916 32788 41972 33182
rect 42252 33122 42308 33134
rect 42252 33070 42254 33122
rect 42306 33070 42308 33122
rect 42028 32788 42084 32798
rect 41916 32732 42028 32788
rect 42028 32722 42084 32732
rect 41804 29426 41860 31948
rect 42140 32562 42196 32574
rect 42140 32510 42142 32562
rect 42194 32510 42196 32562
rect 42140 31220 42196 32510
rect 42252 31778 42308 33070
rect 42252 31726 42254 31778
rect 42306 31726 42308 31778
rect 42252 31714 42308 31726
rect 42140 31154 42196 31164
rect 42364 30882 42420 33292
rect 42476 32450 42532 34300
rect 42588 33346 42644 38612
rect 42700 36372 42756 36382
rect 42700 35810 42756 36316
rect 42700 35758 42702 35810
rect 42754 35758 42756 35810
rect 42700 35746 42756 35758
rect 42700 34244 42756 34254
rect 42700 34150 42756 34188
rect 42588 33294 42590 33346
rect 42642 33294 42644 33346
rect 42588 33282 42644 33294
rect 42700 33796 42756 33806
rect 42476 32398 42478 32450
rect 42530 32398 42532 32450
rect 42476 32386 42532 32398
rect 42700 31780 42756 33740
rect 42812 31892 42868 40348
rect 43148 40404 43204 41020
rect 43484 41076 43540 42702
rect 43820 42642 43876 42654
rect 43820 42590 43822 42642
rect 43874 42590 43876 42642
rect 43820 42196 43876 42590
rect 43820 42130 43876 42140
rect 45724 42196 45780 42206
rect 45724 42102 45780 42140
rect 43484 41010 43540 41020
rect 43148 40338 43204 40348
rect 45052 40404 45108 40414
rect 45052 40310 45108 40348
rect 43708 37828 43764 37838
rect 43484 37826 43764 37828
rect 43484 37774 43710 37826
rect 43762 37774 43764 37826
rect 43484 37772 43764 37774
rect 43484 37492 43540 37772
rect 43708 37762 43764 37772
rect 44156 37826 44212 37838
rect 44156 37774 44158 37826
rect 44210 37774 44212 37826
rect 43148 37380 43204 37390
rect 43148 37286 43204 37324
rect 42924 37268 42980 37278
rect 43372 37268 43428 37278
rect 42924 37266 43092 37268
rect 42924 37214 42926 37266
rect 42978 37214 43092 37266
rect 42924 37212 43092 37214
rect 42924 37202 42980 37212
rect 43036 36706 43092 37212
rect 43372 37174 43428 37212
rect 43036 36654 43038 36706
rect 43090 36654 43092 36706
rect 43036 36642 43092 36654
rect 43372 36708 43428 36718
rect 43484 36708 43540 37436
rect 44044 37380 44100 37390
rect 44044 37266 44100 37324
rect 44044 37214 44046 37266
rect 44098 37214 44100 37266
rect 44044 37202 44100 37214
rect 44156 37268 44212 37774
rect 44156 37202 44212 37212
rect 43372 36706 43540 36708
rect 43372 36654 43374 36706
rect 43426 36654 43540 36706
rect 43372 36652 43540 36654
rect 43708 37156 43764 37166
rect 43372 36642 43428 36652
rect 43260 36372 43316 36382
rect 43260 35922 43316 36316
rect 43708 36370 43764 37100
rect 46508 37154 46564 37166
rect 46508 37102 46510 37154
rect 46562 37102 46564 37154
rect 43708 36318 43710 36370
rect 43762 36318 43764 36370
rect 43708 36306 43764 36318
rect 44156 36372 44212 36382
rect 44156 36278 44212 36316
rect 44828 36372 44884 36382
rect 43260 35870 43262 35922
rect 43314 35870 43316 35922
rect 43260 35858 43316 35870
rect 44828 36260 44884 36316
rect 46508 36372 46564 37102
rect 46508 36306 46564 36316
rect 44940 36260 44996 36270
rect 44828 36258 44996 36260
rect 44828 36206 44942 36258
rect 44994 36206 44996 36258
rect 44828 36204 44996 36206
rect 43036 34804 43092 34814
rect 43372 34804 43428 34814
rect 42924 34692 42980 34702
rect 42924 33348 42980 34636
rect 43036 33796 43092 34748
rect 43036 33730 43092 33740
rect 43148 34802 43428 34804
rect 43148 34750 43374 34802
rect 43426 34750 43428 34802
rect 43148 34748 43428 34750
rect 43036 33572 43092 33582
rect 43148 33572 43204 34748
rect 43372 34738 43428 34748
rect 43708 34690 43764 34702
rect 43708 34638 43710 34690
rect 43762 34638 43764 34690
rect 43260 34130 43316 34142
rect 43260 34078 43262 34130
rect 43314 34078 43316 34130
rect 43260 33684 43316 34078
rect 43708 34130 43764 34638
rect 44156 34692 44212 34702
rect 44156 34598 44212 34636
rect 43708 34078 43710 34130
rect 43762 34078 43764 34130
rect 43708 34066 43764 34078
rect 43932 34244 43988 34254
rect 43260 33618 43316 33628
rect 43036 33570 43204 33572
rect 43036 33518 43038 33570
rect 43090 33518 43204 33570
rect 43036 33516 43204 33518
rect 43036 33506 43092 33516
rect 43372 33348 43428 33358
rect 42924 33292 43204 33348
rect 43036 32788 43092 32798
rect 43036 32694 43092 32732
rect 43036 31892 43092 31902
rect 42812 31890 43092 31892
rect 42812 31838 43038 31890
rect 43090 31838 43092 31890
rect 42812 31836 43092 31838
rect 43036 31826 43092 31836
rect 43148 31892 43204 33292
rect 43372 33254 43428 33292
rect 43820 33346 43876 33358
rect 43820 33294 43822 33346
rect 43874 33294 43876 33346
rect 43148 31826 43204 31836
rect 42700 31724 42868 31780
rect 42700 31556 42756 31566
rect 42700 31462 42756 31500
rect 42364 30830 42366 30882
rect 42418 30830 42420 30882
rect 41916 30324 41972 30334
rect 41916 30098 41972 30268
rect 41916 30046 41918 30098
rect 41970 30046 41972 30098
rect 41916 30034 41972 30046
rect 42364 30100 42420 30830
rect 42364 30034 42420 30044
rect 42476 29876 42532 29886
rect 41804 29374 41806 29426
rect 41858 29374 41860 29426
rect 41804 29362 41860 29374
rect 41916 29764 41972 29774
rect 41692 28590 41694 28642
rect 41746 28590 41748 28642
rect 41692 28578 41748 28590
rect 41916 28530 41972 29708
rect 41916 28478 41918 28530
rect 41970 28478 41972 28530
rect 41580 27972 41636 27982
rect 41244 27074 41412 27076
rect 41244 27022 41246 27074
rect 41298 27022 41412 27074
rect 41244 27020 41412 27022
rect 41468 27188 41524 27198
rect 41244 26964 41300 27020
rect 41244 26898 41300 26908
rect 41132 26798 41134 26850
rect 41186 26798 41188 26850
rect 41132 26786 41188 26798
rect 40908 26238 40910 26290
rect 40962 26238 40964 26290
rect 40908 26226 40964 26238
rect 41468 26180 41524 27132
rect 41580 27074 41636 27916
rect 41580 27022 41582 27074
rect 41634 27022 41636 27074
rect 41580 27010 41636 27022
rect 41916 27074 41972 28478
rect 42476 28082 42532 29820
rect 42588 29428 42644 29438
rect 42588 29426 42756 29428
rect 42588 29374 42590 29426
rect 42642 29374 42756 29426
rect 42588 29372 42756 29374
rect 42588 29362 42644 29372
rect 42700 28530 42756 29372
rect 42700 28478 42702 28530
rect 42754 28478 42756 28530
rect 42700 28466 42756 28478
rect 42476 28030 42478 28082
rect 42530 28030 42532 28082
rect 42476 28018 42532 28030
rect 42364 27858 42420 27870
rect 42364 27806 42366 27858
rect 42418 27806 42420 27858
rect 42364 27524 42420 27806
rect 42700 27858 42756 27870
rect 42700 27806 42702 27858
rect 42754 27806 42756 27858
rect 42700 27748 42756 27806
rect 42700 27682 42756 27692
rect 42364 27458 42420 27468
rect 42700 27188 42756 27198
rect 42700 27094 42756 27132
rect 41916 27022 41918 27074
rect 41970 27022 41972 27074
rect 41916 27010 41972 27022
rect 42252 27076 42308 27086
rect 42252 26982 42308 27020
rect 42028 26852 42084 26862
rect 42028 26850 42644 26852
rect 42028 26798 42030 26850
rect 42082 26798 42644 26850
rect 42028 26796 42644 26798
rect 42028 26786 42084 26796
rect 41916 26740 41972 26750
rect 41916 26516 41972 26684
rect 41916 26460 42084 26516
rect 42028 26402 42084 26460
rect 42028 26350 42030 26402
rect 42082 26350 42084 26402
rect 42028 26338 42084 26350
rect 42588 26404 42644 26796
rect 42812 26516 42868 31724
rect 43260 31668 43316 31678
rect 43148 31666 43316 31668
rect 43148 31614 43262 31666
rect 43314 31614 43316 31666
rect 43148 31612 43316 31614
rect 43036 30436 43092 30446
rect 43036 30210 43092 30380
rect 43036 30158 43038 30210
rect 43090 30158 43092 30210
rect 43036 30146 43092 30158
rect 43148 30324 43204 31612
rect 43260 31602 43316 31612
rect 43596 31666 43652 31678
rect 43596 31614 43598 31666
rect 43650 31614 43652 31666
rect 43596 30436 43652 31614
rect 43820 30772 43876 33294
rect 43932 33234 43988 34188
rect 43932 33182 43934 33234
rect 43986 33182 43988 33234
rect 43932 33170 43988 33182
rect 43932 31554 43988 31566
rect 43932 31502 43934 31554
rect 43986 31502 43988 31554
rect 43932 30996 43988 31502
rect 44716 30996 44772 31006
rect 43932 30994 44772 30996
rect 43932 30942 44718 30994
rect 44770 30942 44772 30994
rect 43932 30940 44772 30942
rect 44716 30930 44772 30940
rect 43820 30716 44100 30772
rect 43596 30370 43652 30380
rect 43036 28530 43092 28542
rect 43036 28478 43038 28530
rect 43090 28478 43092 28530
rect 43036 28084 43092 28478
rect 43036 28018 43092 28028
rect 43036 27412 43092 27422
rect 43036 27298 43092 27356
rect 43036 27246 43038 27298
rect 43090 27246 43092 27298
rect 43036 27234 43092 27246
rect 43148 26908 43204 30268
rect 43372 30322 43428 30334
rect 43372 30270 43374 30322
rect 43426 30270 43428 30322
rect 43372 29428 43428 30270
rect 44044 30212 44100 30716
rect 44156 30212 44212 30222
rect 44044 30156 44156 30212
rect 44156 30118 44212 30156
rect 43932 30100 43988 30110
rect 43932 30006 43988 30044
rect 43372 29362 43428 29372
rect 44044 29988 44100 29998
rect 44044 28196 44100 29932
rect 43596 27972 43652 27982
rect 43484 27524 43540 27534
rect 42924 26852 43204 26908
rect 43372 27074 43428 27086
rect 43372 27022 43374 27074
rect 43426 27022 43428 27074
rect 43372 26964 43428 27022
rect 43372 26898 43428 26908
rect 42924 26628 42980 26852
rect 42924 26572 43204 26628
rect 42812 26460 42980 26516
rect 42700 26404 42756 26414
rect 42588 26402 42756 26404
rect 42588 26350 42702 26402
rect 42754 26350 42756 26402
rect 42588 26348 42756 26350
rect 42700 26338 42756 26348
rect 41916 26292 41972 26302
rect 41468 26114 41524 26124
rect 41580 26290 41972 26292
rect 41580 26238 41918 26290
rect 41970 26238 41972 26290
rect 41580 26236 41972 26238
rect 40796 25890 40852 25900
rect 40348 24946 40964 24948
rect 40348 24894 40350 24946
rect 40402 24894 40964 24946
rect 40348 24892 40964 24894
rect 40348 24882 40404 24892
rect 40908 24834 40964 24892
rect 40908 24782 40910 24834
rect 40962 24782 40964 24834
rect 40908 24770 40964 24782
rect 41132 24724 41188 24734
rect 41132 24630 41188 24668
rect 41468 24500 41524 24510
rect 41244 24498 41524 24500
rect 41244 24446 41470 24498
rect 41522 24446 41524 24498
rect 41244 24444 41524 24446
rect 41244 24276 41300 24444
rect 41468 24434 41524 24444
rect 40684 24220 41300 24276
rect 39900 23874 39956 23884
rect 40460 23938 40516 23950
rect 40460 23886 40462 23938
rect 40514 23886 40516 23938
rect 40348 23266 40404 23278
rect 40348 23214 40350 23266
rect 40402 23214 40404 23266
rect 40124 23156 40180 23166
rect 40124 23062 40180 23100
rect 39676 23042 39844 23044
rect 39676 22990 39678 23042
rect 39730 22990 39844 23042
rect 39676 22988 39844 22990
rect 39676 22978 39732 22988
rect 39676 22372 39732 22382
rect 39564 22370 39732 22372
rect 39564 22318 39678 22370
rect 39730 22318 39732 22370
rect 39564 22316 39732 22318
rect 39676 22306 39732 22316
rect 39452 22148 39508 22158
rect 39452 22054 39508 22092
rect 39788 22148 39844 22988
rect 40348 22370 40404 23214
rect 40348 22318 40350 22370
rect 40402 22318 40404 22370
rect 40348 22306 40404 22318
rect 39788 22082 39844 22092
rect 40460 22148 40516 23886
rect 40684 23938 40740 24220
rect 41356 24164 41412 24174
rect 41580 24164 41636 26236
rect 41916 26226 41972 26236
rect 42700 25732 42756 25742
rect 41916 25730 42756 25732
rect 41916 25678 42702 25730
rect 42754 25678 42756 25730
rect 41916 25676 42756 25678
rect 41916 25506 41972 25676
rect 42700 25666 42756 25676
rect 41916 25454 41918 25506
rect 41970 25454 41972 25506
rect 41916 25442 41972 25454
rect 41356 24162 41636 24164
rect 41356 24110 41358 24162
rect 41410 24110 41636 24162
rect 41356 24108 41636 24110
rect 42028 25284 42084 25294
rect 42028 24722 42084 25228
rect 42252 25282 42308 25294
rect 42252 25230 42254 25282
rect 42306 25230 42308 25282
rect 42028 24670 42030 24722
rect 42082 24670 42084 24722
rect 41356 24098 41412 24108
rect 40684 23886 40686 23938
rect 40738 23886 40740 23938
rect 40684 23874 40740 23886
rect 41468 23938 41524 23950
rect 41468 23886 41470 23938
rect 41522 23886 41524 23938
rect 41356 23268 41412 23278
rect 41020 23156 41076 23166
rect 41020 23062 41076 23100
rect 41356 23154 41412 23212
rect 41356 23102 41358 23154
rect 41410 23102 41412 23154
rect 41356 23090 41412 23102
rect 40460 22082 40516 22092
rect 41132 22148 41188 22158
rect 39340 21868 39620 21924
rect 39452 21700 39508 21710
rect 39452 21606 39508 21644
rect 39116 21588 39172 21598
rect 39116 20242 39172 21532
rect 39340 21476 39396 21486
rect 39340 21382 39396 21420
rect 39228 21364 39284 21374
rect 39228 21270 39284 21308
rect 39228 20804 39284 20814
rect 39228 20802 39396 20804
rect 39228 20750 39230 20802
rect 39282 20750 39396 20802
rect 39228 20748 39396 20750
rect 39228 20738 39284 20748
rect 39116 20190 39118 20242
rect 39170 20190 39172 20242
rect 39116 20178 39172 20190
rect 39004 20066 39060 20076
rect 38892 20020 38948 20030
rect 38892 18676 38948 19964
rect 39340 19572 39396 20748
rect 39452 19796 39508 19806
rect 39452 19702 39508 19740
rect 39340 19516 39508 19572
rect 38892 16882 38948 18620
rect 39340 19346 39396 19358
rect 39340 19294 39342 19346
rect 39394 19294 39396 19346
rect 39004 18450 39060 18462
rect 39004 18398 39006 18450
rect 39058 18398 39060 18450
rect 39004 18116 39060 18398
rect 39228 18452 39284 18462
rect 39228 18358 39284 18396
rect 39004 18050 39060 18060
rect 39004 17668 39060 17678
rect 39004 17574 39060 17612
rect 39340 17668 39396 19294
rect 39452 18450 39508 19516
rect 39452 18398 39454 18450
rect 39506 18398 39508 18450
rect 39452 18386 39508 18398
rect 39228 17332 39284 17342
rect 39228 16996 39284 17276
rect 39228 16930 39284 16940
rect 38892 16830 38894 16882
rect 38946 16830 38948 16882
rect 38892 16818 38948 16830
rect 39340 16884 39396 17612
rect 39452 16996 39508 17006
rect 39452 16902 39508 16940
rect 39340 16818 39396 16828
rect 39564 16772 39620 21868
rect 40124 21700 40180 21710
rect 40124 21606 40180 21644
rect 41132 21586 41188 22092
rect 41468 21700 41524 23886
rect 42028 23940 42084 24670
rect 41692 23826 41748 23838
rect 41692 23774 41694 23826
rect 41746 23774 41748 23826
rect 41692 23268 41748 23774
rect 41692 23202 41748 23212
rect 41916 23492 41972 23502
rect 41916 23154 41972 23436
rect 41916 23102 41918 23154
rect 41970 23102 41972 23154
rect 41916 23090 41972 23102
rect 42028 22484 42084 23884
rect 42140 24724 42196 24734
rect 42252 24724 42308 25230
rect 42700 24724 42756 24734
rect 42252 24722 42756 24724
rect 42252 24670 42702 24722
rect 42754 24670 42756 24722
rect 42252 24668 42756 24670
rect 42140 23268 42196 24668
rect 42700 24658 42756 24668
rect 42140 23266 42868 23268
rect 42140 23214 42142 23266
rect 42194 23214 42868 23266
rect 42140 23212 42868 23214
rect 42140 23202 42196 23212
rect 41916 22428 42028 22484
rect 41468 21634 41524 21644
rect 41804 21700 41860 21710
rect 41132 21534 41134 21586
rect 41186 21534 41188 21586
rect 41132 21522 41188 21534
rect 40124 21474 40180 21486
rect 40124 21422 40126 21474
rect 40178 21422 40180 21474
rect 39900 21362 39956 21374
rect 39900 21310 39902 21362
rect 39954 21310 39956 21362
rect 39676 21252 39732 21262
rect 39900 21252 39956 21310
rect 39732 21196 39956 21252
rect 39676 21186 39732 21196
rect 40124 20802 40180 21422
rect 40124 20750 40126 20802
rect 40178 20750 40180 20802
rect 40124 20738 40180 20750
rect 41580 20914 41636 20926
rect 41580 20862 41582 20914
rect 41634 20862 41636 20914
rect 39676 20580 39732 20590
rect 39676 20130 39732 20524
rect 39676 20078 39678 20130
rect 39730 20078 39732 20130
rect 39676 20066 39732 20078
rect 40012 20130 40068 20142
rect 40012 20078 40014 20130
rect 40066 20078 40068 20130
rect 40012 18788 40068 20078
rect 40348 19236 40404 19246
rect 40348 19142 40404 19180
rect 41020 19234 41076 19246
rect 41020 19182 41022 19234
rect 41074 19182 41076 19234
rect 41020 19012 41076 19182
rect 41020 18946 41076 18956
rect 39900 18732 40068 18788
rect 39676 18452 39732 18462
rect 39676 18358 39732 18396
rect 39900 17778 39956 18732
rect 41020 18564 41076 18574
rect 41020 18470 41076 18508
rect 40908 18452 40964 18462
rect 40908 18358 40964 18396
rect 40012 18338 40068 18350
rect 40012 18286 40014 18338
rect 40066 18286 40068 18338
rect 40012 18004 40068 18286
rect 40012 17938 40068 17948
rect 40796 18340 40852 18350
rect 39900 17726 39902 17778
rect 39954 17726 39956 17778
rect 39900 17714 39956 17726
rect 40796 17778 40852 18284
rect 41468 18340 41524 18350
rect 40796 17726 40798 17778
rect 40850 17726 40852 17778
rect 40796 17714 40852 17726
rect 41020 18226 41076 18238
rect 41020 18174 41022 18226
rect 41074 18174 41076 18226
rect 40572 17666 40628 17678
rect 40572 17614 40574 17666
rect 40626 17614 40628 17666
rect 40012 17332 40068 17342
rect 40012 17106 40068 17276
rect 40012 17054 40014 17106
rect 40066 17054 40068 17106
rect 40012 17042 40068 17054
rect 40572 16996 40628 17614
rect 41020 17332 41076 18174
rect 41132 17668 41188 17678
rect 41132 17574 41188 17612
rect 41020 17266 41076 17276
rect 41356 17220 41412 17230
rect 40908 17108 40964 17118
rect 40908 17014 40964 17052
rect 41356 17106 41412 17164
rect 41356 17054 41358 17106
rect 41410 17054 41412 17106
rect 41356 17042 41412 17054
rect 40572 16884 40628 16940
rect 41468 16994 41524 18284
rect 41468 16942 41470 16994
rect 41522 16942 41524 16994
rect 41020 16884 41076 16894
rect 41468 16884 41524 16942
rect 40572 16882 41076 16884
rect 40572 16830 41022 16882
rect 41074 16830 41076 16882
rect 40572 16828 41076 16830
rect 39452 16716 39620 16772
rect 39900 16770 39956 16782
rect 39900 16718 39902 16770
rect 39954 16718 39956 16770
rect 39340 16548 39396 16558
rect 38780 16482 38836 16492
rect 39116 16492 39340 16548
rect 38556 16380 38724 16436
rect 38556 15764 38612 16380
rect 38668 16324 38724 16380
rect 38668 16268 38948 16324
rect 38556 15698 38612 15708
rect 38780 15540 38836 15550
rect 38892 15540 38948 16268
rect 39116 16210 39172 16492
rect 39340 16482 39396 16492
rect 39116 16158 39118 16210
rect 39170 16158 39172 16210
rect 39116 16146 39172 16158
rect 39004 15540 39060 15550
rect 38892 15538 39060 15540
rect 38892 15486 39006 15538
rect 39058 15486 39060 15538
rect 38892 15484 39060 15486
rect 38780 15426 38836 15484
rect 39004 15474 39060 15484
rect 38780 15374 38782 15426
rect 38834 15374 38836 15426
rect 38780 15362 38836 15374
rect 38108 15092 38276 15148
rect 38332 15204 38388 15242
rect 38332 15138 38388 15148
rect 38444 15204 38500 15214
rect 38892 15204 38948 15242
rect 38444 15202 38724 15204
rect 38444 15150 38446 15202
rect 38498 15150 38724 15202
rect 38444 15148 38724 15150
rect 39452 15148 39508 16716
rect 39788 16660 39844 16670
rect 39788 16566 39844 16604
rect 39900 16548 39956 16718
rect 39900 16482 39956 16492
rect 38444 15138 38500 15148
rect 38668 15092 38836 15148
rect 38892 15138 38948 15148
rect 37884 14980 37940 14990
rect 37884 14642 37940 14924
rect 37884 14590 37886 14642
rect 37938 14590 37940 14642
rect 37884 14578 37940 14590
rect 37884 13972 37940 13982
rect 37660 13970 37940 13972
rect 37660 13918 37886 13970
rect 37938 13918 37940 13970
rect 37660 13916 37940 13918
rect 37884 13906 37940 13916
rect 37436 12786 37492 12796
rect 37548 13636 37604 13646
rect 37548 12404 37604 13580
rect 37996 13076 38052 13086
rect 37996 12982 38052 13020
rect 37884 12852 37940 12862
rect 38108 12852 38164 15092
rect 38780 14756 38836 15092
rect 39340 15092 39508 15148
rect 39564 15202 39620 15214
rect 39564 15150 39566 15202
rect 39618 15150 39620 15202
rect 38780 14700 39172 14756
rect 38556 14644 38612 14654
rect 38444 14530 38500 14542
rect 38444 14478 38446 14530
rect 38498 14478 38500 14530
rect 38444 13972 38500 14478
rect 38444 13906 38500 13916
rect 38220 13748 38276 13758
rect 38220 13654 38276 13692
rect 37940 12796 38164 12852
rect 37660 12740 37716 12750
rect 37884 12740 37940 12796
rect 37660 12738 37940 12740
rect 37660 12686 37662 12738
rect 37714 12686 37940 12738
rect 37660 12684 37940 12686
rect 37660 12674 37716 12684
rect 37436 12348 37604 12404
rect 37436 12178 37492 12348
rect 37436 12126 37438 12178
rect 37490 12126 37492 12178
rect 37436 12114 37492 12126
rect 37548 12180 37604 12190
rect 37324 11116 37492 11172
rect 37324 10724 37380 10734
rect 37100 10668 37324 10724
rect 37324 10630 37380 10668
rect 37436 10500 37492 11116
rect 37548 10722 37604 12124
rect 37548 10670 37550 10722
rect 37602 10670 37604 10722
rect 37548 10658 37604 10670
rect 37772 11282 37828 11294
rect 37772 11230 37774 11282
rect 37826 11230 37828 11282
rect 37324 10444 37492 10500
rect 37772 10612 37828 11230
rect 37212 10052 37268 10062
rect 36988 9986 37044 9996
rect 37100 9996 37212 10052
rect 37100 9826 37156 9996
rect 37212 9986 37268 9996
rect 37100 9774 37102 9826
rect 37154 9774 37156 9826
rect 37100 9762 37156 9774
rect 37212 9714 37268 9726
rect 37212 9662 37214 9714
rect 37266 9662 37268 9714
rect 37212 9604 37268 9662
rect 37212 9538 37268 9548
rect 36428 8642 36484 8652
rect 37212 9156 37268 9166
rect 37324 9156 37380 10444
rect 37660 9828 37716 9838
rect 37772 9828 37828 10556
rect 37884 10610 37940 12684
rect 37996 12178 38052 12190
rect 37996 12126 37998 12178
rect 38050 12126 38052 12178
rect 37996 11172 38052 12126
rect 38108 12068 38164 12078
rect 38444 12068 38500 12078
rect 38108 12066 38500 12068
rect 38108 12014 38110 12066
rect 38162 12014 38446 12066
rect 38498 12014 38500 12066
rect 38108 12012 38500 12014
rect 38108 12002 38164 12012
rect 38444 12002 38500 12012
rect 38556 11844 38612 14588
rect 39116 14642 39172 14700
rect 39116 14590 39118 14642
rect 39170 14590 39172 14642
rect 39116 14578 39172 14590
rect 38668 13636 38724 13646
rect 38668 13542 38724 13580
rect 38668 12852 38724 12862
rect 38668 12402 38724 12796
rect 38668 12350 38670 12402
rect 38722 12350 38724 12402
rect 38668 12338 38724 12350
rect 39228 12404 39284 12414
rect 39228 12310 39284 12348
rect 38780 12068 38836 12078
rect 38780 11974 38836 12012
rect 38220 11788 38612 11844
rect 38108 11396 38164 11406
rect 38108 11302 38164 11340
rect 38220 11282 38276 11788
rect 38220 11230 38222 11282
rect 38274 11230 38276 11282
rect 38220 11218 38276 11230
rect 39004 11506 39060 11518
rect 39004 11454 39006 11506
rect 39058 11454 39060 11506
rect 37996 11106 38052 11116
rect 38444 11172 38500 11182
rect 38444 11170 38724 11172
rect 38444 11118 38446 11170
rect 38498 11118 38724 11170
rect 38444 11116 38724 11118
rect 38444 11106 38500 11116
rect 38108 10836 38164 10846
rect 38108 10742 38164 10780
rect 38556 10724 38612 10734
rect 37884 10558 37886 10610
rect 37938 10558 37940 10610
rect 37884 10546 37940 10558
rect 38332 10722 38612 10724
rect 38332 10670 38558 10722
rect 38610 10670 38612 10722
rect 38332 10668 38612 10670
rect 37996 10052 38052 10062
rect 37996 9938 38052 9996
rect 37996 9886 37998 9938
rect 38050 9886 38052 9938
rect 37996 9874 38052 9886
rect 37660 9826 37828 9828
rect 37660 9774 37662 9826
rect 37714 9774 37828 9826
rect 37660 9772 37828 9774
rect 37660 9762 37716 9772
rect 37268 9100 37380 9156
rect 37436 9602 37492 9614
rect 37436 9550 37438 9602
rect 37490 9550 37492 9602
rect 37436 9156 37492 9550
rect 37772 9604 37828 9772
rect 37884 9604 37940 9614
rect 37772 9602 37940 9604
rect 37772 9550 37886 9602
rect 37938 9550 37940 9602
rect 37772 9548 37940 9550
rect 37884 9538 37940 9548
rect 38108 9604 38164 9614
rect 38332 9604 38388 10668
rect 38556 10658 38612 10668
rect 38668 10722 38724 11116
rect 38668 10670 38670 10722
rect 38722 10670 38724 10722
rect 38668 10658 38724 10670
rect 38780 10724 38836 10734
rect 38780 10630 38836 10668
rect 38108 9510 38164 9548
rect 38220 9602 38388 9604
rect 38220 9550 38334 9602
rect 38386 9550 38388 9602
rect 38220 9548 38388 9550
rect 37548 9156 37604 9166
rect 37436 9154 37604 9156
rect 37436 9102 37550 9154
rect 37602 9102 37604 9154
rect 37436 9100 37604 9102
rect 37212 8370 37268 9100
rect 37548 9090 37604 9100
rect 37324 8932 37380 8942
rect 37324 8482 37380 8876
rect 38108 8932 38164 8942
rect 38220 8932 38276 9548
rect 38332 9538 38388 9548
rect 38444 10500 38500 10510
rect 38332 9044 38388 9054
rect 38444 9044 38500 10444
rect 39004 9716 39060 11454
rect 39340 10948 39396 15092
rect 39564 14868 39620 15150
rect 41020 15148 41076 16828
rect 41244 16828 41524 16884
rect 41244 16210 41300 16828
rect 41580 16772 41636 20862
rect 41804 19348 41860 21644
rect 41916 19906 41972 22428
rect 42028 22418 42084 22428
rect 42812 22482 42868 23212
rect 42812 22430 42814 22482
rect 42866 22430 42868 22482
rect 42812 22418 42868 22430
rect 42812 21700 42868 21710
rect 42364 21588 42420 21598
rect 42364 21494 42420 21532
rect 42812 21586 42868 21644
rect 42812 21534 42814 21586
rect 42866 21534 42868 21586
rect 42812 21522 42868 21534
rect 42924 21028 42980 26460
rect 43036 26292 43092 26302
rect 43036 26198 43092 26236
rect 43036 25506 43092 25518
rect 43036 25454 43038 25506
rect 43090 25454 43092 25506
rect 43036 24724 43092 25454
rect 43036 24658 43092 24668
rect 41916 19854 41918 19906
rect 41970 19854 41972 19906
rect 41916 19842 41972 19854
rect 42252 20972 42980 21028
rect 43036 21474 43092 21486
rect 43036 21422 43038 21474
rect 43090 21422 43092 21474
rect 41804 19254 41860 19292
rect 41916 18450 41972 18462
rect 41916 18398 41918 18450
rect 41970 18398 41972 18450
rect 41916 18340 41972 18398
rect 41916 18274 41972 18284
rect 41916 18116 41972 18126
rect 41804 18060 41916 18116
rect 41804 17666 41860 18060
rect 41916 18050 41972 18060
rect 41804 17614 41806 17666
rect 41858 17614 41860 17666
rect 41804 17602 41860 17614
rect 41916 17668 41972 17678
rect 41916 17108 41972 17612
rect 41244 16158 41246 16210
rect 41298 16158 41300 16210
rect 41244 16146 41300 16158
rect 41356 16212 41412 16222
rect 41020 15092 41300 15148
rect 39564 14802 39620 14812
rect 41244 14642 41300 15092
rect 41244 14590 41246 14642
rect 41298 14590 41300 14642
rect 41244 14578 41300 14590
rect 40796 13972 40852 13982
rect 40796 12962 40852 13916
rect 41132 13972 41188 13982
rect 41132 13878 41188 13916
rect 40796 12910 40798 12962
rect 40850 12910 40852 12962
rect 40124 12850 40180 12862
rect 40124 12798 40126 12850
rect 40178 12798 40180 12850
rect 40124 12068 40180 12798
rect 40124 12002 40180 12012
rect 39340 10882 39396 10892
rect 39452 11172 39508 11182
rect 39452 10834 39508 11116
rect 39452 10782 39454 10834
rect 39506 10782 39508 10834
rect 39452 10770 39508 10782
rect 39676 10722 39732 10734
rect 39676 10670 39678 10722
rect 39730 10670 39732 10722
rect 39228 10386 39284 10398
rect 39228 10334 39230 10386
rect 39282 10334 39284 10386
rect 39116 9940 39172 9950
rect 39116 9846 39172 9884
rect 39004 9650 39060 9660
rect 38332 9042 38612 9044
rect 38332 8990 38334 9042
rect 38386 8990 38612 9042
rect 38332 8988 38612 8990
rect 38332 8978 38388 8988
rect 38164 8876 38276 8932
rect 38108 8866 38164 8876
rect 37324 8430 37326 8482
rect 37378 8430 37380 8482
rect 37324 8418 37380 8430
rect 38108 8708 38164 8718
rect 37212 8318 37214 8370
rect 37266 8318 37268 8370
rect 35868 7698 36036 7700
rect 35868 7646 35870 7698
rect 35922 7646 36036 7698
rect 35868 7644 36036 7646
rect 35868 7634 35924 7644
rect 35532 6862 35534 6914
rect 35586 6862 35588 6914
rect 35532 6850 35588 6862
rect 34748 6802 34916 6804
rect 34748 6750 34750 6802
rect 34802 6750 34916 6802
rect 34748 6748 34916 6750
rect 34748 6738 34804 6748
rect 35196 6468 35252 6478
rect 35196 6374 35252 6412
rect 35980 6468 36036 7644
rect 36092 8148 36148 8158
rect 36092 6692 36148 8092
rect 36204 8036 36260 8046
rect 37212 8036 37268 8318
rect 37660 8260 37716 8270
rect 37716 8204 37828 8260
rect 37660 8194 37716 8204
rect 36204 8034 36596 8036
rect 36204 7982 36206 8034
rect 36258 7982 36596 8034
rect 36204 7980 36596 7982
rect 36204 7970 36260 7980
rect 36092 6598 36148 6636
rect 36316 6580 36372 6590
rect 36316 6486 36372 6524
rect 33740 6132 33796 6142
rect 33740 6130 34244 6132
rect 33740 6078 33742 6130
rect 33794 6078 34244 6130
rect 33740 6076 34244 6078
rect 33740 6066 33796 6076
rect 34076 5908 34132 5918
rect 34188 5908 34244 6076
rect 34636 5908 34692 5918
rect 34188 5906 34692 5908
rect 34188 5854 34638 5906
rect 34690 5854 34692 5906
rect 34188 5852 34692 5854
rect 34076 5236 34132 5852
rect 34636 5842 34692 5852
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34076 5170 34132 5180
rect 34636 5236 34692 5246
rect 33628 5058 33684 5068
rect 34636 5122 34692 5180
rect 35532 5236 35588 5246
rect 35980 5236 36036 6412
rect 36428 5236 36484 5246
rect 35588 5234 36484 5236
rect 35588 5182 35982 5234
rect 36034 5182 36430 5234
rect 36482 5182 36484 5234
rect 35588 5180 36484 5182
rect 35532 5142 35588 5180
rect 34636 5070 34638 5122
rect 34690 5070 34692 5122
rect 34636 5058 34692 5070
rect 35084 5124 35140 5134
rect 35084 5030 35140 5068
rect 30268 4958 30270 5010
rect 30322 4958 30324 5010
rect 29596 4946 29652 4956
rect 30268 4946 30324 4958
rect 33852 5012 33908 5022
rect 33852 5010 34132 5012
rect 33852 4958 33854 5010
rect 33906 4958 34132 5010
rect 33852 4956 34132 4958
rect 33852 4946 33908 4956
rect 31388 4900 31444 4910
rect 31388 4806 31444 4844
rect 33740 4900 33796 4910
rect 33292 4788 33348 4798
rect 32284 4452 32340 4462
rect 33068 4452 33124 4462
rect 31948 4340 32004 4350
rect 31612 4338 32004 4340
rect 31612 4286 31950 4338
rect 32002 4286 32004 4338
rect 31612 4284 32004 4286
rect 30044 4116 30100 4126
rect 30044 4022 30100 4060
rect 31164 3892 31220 3902
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 29148 3490 29204 3500
rect 30044 3444 30100 3454
rect 30044 800 30100 3388
rect 31164 800 31220 3836
rect 31276 3556 31332 3566
rect 31276 3462 31332 3500
rect 31612 3442 31668 4284
rect 31948 4274 32004 4284
rect 31612 3390 31614 3442
rect 31666 3390 31668 3442
rect 31612 3378 31668 3390
rect 32284 800 32340 4396
rect 32620 4450 33124 4452
rect 32620 4398 33070 4450
rect 33122 4398 33124 4450
rect 32620 4396 33124 4398
rect 32620 3554 32676 4396
rect 33068 4386 33124 4396
rect 33292 4338 33348 4732
rect 33740 4450 33796 4844
rect 34076 4562 34132 4956
rect 34076 4510 34078 4562
rect 34130 4510 34132 4562
rect 34076 4498 34132 4510
rect 33740 4398 33742 4450
rect 33794 4398 33796 4450
rect 33740 4386 33796 4398
rect 34412 4450 34468 4462
rect 34412 4398 34414 4450
rect 34466 4398 34468 4450
rect 33292 4286 33294 4338
rect 33346 4286 33348 4338
rect 33292 4274 33348 4286
rect 32620 3502 32622 3554
rect 32674 3502 32676 3554
rect 32620 3490 32676 3502
rect 33404 4116 33460 4126
rect 33404 800 33460 4060
rect 34412 3892 34468 4398
rect 34860 4452 34916 4462
rect 34860 4358 34916 4396
rect 35868 4450 35924 5180
rect 35980 5170 36036 5180
rect 35868 4398 35870 4450
rect 35922 4398 35924 4450
rect 35868 4386 35924 4398
rect 36428 4338 36484 5180
rect 36428 4286 36430 4338
rect 36482 4286 36484 4338
rect 36428 4274 36484 4286
rect 35308 4116 35364 4154
rect 35756 4116 35812 4126
rect 35308 4050 35364 4060
rect 35532 4114 35812 4116
rect 35532 4062 35758 4114
rect 35810 4062 35812 4114
rect 35532 4060 35812 4062
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34412 3826 34468 3836
rect 35532 3780 35588 4060
rect 35756 4050 35812 4060
rect 35196 3724 35588 3780
rect 34524 3668 34580 3678
rect 33740 3444 33796 3482
rect 33740 3378 33796 3388
rect 34524 800 34580 3612
rect 35196 3554 35252 3724
rect 35196 3502 35198 3554
rect 35250 3502 35252 3554
rect 35196 3490 35252 3502
rect 36428 3556 36484 3566
rect 36540 3556 36596 7980
rect 37212 7970 37268 7980
rect 37548 8148 37604 8158
rect 37212 7812 37268 7822
rect 36652 7700 36708 7710
rect 36652 7606 36708 7644
rect 37100 7362 37156 7374
rect 37100 7310 37102 7362
rect 37154 7310 37156 7362
rect 37100 6580 37156 7310
rect 37212 6690 37268 7756
rect 37548 7474 37604 8092
rect 37548 7422 37550 7474
rect 37602 7422 37604 7474
rect 37548 7410 37604 7422
rect 37212 6638 37214 6690
rect 37266 6638 37268 6690
rect 37212 6626 37268 6638
rect 37548 6692 37604 6702
rect 37772 6692 37828 8204
rect 37884 8036 37940 8046
rect 37884 7942 37940 7980
rect 37884 7700 37940 7710
rect 37884 7474 37940 7644
rect 38108 7698 38164 8652
rect 38556 8370 38612 8988
rect 39228 9042 39284 10334
rect 39676 9492 39732 10670
rect 39788 10612 39844 10622
rect 39788 10518 39844 10556
rect 40796 10500 40852 12910
rect 41132 12964 41188 12974
rect 41356 12964 41412 16156
rect 41468 15652 41524 15662
rect 41468 15148 41524 15596
rect 41580 15540 41636 16716
rect 41692 17106 41972 17108
rect 41692 17054 41918 17106
rect 41970 17054 41972 17106
rect 41692 17052 41972 17054
rect 41692 16212 41748 17052
rect 41916 17042 41972 17052
rect 41692 16118 41748 16156
rect 41580 15484 41748 15540
rect 41692 15314 41748 15484
rect 41692 15262 41694 15314
rect 41746 15262 41748 15314
rect 41468 15092 41636 15148
rect 41132 12962 41412 12964
rect 41132 12910 41134 12962
rect 41186 12910 41412 12962
rect 41132 12908 41412 12910
rect 41132 12740 41188 12908
rect 41020 12068 41076 12078
rect 41132 12068 41188 12684
rect 41020 12066 41188 12068
rect 41020 12014 41022 12066
rect 41074 12014 41188 12066
rect 41020 12012 41188 12014
rect 41020 11396 41076 12012
rect 41020 11330 41076 11340
rect 41132 11282 41188 11294
rect 41132 11230 41134 11282
rect 41186 11230 41188 11282
rect 41132 10836 41188 11230
rect 41132 10770 41188 10780
rect 40796 10434 40852 10444
rect 39676 9426 39732 9436
rect 40796 9716 40852 9726
rect 39452 9268 39508 9278
rect 39452 9174 39508 9212
rect 39228 8990 39230 9042
rect 39282 8990 39284 9042
rect 39228 8978 39284 8990
rect 38780 8932 38836 8942
rect 38780 8838 38836 8876
rect 40796 8932 40852 9660
rect 41244 9714 41300 9726
rect 41244 9662 41246 9714
rect 41298 9662 41300 9714
rect 41244 9268 41300 9662
rect 41244 9202 41300 9212
rect 41580 8932 41636 15092
rect 41692 14306 41748 15262
rect 42252 15148 42308 20972
rect 42924 20802 42980 20814
rect 42924 20750 42926 20802
rect 42978 20750 42980 20802
rect 42476 20356 42532 20366
rect 42364 19796 42420 19806
rect 42364 18338 42420 19740
rect 42476 19124 42532 20300
rect 42588 20244 42644 20254
rect 42588 19346 42644 20188
rect 42588 19294 42590 19346
rect 42642 19294 42644 19346
rect 42588 19282 42644 19294
rect 42924 20018 42980 20750
rect 42924 19966 42926 20018
rect 42978 19966 42980 20018
rect 42812 19236 42868 19246
rect 42700 19234 42868 19236
rect 42700 19182 42814 19234
rect 42866 19182 42868 19234
rect 42700 19180 42868 19182
rect 42476 19068 42644 19124
rect 42364 18286 42366 18338
rect 42418 18286 42420 18338
rect 42364 18274 42420 18286
rect 42364 17332 42420 17342
rect 42364 17106 42420 17276
rect 42364 17054 42366 17106
rect 42418 17054 42420 17106
rect 42364 17042 42420 17054
rect 42476 15314 42532 15326
rect 42476 15262 42478 15314
rect 42530 15262 42532 15314
rect 42252 15092 42420 15148
rect 41692 14254 41694 14306
rect 41746 14254 41748 14306
rect 41692 13972 41748 14254
rect 41692 13906 41748 13916
rect 41916 12964 41972 12974
rect 41916 12962 42308 12964
rect 41916 12910 41918 12962
rect 41970 12910 42308 12962
rect 41916 12908 42308 12910
rect 41916 12898 41972 12908
rect 42252 12402 42308 12908
rect 42252 12350 42254 12402
rect 42306 12350 42308 12402
rect 42252 12338 42308 12350
rect 41916 11396 41972 11406
rect 42364 11396 42420 15092
rect 42476 14418 42532 15262
rect 42476 14366 42478 14418
rect 42530 14366 42532 14418
rect 42476 14354 42532 14366
rect 42588 12404 42644 19068
rect 42700 15988 42756 19180
rect 42812 19170 42868 19180
rect 42924 19236 42980 19966
rect 42924 19170 42980 19180
rect 43036 18676 43092 21422
rect 43148 20916 43204 26572
rect 43484 22708 43540 27468
rect 43596 25506 43652 27916
rect 43596 25454 43598 25506
rect 43650 25454 43652 25506
rect 43596 23492 43652 25454
rect 43820 26964 43876 26974
rect 43820 25394 43876 26908
rect 44044 26962 44100 28140
rect 44492 27970 44548 27982
rect 44492 27918 44494 27970
rect 44546 27918 44548 27970
rect 44156 27188 44212 27198
rect 44156 27074 44212 27132
rect 44156 27022 44158 27074
rect 44210 27022 44212 27074
rect 44156 27010 44212 27022
rect 44044 26910 44046 26962
rect 44098 26910 44100 26962
rect 44044 26898 44100 26910
rect 44492 26908 44548 27918
rect 44716 27860 44772 27870
rect 44716 27766 44772 27804
rect 44492 26852 44660 26908
rect 43820 25342 43822 25394
rect 43874 25342 43876 25394
rect 43820 25330 43876 25342
rect 44268 26292 44324 26302
rect 43652 23436 44212 23492
rect 43596 23398 43652 23436
rect 44156 23266 44212 23436
rect 44156 23214 44158 23266
rect 44210 23214 44212 23266
rect 44156 23202 44212 23214
rect 43596 22932 43652 22942
rect 43596 22930 43764 22932
rect 43596 22878 43598 22930
rect 43650 22878 43764 22930
rect 43596 22876 43764 22878
rect 43596 22866 43652 22876
rect 43484 22652 43652 22708
rect 43260 22484 43316 22494
rect 43260 22390 43316 22428
rect 43484 21588 43540 21598
rect 43484 21026 43540 21532
rect 43596 21362 43652 22652
rect 43708 22370 43764 22876
rect 43708 22318 43710 22370
rect 43762 22318 43764 22370
rect 43708 22306 43764 22318
rect 43932 22930 43988 22942
rect 43932 22878 43934 22930
rect 43986 22878 43988 22930
rect 43596 21310 43598 21362
rect 43650 21310 43652 21362
rect 43596 21298 43652 21310
rect 43484 20974 43486 21026
rect 43538 20974 43540 21026
rect 43484 20962 43540 20974
rect 43148 20850 43204 20860
rect 43596 20916 43652 20926
rect 43596 20804 43652 20860
rect 43484 20748 43652 20804
rect 43820 20802 43876 20814
rect 43820 20750 43822 20802
rect 43874 20750 43876 20802
rect 43484 20244 43540 20748
rect 43148 20020 43204 20030
rect 43148 19458 43204 19964
rect 43148 19406 43150 19458
rect 43202 19406 43204 19458
rect 43148 19394 43204 19406
rect 43484 19346 43540 20188
rect 43820 20242 43876 20750
rect 43820 20190 43822 20242
rect 43874 20190 43876 20242
rect 43820 20178 43876 20190
rect 43484 19294 43486 19346
rect 43538 19294 43540 19346
rect 43484 19282 43540 19294
rect 43036 18610 43092 18620
rect 43596 19236 43652 19246
rect 43596 18674 43652 19180
rect 43708 19234 43764 19246
rect 43708 19182 43710 19234
rect 43762 19182 43764 19234
rect 43708 19124 43764 19182
rect 43932 19124 43988 22878
rect 44044 22260 44100 22270
rect 44044 22166 44100 22204
rect 44268 22148 44324 26236
rect 44268 22082 44324 22092
rect 44492 22484 44548 22494
rect 44492 21586 44548 22428
rect 44492 21534 44494 21586
rect 44546 21534 44548 21586
rect 44492 21522 44548 21534
rect 44044 20916 44100 20926
rect 44044 20822 44100 20860
rect 44156 20130 44212 20142
rect 44156 20078 44158 20130
rect 44210 20078 44212 20130
rect 43708 19068 43988 19124
rect 43596 18622 43598 18674
rect 43650 18622 43652 18674
rect 43596 18610 43652 18622
rect 42812 18562 42868 18574
rect 42812 18510 42814 18562
rect 42866 18510 42868 18562
rect 42812 18116 42868 18510
rect 43036 18452 43092 18462
rect 42812 18050 42868 18060
rect 42924 18450 43092 18452
rect 42924 18398 43038 18450
rect 43090 18398 43092 18450
rect 42924 18396 43092 18398
rect 42812 17108 42868 17118
rect 42924 17108 42980 18396
rect 43036 18386 43092 18396
rect 43820 17780 43876 17790
rect 43820 17108 43876 17724
rect 42812 17106 42980 17108
rect 42812 17054 42814 17106
rect 42866 17054 42980 17106
rect 42812 17052 42980 17054
rect 43260 17052 43876 17108
rect 42812 17042 42868 17052
rect 43148 16660 43204 16670
rect 43148 16566 43204 16604
rect 43260 16322 43316 17052
rect 43820 16994 43876 17052
rect 43820 16942 43822 16994
rect 43874 16942 43876 16994
rect 43820 16930 43876 16942
rect 43596 16884 43652 16894
rect 43596 16772 43652 16828
rect 43596 16716 43764 16772
rect 43260 16270 43262 16322
rect 43314 16270 43316 16322
rect 43260 16258 43316 16270
rect 43708 16098 43764 16716
rect 43708 16046 43710 16098
rect 43762 16046 43764 16098
rect 43708 16034 43764 16046
rect 42700 15922 42756 15932
rect 43820 15988 43876 15998
rect 43820 15894 43876 15932
rect 42924 15874 42980 15886
rect 42924 15822 42926 15874
rect 42978 15822 42980 15874
rect 42924 15148 42980 15822
rect 42812 15092 42980 15148
rect 43932 15148 43988 19068
rect 44044 19124 44100 19134
rect 44044 19010 44100 19068
rect 44044 18958 44046 19010
rect 44098 18958 44100 19010
rect 44044 18946 44100 18958
rect 44044 18338 44100 18350
rect 44044 18286 44046 18338
rect 44098 18286 44100 18338
rect 44044 17892 44100 18286
rect 44156 18340 44212 20078
rect 44156 18274 44212 18284
rect 44268 20018 44324 20030
rect 44268 19966 44270 20018
rect 44322 19966 44324 20018
rect 44100 17836 44212 17892
rect 44044 17826 44100 17836
rect 44156 17556 44212 17836
rect 44268 17780 44324 19966
rect 44604 19794 44660 26852
rect 44716 23268 44772 23278
rect 44716 23174 44772 23212
rect 44604 19742 44606 19794
rect 44658 19742 44660 19794
rect 44604 19730 44660 19742
rect 44716 18450 44772 18462
rect 44716 18398 44718 18450
rect 44770 18398 44772 18450
rect 44716 17892 44772 18398
rect 44716 17826 44772 17836
rect 44268 17686 44324 17724
rect 44156 17500 44324 17556
rect 43932 15092 44212 15148
rect 42812 14530 42868 15092
rect 42812 14478 42814 14530
rect 42866 14478 42868 14530
rect 42812 14466 42868 14478
rect 42588 12338 42644 12348
rect 44156 13076 44212 15092
rect 44268 15092 44324 17500
rect 44828 16996 44884 36204
rect 44940 36194 44996 36204
rect 46508 34802 46564 34814
rect 46508 34750 46510 34802
rect 46562 34750 46564 34802
rect 46172 34692 46228 34702
rect 45948 34690 46228 34692
rect 45948 34638 46174 34690
rect 46226 34638 46228 34690
rect 45948 34636 46228 34638
rect 45276 33572 45332 33582
rect 45276 33346 45332 33516
rect 45276 33294 45278 33346
rect 45330 33294 45332 33346
rect 45276 31778 45332 33294
rect 45948 33346 46004 34636
rect 46172 34626 46228 34636
rect 46508 34356 46564 34750
rect 46620 34356 46676 34366
rect 46508 34354 46676 34356
rect 46508 34302 46622 34354
rect 46674 34302 46676 34354
rect 46508 34300 46676 34302
rect 46620 34290 46676 34300
rect 46172 34244 46228 34254
rect 46172 34150 46228 34188
rect 46956 34244 47012 34254
rect 46956 34130 47012 34188
rect 46956 34078 46958 34130
rect 47010 34078 47012 34130
rect 46956 34066 47012 34078
rect 47180 34242 47236 34254
rect 47180 34190 47182 34242
rect 47234 34190 47236 34242
rect 45948 33294 45950 33346
rect 46002 33294 46004 33346
rect 45948 33282 46004 33294
rect 46284 32676 46340 32686
rect 45276 31726 45278 31778
rect 45330 31726 45332 31778
rect 45276 30994 45332 31726
rect 45948 32674 46340 32676
rect 45948 32622 46286 32674
rect 46338 32622 46340 32674
rect 45948 32620 46340 32622
rect 45948 31778 46004 32620
rect 46284 32610 46340 32620
rect 45948 31726 45950 31778
rect 46002 31726 46004 31778
rect 45948 31714 46004 31726
rect 46620 32562 46676 32574
rect 46620 32510 46622 32562
rect 46674 32510 46676 32562
rect 46620 31218 46676 32510
rect 46620 31166 46622 31218
rect 46674 31166 46676 31218
rect 46620 31154 46676 31166
rect 46956 32452 47012 32462
rect 45276 30942 45278 30994
rect 45330 30942 45332 30994
rect 44940 29988 44996 29998
rect 44940 29650 44996 29932
rect 44940 29598 44942 29650
rect 44994 29598 44996 29650
rect 44940 29586 44996 29598
rect 45276 29426 45332 30942
rect 46956 30994 47012 32396
rect 46956 30942 46958 30994
rect 47010 30942 47012 30994
rect 46956 30930 47012 30942
rect 47180 31106 47236 34190
rect 47516 34242 47572 34254
rect 47516 34190 47518 34242
rect 47570 34190 47572 34242
rect 47516 32452 47572 34190
rect 47516 32386 47572 32396
rect 48300 33122 48356 33134
rect 48300 33070 48302 33122
rect 48354 33070 48356 33122
rect 48300 32452 48356 33070
rect 48300 32386 48356 32396
rect 48300 31554 48356 31566
rect 48300 31502 48302 31554
rect 48354 31502 48356 31554
rect 47180 31054 47182 31106
rect 47234 31054 47236 31106
rect 47180 30322 47236 31054
rect 47516 31444 47572 31454
rect 47516 31108 47572 31388
rect 48300 31444 48356 31502
rect 48300 31218 48356 31388
rect 48300 31166 48302 31218
rect 48354 31166 48356 31218
rect 48300 31154 48356 31166
rect 47516 31106 47684 31108
rect 47516 31054 47518 31106
rect 47570 31054 47684 31106
rect 47516 31052 47684 31054
rect 47516 31042 47572 31052
rect 47180 30270 47182 30322
rect 47234 30270 47236 30322
rect 46060 30210 46116 30222
rect 46060 30158 46062 30210
rect 46114 30158 46116 30210
rect 45612 29988 45668 29998
rect 45612 29894 45668 29932
rect 45836 29986 45892 29998
rect 45836 29934 45838 29986
rect 45890 29934 45892 29986
rect 45276 29374 45278 29426
rect 45330 29374 45332 29426
rect 45276 29362 45332 29374
rect 45836 29426 45892 29934
rect 45836 29374 45838 29426
rect 45890 29374 45892 29426
rect 45836 29362 45892 29374
rect 45948 28868 46004 28878
rect 46060 28868 46116 30158
rect 47180 30212 47236 30270
rect 47180 30146 47236 30156
rect 45948 28866 46116 28868
rect 45948 28814 45950 28866
rect 46002 28814 46116 28866
rect 45948 28812 46116 28814
rect 46732 29988 46788 29998
rect 45948 28802 46004 28812
rect 45500 28644 45556 28654
rect 45500 28550 45556 28588
rect 46284 28644 46340 28654
rect 46284 28550 46340 28588
rect 46732 28644 46788 29932
rect 46732 28578 46788 28588
rect 46844 29428 46900 29438
rect 46844 28530 46900 29372
rect 46844 28478 46846 28530
rect 46898 28478 46900 28530
rect 46844 28466 46900 28478
rect 46956 28644 47012 28654
rect 46956 28420 47012 28588
rect 47068 28644 47124 28654
rect 47516 28644 47572 28654
rect 47068 28642 47572 28644
rect 47068 28590 47070 28642
rect 47122 28590 47518 28642
rect 47570 28590 47572 28642
rect 47068 28588 47572 28590
rect 47068 28578 47124 28588
rect 46956 28364 47236 28420
rect 46396 28196 46452 28206
rect 45500 28084 45556 28094
rect 45500 27990 45556 28028
rect 46060 27972 46116 27982
rect 46060 27878 46116 27916
rect 46396 27970 46452 28140
rect 47180 28084 47236 28364
rect 47180 28082 47348 28084
rect 47180 28030 47182 28082
rect 47234 28030 47348 28082
rect 47180 28028 47348 28030
rect 47180 28018 47236 28028
rect 46396 27918 46398 27970
rect 46450 27918 46452 27970
rect 46396 27906 46452 27918
rect 45836 27636 45892 27646
rect 45276 27634 45892 27636
rect 45276 27582 45838 27634
rect 45890 27582 45892 27634
rect 45276 27580 45892 27582
rect 45276 26964 45332 27580
rect 45836 27570 45892 27580
rect 45836 27300 45892 27310
rect 45164 26290 45220 26302
rect 45164 26238 45166 26290
rect 45218 26238 45220 26290
rect 44940 26180 44996 26190
rect 45164 26180 45220 26238
rect 44940 26178 45220 26180
rect 44940 26126 44942 26178
rect 44994 26126 45220 26178
rect 44940 26124 45220 26126
rect 44940 25284 44996 26124
rect 44940 25218 44996 25228
rect 45164 24948 45220 24958
rect 45276 24948 45332 26908
rect 45388 27188 45444 27198
rect 45388 25620 45444 27132
rect 45612 27076 45668 27086
rect 45612 26908 45668 27020
rect 45612 26852 45780 26908
rect 45388 25526 45444 25564
rect 45164 24946 45332 24948
rect 45164 24894 45166 24946
rect 45218 24894 45332 24946
rect 45164 24892 45332 24894
rect 45164 24882 45220 24892
rect 45612 24610 45668 24622
rect 45612 24558 45614 24610
rect 45666 24558 45668 24610
rect 45164 23154 45220 23166
rect 45164 23102 45166 23154
rect 45218 23102 45220 23154
rect 44940 22484 44996 22494
rect 45164 22484 45220 23102
rect 45388 22484 45444 22494
rect 45612 22484 45668 24558
rect 44996 22482 45668 22484
rect 44996 22430 45390 22482
rect 45442 22430 45668 22482
rect 44996 22428 45668 22430
rect 44940 20916 44996 22428
rect 45388 22418 45444 22428
rect 45164 22260 45220 22270
rect 45164 21586 45220 22204
rect 45164 21534 45166 21586
rect 45218 21534 45220 21586
rect 45164 21522 45220 21534
rect 45500 22148 45556 22158
rect 44940 20914 45220 20916
rect 44940 20862 44942 20914
rect 44994 20862 45220 20914
rect 44940 20860 45220 20862
rect 44940 20850 44996 20860
rect 45164 20802 45220 20860
rect 45164 20750 45166 20802
rect 45218 20750 45220 20802
rect 45164 20738 45220 20750
rect 45388 20020 45444 20030
rect 45276 20018 45444 20020
rect 45276 19966 45390 20018
rect 45442 19966 45444 20018
rect 45276 19964 45444 19966
rect 45276 19908 45332 19964
rect 45388 19954 45444 19964
rect 45164 19852 45332 19908
rect 45052 19348 45108 19358
rect 45164 19348 45220 19852
rect 45500 19458 45556 22092
rect 45724 21028 45780 26852
rect 45836 25730 45892 27244
rect 47180 27074 47236 27086
rect 47180 27022 47182 27074
rect 47234 27022 47236 27074
rect 46396 26964 46452 26974
rect 46844 26964 46900 26974
rect 46396 26962 46900 26964
rect 46396 26910 46398 26962
rect 46450 26910 46846 26962
rect 46898 26910 46900 26962
rect 46396 26908 46900 26910
rect 47180 26908 47236 27022
rect 46396 26898 46452 26908
rect 46844 26898 46900 26908
rect 46060 26852 46116 26862
rect 45948 26850 46116 26852
rect 45948 26798 46062 26850
rect 46114 26798 46116 26850
rect 45948 26796 46116 26798
rect 45948 26290 46004 26796
rect 46060 26786 46116 26796
rect 46956 26852 47236 26908
rect 45948 26238 45950 26290
rect 46002 26238 46004 26290
rect 45948 26226 46004 26238
rect 45836 25678 45838 25730
rect 45890 25678 45892 25730
rect 45836 25666 45892 25678
rect 46508 25620 46564 25630
rect 46172 25506 46228 25518
rect 46172 25454 46174 25506
rect 46226 25454 46228 25506
rect 46172 23940 46228 25454
rect 46172 23874 46228 23884
rect 46508 25394 46564 25564
rect 46508 25342 46510 25394
rect 46562 25342 46564 25394
rect 46396 23716 46452 23726
rect 45948 23714 46452 23716
rect 45948 23662 46398 23714
rect 46450 23662 46452 23714
rect 45948 23660 46452 23662
rect 45948 23154 46004 23660
rect 46396 23650 46452 23660
rect 45948 23102 45950 23154
rect 46002 23102 46004 23154
rect 45948 23090 46004 23102
rect 45500 19406 45502 19458
rect 45554 19406 45556 19458
rect 45500 19394 45556 19406
rect 45612 20972 45780 21028
rect 45948 21700 46004 21710
rect 45108 19292 45220 19348
rect 45276 19346 45332 19358
rect 45276 19294 45278 19346
rect 45330 19294 45332 19346
rect 45052 19234 45108 19292
rect 45052 19182 45054 19234
rect 45106 19182 45108 19234
rect 45052 19170 45108 19182
rect 44940 18562 44996 18574
rect 44940 18510 44942 18562
rect 44994 18510 44996 18562
rect 44940 18452 44996 18510
rect 44940 18386 44996 18396
rect 45164 18450 45220 18462
rect 45164 18398 45166 18450
rect 45218 18398 45220 18450
rect 45052 17780 45108 17790
rect 45052 17686 45108 17724
rect 45164 17220 45220 18398
rect 44604 16940 44884 16996
rect 44940 17164 45220 17220
rect 44604 16660 44660 16940
rect 44716 16772 44772 16782
rect 44940 16772 44996 17164
rect 45276 16884 45332 19294
rect 44772 16716 44996 16772
rect 44716 16678 44772 16716
rect 44604 15876 44660 16604
rect 44940 16100 44996 16716
rect 45052 16828 45332 16884
rect 45052 16436 45108 16828
rect 45164 16658 45220 16670
rect 45164 16606 45166 16658
rect 45218 16606 45220 16658
rect 45164 16548 45220 16606
rect 45500 16658 45556 16670
rect 45500 16606 45502 16658
rect 45554 16606 45556 16658
rect 45164 16492 45444 16548
rect 45052 16380 45332 16436
rect 45164 16100 45220 16110
rect 44940 16098 45220 16100
rect 44940 16046 45166 16098
rect 45218 16046 45220 16098
rect 44940 16044 45220 16046
rect 44604 15810 44660 15820
rect 44828 15988 44884 15998
rect 44828 15538 44884 15932
rect 44828 15486 44830 15538
rect 44882 15486 44884 15538
rect 44828 15474 44884 15486
rect 44268 15026 44324 15036
rect 44940 14754 44996 16044
rect 45164 16034 45220 16044
rect 45052 15876 45108 15886
rect 45052 15782 45108 15820
rect 45276 15148 45332 16380
rect 45388 15428 45444 16492
rect 45500 15988 45556 16606
rect 45500 15922 45556 15932
rect 45500 15428 45556 15438
rect 45388 15426 45556 15428
rect 45388 15374 45502 15426
rect 45554 15374 45556 15426
rect 45388 15372 45556 15374
rect 45500 15362 45556 15372
rect 44940 14702 44942 14754
rect 44994 14702 44996 14754
rect 44940 14642 44996 14702
rect 44940 14590 44942 14642
rect 44994 14590 44996 14642
rect 44940 14578 44996 14590
rect 45164 15092 45332 15148
rect 45164 14196 45220 15092
rect 45388 14754 45444 14766
rect 45388 14702 45390 14754
rect 45442 14702 45444 14754
rect 45388 14642 45444 14702
rect 45388 14590 45390 14642
rect 45442 14590 45444 14642
rect 45388 14578 45444 14590
rect 45164 14140 45332 14196
rect 45164 13972 45220 13982
rect 45164 13878 45220 13916
rect 44268 13076 44324 13086
rect 44156 13074 44324 13076
rect 44156 13022 44270 13074
rect 44322 13022 44324 13074
rect 44156 13020 44324 13022
rect 44156 12290 44212 13020
rect 44268 13010 44324 13020
rect 45164 12962 45220 12974
rect 45164 12910 45166 12962
rect 45218 12910 45220 12962
rect 44940 12740 44996 12750
rect 45164 12740 45220 12910
rect 44996 12684 45220 12740
rect 44940 12646 44996 12684
rect 44156 12238 44158 12290
rect 44210 12238 44212 12290
rect 44156 12226 44212 12238
rect 44828 12404 44884 12414
rect 42588 12180 42644 12190
rect 43260 12180 43316 12190
rect 42588 12178 43316 12180
rect 42588 12126 42590 12178
rect 42642 12126 43262 12178
rect 43314 12126 43316 12178
rect 42588 12124 43316 12126
rect 42588 12114 42644 12124
rect 43260 12114 43316 12124
rect 44380 12178 44436 12190
rect 44380 12126 44382 12178
rect 44434 12126 44436 12178
rect 43596 12068 43652 12078
rect 43596 11974 43652 12012
rect 44380 11844 44436 12126
rect 44380 11778 44436 11788
rect 42364 11340 42532 11396
rect 41916 11172 41972 11340
rect 42364 11172 42420 11182
rect 41916 11170 42420 11172
rect 41916 11118 42366 11170
rect 42418 11118 42420 11170
rect 41916 11116 42420 11118
rect 41916 9716 41972 11116
rect 42364 11106 42420 11116
rect 42140 10610 42196 10622
rect 42140 10558 42142 10610
rect 42194 10558 42196 10610
rect 42140 10500 42196 10558
rect 42140 10434 42196 10444
rect 42028 9826 42084 9838
rect 42028 9774 42030 9826
rect 42082 9774 42084 9826
rect 42028 9716 42084 9774
rect 41972 9660 42084 9716
rect 41916 9650 41972 9660
rect 41580 8876 41748 8932
rect 38556 8318 38558 8370
rect 38610 8318 38612 8370
rect 38556 8306 38612 8318
rect 40572 8148 40628 8158
rect 40572 8054 40628 8092
rect 38108 7646 38110 7698
rect 38162 7646 38164 7698
rect 38108 7634 38164 7646
rect 37884 7422 37886 7474
rect 37938 7422 37940 7474
rect 37884 7410 37940 7422
rect 38780 7588 38836 7598
rect 38780 7474 38836 7532
rect 38780 7422 38782 7474
rect 38834 7422 38836 7474
rect 38780 7410 38836 7422
rect 39340 7476 39396 7486
rect 39340 7474 39508 7476
rect 39340 7422 39342 7474
rect 39394 7422 39508 7474
rect 39340 7420 39508 7422
rect 39340 7410 39396 7420
rect 37996 6692 38052 6702
rect 37772 6690 38276 6692
rect 37772 6638 37998 6690
rect 38050 6638 38276 6690
rect 37772 6636 38276 6638
rect 37548 6598 37604 6636
rect 37996 6626 38052 6636
rect 36988 6132 37044 6142
rect 36988 5234 37044 6076
rect 37100 5794 37156 6524
rect 38220 6130 38276 6636
rect 38220 6078 38222 6130
rect 38274 6078 38276 6130
rect 38220 6066 38276 6078
rect 38556 6578 38612 6590
rect 38556 6526 38558 6578
rect 38610 6526 38612 6578
rect 37436 6020 37492 6030
rect 37100 5742 37102 5794
rect 37154 5742 37156 5794
rect 37100 5348 37156 5742
rect 37100 5282 37156 5292
rect 37212 6018 37492 6020
rect 37212 5966 37438 6018
rect 37490 5966 37492 6018
rect 37212 5964 37492 5966
rect 36988 5182 36990 5234
rect 37042 5182 37044 5234
rect 36988 5170 37044 5182
rect 37100 4898 37156 4910
rect 37100 4846 37102 4898
rect 37154 4846 37156 4898
rect 36988 3668 37044 3678
rect 36988 3574 37044 3612
rect 36484 3500 36596 3556
rect 37100 3556 37156 4846
rect 37212 4338 37268 5964
rect 37436 5954 37492 5964
rect 38556 6020 38612 6526
rect 38668 6468 38724 6478
rect 38668 6130 38724 6412
rect 38668 6078 38670 6130
rect 38722 6078 38724 6130
rect 38668 6066 38724 6078
rect 39004 6466 39060 6478
rect 39004 6414 39006 6466
rect 39058 6414 39060 6466
rect 39004 6244 39060 6414
rect 37660 5906 37716 5918
rect 37660 5854 37662 5906
rect 37714 5854 37716 5906
rect 37660 5346 37716 5854
rect 37660 5294 37662 5346
rect 37714 5294 37716 5346
rect 37660 5282 37716 5294
rect 37996 5348 38052 5358
rect 37996 5254 38052 5292
rect 37212 4286 37214 4338
rect 37266 4286 37268 4338
rect 37212 4274 37268 4286
rect 38444 5124 38500 5134
rect 36428 3462 36484 3500
rect 37100 3490 37156 3500
rect 37884 3668 37940 3678
rect 35420 3332 35476 3342
rect 36764 3332 36820 3342
rect 35420 3330 35700 3332
rect 35420 3278 35422 3330
rect 35474 3278 35700 3330
rect 35420 3276 35700 3278
rect 35420 3266 35476 3276
rect 35644 800 35700 3276
rect 36764 800 36820 3276
rect 37884 800 37940 3612
rect 38444 2996 38500 5068
rect 38556 5122 38612 5964
rect 39004 5908 39060 6188
rect 39004 5852 39284 5908
rect 38556 5070 38558 5122
rect 38610 5070 38612 5122
rect 38556 5058 38612 5070
rect 39116 5682 39172 5694
rect 39116 5630 39118 5682
rect 39170 5630 39172 5682
rect 38780 5012 38836 5022
rect 38780 4918 38836 4956
rect 39116 4452 39172 5630
rect 39228 5122 39284 5852
rect 39228 5070 39230 5122
rect 39282 5070 39284 5122
rect 39228 5058 39284 5070
rect 39452 5906 39508 7420
rect 40236 7474 40292 7486
rect 40236 7422 40238 7474
rect 40290 7422 40292 7474
rect 40236 7252 40292 7422
rect 39788 6468 39844 6478
rect 39788 6374 39844 6412
rect 39676 6020 39732 6030
rect 39676 5926 39732 5964
rect 40236 6018 40292 7196
rect 40348 6692 40404 6702
rect 40796 6692 40852 8876
rect 41580 8260 41636 8270
rect 41244 8258 41636 8260
rect 41244 8206 41582 8258
rect 41634 8206 41636 8258
rect 41244 8204 41636 8206
rect 41244 7698 41300 8204
rect 41580 8194 41636 8204
rect 41692 8260 41748 8876
rect 42476 8260 42532 11340
rect 42924 10612 42980 10622
rect 42924 10610 43204 10612
rect 42924 10558 42926 10610
rect 42978 10558 43204 10610
rect 42924 10556 43204 10558
rect 42924 10546 42980 10556
rect 43148 9714 43204 10556
rect 43484 10388 43540 10398
rect 43484 9826 43540 10332
rect 43484 9774 43486 9826
rect 43538 9774 43540 9826
rect 43484 9762 43540 9774
rect 43148 9662 43150 9714
rect 43202 9662 43204 9714
rect 43148 9650 43204 9662
rect 41692 8194 41748 8204
rect 42364 8204 42532 8260
rect 43820 8372 43876 8382
rect 42364 8148 42420 8204
rect 42364 8082 42420 8092
rect 43148 8148 43204 8158
rect 41244 7646 41246 7698
rect 41298 7646 41300 7698
rect 41244 7634 41300 7646
rect 41356 8034 41412 8046
rect 41356 7982 41358 8034
rect 41410 7982 41412 8034
rect 40348 6690 40852 6692
rect 40348 6638 40350 6690
rect 40402 6638 40798 6690
rect 40850 6638 40852 6690
rect 40348 6636 40852 6638
rect 40348 6626 40404 6636
rect 40236 5966 40238 6018
rect 40290 5966 40292 6018
rect 39452 5854 39454 5906
rect 39506 5854 39508 5906
rect 39452 5012 39508 5854
rect 40236 5908 40292 5966
rect 40236 5852 40516 5908
rect 39452 4564 39508 4956
rect 40236 4900 40292 4910
rect 39900 4898 40292 4900
rect 39900 4846 40238 4898
rect 40290 4846 40292 4898
rect 39900 4844 40292 4846
rect 39564 4564 39620 4574
rect 39452 4562 39620 4564
rect 39452 4510 39566 4562
rect 39618 4510 39620 4562
rect 39452 4508 39620 4510
rect 39564 4498 39620 4508
rect 39116 4386 39172 4396
rect 39788 3556 39844 3566
rect 39788 3462 39844 3500
rect 38892 3332 38948 3342
rect 38892 3238 38948 3276
rect 38444 2930 38500 2940
rect 39004 924 39284 980
rect 39004 800 39060 924
rect 25900 700 26292 756
rect 26656 0 26768 800
rect 27776 0 27888 800
rect 28896 0 29008 800
rect 30016 0 30128 800
rect 31136 0 31248 800
rect 32256 0 32368 800
rect 33376 0 33488 800
rect 34496 0 34608 800
rect 35616 0 35728 800
rect 36736 0 36848 800
rect 37856 0 37968 800
rect 38976 0 39088 800
rect 39228 756 39284 924
rect 39900 756 39956 4844
rect 40236 4834 40292 4844
rect 40460 4564 40516 5852
rect 40796 5796 40852 6636
rect 41356 6690 41412 7982
rect 42476 8034 42532 8046
rect 42476 7982 42478 8034
rect 42530 7982 42532 8034
rect 42364 7586 42420 7598
rect 42364 7534 42366 7586
rect 42418 7534 42420 7586
rect 42028 7474 42084 7486
rect 42028 7422 42030 7474
rect 42082 7422 42084 7474
rect 41580 7252 41636 7262
rect 41580 7158 41636 7196
rect 41356 6638 41358 6690
rect 41410 6638 41412 6690
rect 41356 6626 41412 6638
rect 41468 6020 41524 6030
rect 41244 6018 41524 6020
rect 41244 5966 41470 6018
rect 41522 5966 41524 6018
rect 41244 5964 41524 5966
rect 41020 5796 41076 5806
rect 40796 5794 41076 5796
rect 40796 5742 41022 5794
rect 41074 5742 41076 5794
rect 40796 5740 41076 5742
rect 40908 4564 40964 4574
rect 40460 4562 40964 4564
rect 40460 4510 40910 4562
rect 40962 4510 40964 4562
rect 40460 4508 40964 4510
rect 40908 4498 40964 4508
rect 40012 4452 40068 4462
rect 40012 4358 40068 4396
rect 40348 4452 40404 4462
rect 40348 4358 40404 4396
rect 41020 4340 41076 5740
rect 41020 4274 41076 4284
rect 40796 3668 40852 3678
rect 40796 3574 40852 3612
rect 40124 3332 40180 3342
rect 40124 800 40180 3276
rect 41244 800 41300 5964
rect 41468 5954 41524 5964
rect 42028 6020 42084 7422
rect 42364 6692 42420 7534
rect 42476 7588 42532 7982
rect 42476 7522 42532 7532
rect 43148 7476 43204 8092
rect 43820 7698 43876 8316
rect 43820 7646 43822 7698
rect 43874 7646 43876 7698
rect 43820 7634 43876 7646
rect 44268 7588 44324 7598
rect 44268 7494 44324 7532
rect 43148 7382 43204 7420
rect 43596 7474 43652 7486
rect 43596 7422 43598 7474
rect 43650 7422 43652 7474
rect 42812 7362 42868 7374
rect 42812 7310 42814 7362
rect 42866 7310 42868 7362
rect 42812 6804 42868 7310
rect 43148 6804 43204 6814
rect 42812 6748 43148 6804
rect 42364 6626 42420 6636
rect 42028 5954 42084 5964
rect 42924 6020 42980 6030
rect 42924 5906 42980 5964
rect 43148 6018 43204 6748
rect 43596 6692 43652 7422
rect 43708 6692 43764 6702
rect 43596 6636 43708 6692
rect 43148 5966 43150 6018
rect 43202 5966 43204 6018
rect 43148 5954 43204 5966
rect 43260 6132 43316 6142
rect 42924 5854 42926 5906
rect 42978 5854 42980 5906
rect 42924 5842 42980 5854
rect 42140 5794 42196 5806
rect 42140 5742 42142 5794
rect 42194 5742 42196 5794
rect 42140 5124 42196 5742
rect 43260 5234 43316 6076
rect 43708 5906 43764 6636
rect 44828 6692 44884 12348
rect 45276 12068 45332 14140
rect 45500 13972 45556 13982
rect 45612 13972 45668 20972
rect 45948 20802 46004 21644
rect 45948 20750 45950 20802
rect 46002 20750 46004 20802
rect 45948 20738 46004 20750
rect 46060 20020 46116 20030
rect 46060 19926 46116 19964
rect 46284 20018 46340 20030
rect 46284 19966 46286 20018
rect 46338 19966 46340 20018
rect 46284 19234 46340 19966
rect 46284 19182 46286 19234
rect 46338 19182 46340 19234
rect 45836 19124 45892 19134
rect 45836 19030 45892 19068
rect 46060 18676 46116 18686
rect 45836 18452 45892 18462
rect 45836 18358 45892 18396
rect 45724 17892 45780 17902
rect 45724 17798 45780 17836
rect 46060 17890 46116 18620
rect 46060 17838 46062 17890
rect 46114 17838 46116 17890
rect 45724 16994 45780 17006
rect 45724 16942 45726 16994
rect 45778 16942 45780 16994
rect 45724 16884 45780 16942
rect 45724 16818 45780 16828
rect 46060 16994 46116 17838
rect 46284 17780 46340 19182
rect 46284 17714 46340 17724
rect 46060 16942 46062 16994
rect 46114 16942 46116 16994
rect 46060 16212 46116 16942
rect 46060 16146 46116 16156
rect 45836 16098 45892 16110
rect 45836 16046 45838 16098
rect 45890 16046 45892 16098
rect 45836 15538 45892 16046
rect 45836 15486 45838 15538
rect 45890 15486 45892 15538
rect 45836 15474 45892 15486
rect 45500 13970 45668 13972
rect 45500 13918 45502 13970
rect 45554 13918 45668 13970
rect 45500 13916 45668 13918
rect 46508 13972 46564 25342
rect 46956 25396 47012 26852
rect 46956 25302 47012 25340
rect 47180 23940 47236 23950
rect 46732 23828 46788 23838
rect 46732 23826 46900 23828
rect 46732 23774 46734 23826
rect 46786 23774 46900 23826
rect 46732 23772 46900 23774
rect 46732 23762 46788 23772
rect 46844 22594 46900 23772
rect 46844 22542 46846 22594
rect 46898 22542 46900 22594
rect 46844 22530 46900 22542
rect 47180 22594 47236 23884
rect 47180 22542 47182 22594
rect 47234 22542 47236 22594
rect 47180 19122 47236 22542
rect 47180 19070 47182 19122
rect 47234 19070 47236 19122
rect 47180 19058 47236 19070
rect 47292 23716 47348 28028
rect 46620 18340 46676 18350
rect 46620 17554 46676 18284
rect 46620 17502 46622 17554
rect 46674 17502 46676 17554
rect 46620 17490 46676 17502
rect 46732 17666 46788 17678
rect 46732 17614 46734 17666
rect 46786 17614 46788 17666
rect 46732 16884 46788 17614
rect 46732 16790 46788 16828
rect 47292 17106 47348 23660
rect 47404 26962 47460 28588
rect 47516 28578 47572 28588
rect 47404 26910 47406 26962
rect 47458 26910 47460 26962
rect 47404 22258 47460 26910
rect 47628 26908 47684 31052
rect 48300 29428 48356 29438
rect 48300 29334 48356 29372
rect 47964 28644 48020 28654
rect 47964 28550 48020 28588
rect 48300 27746 48356 27758
rect 48300 27694 48302 27746
rect 48354 27694 48356 27746
rect 47964 26964 48020 26974
rect 48300 26964 48356 27694
rect 47404 22206 47406 22258
rect 47458 22206 47460 22258
rect 47404 19122 47460 22206
rect 47404 19070 47406 19122
rect 47458 19070 47460 19122
rect 47404 19058 47460 19070
rect 47516 26852 47684 26908
rect 47740 26962 48356 26964
rect 47740 26910 47966 26962
rect 48018 26910 48356 26962
rect 47740 26908 48356 26910
rect 47292 17054 47294 17106
rect 47346 17054 47348 17106
rect 47292 16772 47348 17054
rect 46620 15540 46676 15550
rect 46620 15446 46676 15484
rect 47292 15540 47348 16716
rect 47292 15314 47348 15484
rect 47292 15262 47294 15314
rect 47346 15262 47348 15314
rect 47292 15250 47348 15262
rect 46956 15202 47012 15214
rect 46956 15150 46958 15202
rect 47010 15150 47012 15202
rect 46956 14420 47012 15150
rect 47516 15148 47572 26852
rect 47740 26068 47796 26908
rect 47964 26898 48020 26908
rect 48300 26514 48356 26908
rect 48300 26462 48302 26514
rect 48354 26462 48356 26514
rect 48300 26450 48356 26462
rect 47740 26002 47796 26012
rect 48300 25396 48356 25406
rect 48300 23380 48356 25340
rect 47964 23378 48356 23380
rect 47964 23326 48302 23378
rect 48354 23326 48356 23378
rect 47964 23324 48356 23326
rect 47628 23268 47684 23278
rect 47628 21810 47684 23212
rect 47964 22258 48020 23324
rect 48300 23314 48356 23324
rect 48412 23940 48468 23950
rect 47964 22206 47966 22258
rect 48018 22206 48020 22258
rect 47964 22194 48020 22206
rect 47628 21758 47630 21810
rect 47682 21758 47684 21810
rect 47628 21746 47684 21758
rect 47964 21700 48020 21710
rect 47964 21606 48020 21644
rect 48188 21588 48244 21598
rect 48076 21586 48244 21588
rect 48076 21534 48190 21586
rect 48242 21534 48244 21586
rect 48076 21532 48244 21534
rect 48076 19458 48132 21532
rect 48188 21522 48244 21532
rect 48300 20916 48356 20926
rect 48412 20916 48468 23884
rect 48300 20914 48468 20916
rect 48300 20862 48302 20914
rect 48354 20862 48468 20914
rect 48300 20860 48468 20862
rect 48300 20850 48356 20860
rect 48076 19406 48078 19458
rect 48130 19406 48132 19458
rect 48076 19394 48132 19406
rect 47740 19234 47796 19246
rect 47740 19182 47742 19234
rect 47794 19182 47796 19234
rect 47740 18340 47796 19182
rect 47740 18274 47796 18284
rect 48300 18340 48356 18350
rect 48300 18246 48356 18284
rect 47740 16772 47796 16782
rect 47740 16678 47796 16716
rect 48300 16212 48356 16222
rect 48300 16118 48356 16156
rect 47180 15092 48356 15148
rect 47180 14754 47236 15092
rect 47180 14702 47182 14754
rect 47234 14702 47236 14754
rect 47180 14690 47236 14702
rect 47404 14420 47460 14430
rect 46956 14418 47460 14420
rect 46956 14366 47406 14418
rect 47458 14366 47460 14418
rect 46956 14364 47460 14366
rect 46844 14308 46900 14318
rect 45500 13906 45556 13916
rect 46396 13858 46452 13870
rect 46396 13806 46398 13858
rect 46450 13806 46452 13858
rect 45836 13748 45892 13758
rect 45836 13654 45892 13692
rect 45948 12964 46004 12974
rect 45948 12962 46340 12964
rect 45948 12910 45950 12962
rect 46002 12910 46340 12962
rect 45948 12908 46340 12910
rect 45948 12898 46004 12908
rect 46284 12402 46340 12908
rect 46284 12350 46286 12402
rect 46338 12350 46340 12402
rect 46284 12338 46340 12350
rect 45276 10836 45332 12012
rect 46284 11844 46340 11854
rect 45276 10742 45332 10780
rect 45500 11170 45556 11182
rect 45500 11118 45502 11170
rect 45554 11118 45556 11170
rect 44828 6626 44884 6636
rect 44940 10500 44996 10510
rect 44940 9940 44996 10444
rect 45500 10500 45556 11118
rect 45724 10836 45780 10846
rect 45724 10722 45780 10780
rect 45724 10670 45726 10722
rect 45778 10670 45780 10722
rect 45724 10658 45780 10670
rect 45948 10724 46004 10734
rect 45500 10434 45556 10444
rect 44940 9938 45220 9940
rect 44940 9886 44942 9938
rect 44994 9886 45220 9938
rect 44940 9884 45220 9886
rect 44940 8372 44996 9884
rect 45164 9826 45220 9884
rect 45164 9774 45166 9826
rect 45218 9774 45220 9826
rect 45164 9762 45220 9774
rect 45948 9826 46004 10668
rect 46284 10722 46340 11788
rect 46396 11284 46452 13806
rect 46508 13746 46564 13916
rect 46508 13694 46510 13746
rect 46562 13694 46564 13746
rect 46508 13682 46564 13694
rect 46620 14306 46900 14308
rect 46620 14254 46846 14306
rect 46898 14254 46900 14306
rect 46620 14252 46900 14254
rect 46620 12290 46676 14252
rect 46844 14242 46900 14252
rect 46620 12238 46622 12290
rect 46674 12238 46676 12290
rect 46620 12226 46676 12238
rect 46956 11844 47012 14364
rect 47404 14354 47460 14364
rect 47740 14418 47796 14430
rect 47740 14366 47742 14418
rect 47794 14366 47796 14418
rect 46956 11394 47012 11788
rect 47404 13748 47460 13758
rect 47404 11618 47460 13692
rect 47740 13748 47796 14366
rect 48300 13970 48356 15092
rect 48300 13918 48302 13970
rect 48354 13918 48356 13970
rect 48300 13906 48356 13918
rect 47740 13682 47796 13692
rect 48300 13748 48356 13758
rect 48300 13074 48356 13692
rect 48300 13022 48302 13074
rect 48354 13022 48356 13074
rect 48300 13010 48356 13022
rect 47404 11566 47406 11618
rect 47458 11566 47460 11618
rect 47404 11554 47460 11566
rect 46956 11342 46958 11394
rect 47010 11342 47012 11394
rect 46956 11330 47012 11342
rect 46620 11284 46676 11294
rect 46396 11282 46676 11284
rect 46396 11230 46622 11282
rect 46674 11230 46676 11282
rect 46396 11228 46676 11230
rect 46284 10670 46286 10722
rect 46338 10670 46340 10722
rect 46284 10658 46340 10670
rect 46508 10610 46564 11228
rect 46620 11218 46676 11228
rect 47740 11172 47796 11182
rect 47628 11170 47796 11172
rect 47628 11118 47742 11170
rect 47794 11118 47796 11170
rect 47628 11116 47796 11118
rect 47292 10724 47348 10734
rect 47292 10630 47348 10668
rect 47628 10722 47684 11116
rect 47740 11106 47796 11116
rect 47628 10670 47630 10722
rect 47682 10670 47684 10722
rect 47628 10658 47684 10670
rect 46508 10558 46510 10610
rect 46562 10558 46564 10610
rect 46508 9940 46564 10558
rect 46844 10388 46900 10398
rect 46844 10294 46900 10332
rect 46508 9874 46564 9884
rect 48300 9940 48356 9950
rect 48300 9846 48356 9884
rect 45948 9774 45950 9826
rect 46002 9774 46004 9826
rect 45948 9762 46004 9774
rect 45948 9154 46004 9166
rect 45948 9102 45950 9154
rect 46002 9102 46004 9154
rect 44940 8370 45220 8372
rect 44940 8318 44942 8370
rect 44994 8318 45220 8370
rect 44940 8316 45220 8318
rect 43708 5854 43710 5906
rect 43762 5854 43764 5906
rect 43708 5842 43764 5854
rect 44156 6132 44212 6142
rect 44044 5684 44100 5694
rect 43260 5182 43262 5234
rect 43314 5182 43316 5234
rect 43260 5170 43316 5182
rect 43820 5682 44100 5684
rect 43820 5630 44046 5682
rect 44098 5630 44100 5682
rect 43820 5628 44100 5630
rect 42140 5030 42196 5068
rect 43708 5124 43764 5134
rect 43820 5124 43876 5628
rect 44044 5618 44100 5628
rect 43708 5122 43876 5124
rect 43708 5070 43710 5122
rect 43762 5070 43876 5122
rect 43708 5068 43876 5070
rect 43708 5058 43764 5068
rect 42476 4898 42532 4910
rect 42476 4846 42478 4898
rect 42530 4846 42532 4898
rect 42364 3668 42420 3678
rect 42364 800 42420 3612
rect 42476 3556 42532 4846
rect 43932 4898 43988 4910
rect 43932 4846 43934 4898
rect 43986 4846 43988 4898
rect 43260 4452 43316 4462
rect 43260 4338 43316 4396
rect 43260 4286 43262 4338
rect 43314 4286 43316 4338
rect 43260 4274 43316 4286
rect 43820 4340 43876 4350
rect 43820 4246 43876 4284
rect 43932 4116 43988 4846
rect 44156 4338 44212 6076
rect 44940 6132 44996 8316
rect 45164 8258 45220 8316
rect 45164 8206 45166 8258
rect 45218 8206 45220 8258
rect 45164 8194 45220 8206
rect 45388 8260 45444 8270
rect 45052 7588 45108 7598
rect 45052 7474 45108 7532
rect 45052 7422 45054 7474
rect 45106 7422 45108 7474
rect 45052 7410 45108 7422
rect 45052 6692 45108 6702
rect 45052 6598 45108 6636
rect 45388 6132 45444 8204
rect 45948 8258 46004 9102
rect 46284 9044 46340 9054
rect 46284 9042 46564 9044
rect 46284 8990 46286 9042
rect 46338 8990 46564 9042
rect 46284 8988 46564 8990
rect 46284 8978 46340 8988
rect 45948 8206 45950 8258
rect 46002 8206 46004 8258
rect 45948 8194 46004 8206
rect 46508 7698 46564 8988
rect 46508 7646 46510 7698
rect 46562 7646 46564 7698
rect 46508 7634 46564 7646
rect 48300 8034 48356 8046
rect 48300 7982 48302 8034
rect 48354 7982 48356 8034
rect 46956 7588 47012 7598
rect 45500 7476 45556 7486
rect 45500 6690 45556 7420
rect 45500 6638 45502 6690
rect 45554 6638 45556 6690
rect 45500 6626 45556 6638
rect 45948 7474 46004 7486
rect 45948 7422 45950 7474
rect 46002 7422 46004 7474
rect 45948 6580 46004 7422
rect 46844 7250 46900 7262
rect 46844 7198 46846 7250
rect 46898 7198 46900 7250
rect 46844 6804 46900 7198
rect 46956 6914 47012 7532
rect 46956 6862 46958 6914
rect 47010 6862 47012 6914
rect 46956 6850 47012 6862
rect 47180 7586 47236 7598
rect 47180 7534 47182 7586
rect 47234 7534 47236 7586
rect 46844 6692 46900 6748
rect 47180 6692 47236 7534
rect 47628 7588 47684 7598
rect 47628 7494 47684 7532
rect 48300 7588 48356 7982
rect 48300 7522 48356 7532
rect 46844 6636 47124 6692
rect 45948 6514 46004 6524
rect 46172 6580 46228 6590
rect 46620 6580 46676 6590
rect 46172 6578 46676 6580
rect 46172 6526 46174 6578
rect 46226 6526 46622 6578
rect 46674 6526 46676 6578
rect 46172 6524 46676 6526
rect 46172 6514 46228 6524
rect 46620 6514 46676 6524
rect 45836 6466 45892 6478
rect 45836 6414 45838 6466
rect 45890 6414 45892 6466
rect 44996 6076 45220 6132
rect 44940 6038 44996 6076
rect 44828 5236 44884 5246
rect 44828 5234 44996 5236
rect 44828 5182 44830 5234
rect 44882 5182 44996 5234
rect 44828 5180 44996 5182
rect 44828 5170 44884 5180
rect 44828 4340 44884 4350
rect 44156 4286 44158 4338
rect 44210 4286 44212 4338
rect 44156 4274 44212 4286
rect 44268 4338 44884 4340
rect 44268 4286 44830 4338
rect 44882 4286 44884 4338
rect 44268 4284 44884 4286
rect 44268 4116 44324 4284
rect 44828 4274 44884 4284
rect 43932 4060 44324 4116
rect 44604 3668 44660 3678
rect 44604 3574 44660 3612
rect 42476 3490 42532 3500
rect 43596 3556 43652 3566
rect 43596 3462 43652 3500
rect 43484 3444 43540 3454
rect 42700 3332 42756 3342
rect 42700 3238 42756 3276
rect 43484 800 43540 3388
rect 44940 980 44996 5180
rect 45164 5122 45220 6076
rect 45388 6130 45780 6132
rect 45388 6078 45390 6130
rect 45442 6078 45780 6130
rect 45388 6076 45780 6078
rect 45388 6066 45444 6076
rect 45724 5906 45780 6076
rect 45724 5854 45726 5906
rect 45778 5854 45780 5906
rect 45724 5842 45780 5854
rect 45164 5070 45166 5122
rect 45218 5070 45220 5122
rect 45164 5058 45220 5070
rect 45836 5122 45892 6414
rect 45836 5070 45838 5122
rect 45890 5070 45892 5122
rect 45836 5058 45892 5070
rect 46844 5794 46900 5806
rect 46844 5742 46846 5794
rect 46898 5742 46900 5794
rect 46508 3666 46564 3678
rect 46508 3614 46510 3666
rect 46562 3614 46564 3666
rect 46508 3444 46564 3614
rect 46508 3378 46564 3388
rect 44604 924 44996 980
rect 45724 3332 45780 3342
rect 44604 800 44660 924
rect 45724 800 45780 3276
rect 46844 800 46900 5742
rect 47068 4564 47124 6636
rect 47180 6578 47236 6636
rect 48188 7362 48244 7374
rect 48188 7310 48190 7362
rect 48242 7310 48244 7362
rect 48188 6692 48244 7310
rect 48188 6626 48244 6636
rect 47180 6526 47182 6578
rect 47234 6526 47236 6578
rect 47180 6514 47236 6526
rect 47516 6580 47572 6590
rect 47516 6486 47572 6524
rect 48300 6580 48356 6590
rect 48300 5234 48356 6524
rect 48300 5182 48302 5234
rect 48354 5182 48356 5234
rect 48300 5170 48356 5182
rect 47292 4564 47348 4574
rect 47068 4562 47348 4564
rect 47068 4510 47294 4562
rect 47346 4510 47348 4562
rect 47068 4508 47348 4510
rect 47292 4498 47348 4508
rect 48188 3666 48244 3678
rect 48188 3614 48190 3666
rect 48242 3614 48244 3666
rect 48188 3388 48244 3614
rect 47404 3332 47460 3342
rect 47404 3238 47460 3276
rect 47964 3332 48244 3388
rect 47964 800 48020 3332
rect 39228 700 39956 756
rect 40096 0 40208 800
rect 41216 0 41328 800
rect 42336 0 42448 800
rect 43456 0 43568 800
rect 44576 0 44688 800
rect 45696 0 45808 800
rect 46816 0 46928 800
rect 47936 0 48048 800
<< via2 >>
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 14476 49026 14532 49028
rect 14476 48974 14478 49026
rect 14478 48974 14530 49026
rect 14530 48974 14532 49026
rect 14476 48972 14532 48974
rect 16828 48972 16884 49028
rect 15036 48748 15092 48804
rect 16268 48748 16324 48804
rect 16604 48242 16660 48244
rect 16604 48190 16606 48242
rect 16606 48190 16658 48242
rect 16658 48190 16660 48242
rect 16604 48188 16660 48190
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 9996 46844 10052 46900
rect 11004 46844 11060 46900
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 7532 43372 7588 43428
rect 11676 46898 11732 46900
rect 11676 46846 11678 46898
rect 11678 46846 11730 46898
rect 11730 46846 11732 46898
rect 11676 46844 11732 46846
rect 11116 45724 11172 45780
rect 11676 45724 11732 45780
rect 11228 45666 11284 45668
rect 11228 45614 11230 45666
rect 11230 45614 11282 45666
rect 11282 45614 11284 45666
rect 11228 45612 11284 45614
rect 8316 43372 8372 43428
rect 8876 43426 8932 43428
rect 8876 43374 8878 43426
rect 8878 43374 8930 43426
rect 8930 43374 8932 43426
rect 8876 43372 8932 43374
rect 7644 42700 7700 42756
rect 8988 42754 9044 42756
rect 8988 42702 8990 42754
rect 8990 42702 9042 42754
rect 9042 42702 9044 42754
rect 8988 42700 9044 42702
rect 9660 42140 9716 42196
rect 9772 42588 9828 42644
rect 10220 42700 10276 42756
rect 9772 42028 9828 42084
rect 9884 42252 9940 42308
rect 7532 41970 7588 41972
rect 7532 41918 7534 41970
rect 7534 41918 7586 41970
rect 7586 41918 7588 41970
rect 7532 41916 7588 41918
rect 6860 41746 6916 41748
rect 6860 41694 6862 41746
rect 6862 41694 6914 41746
rect 6914 41694 6916 41746
rect 6860 41692 6916 41694
rect 4844 40348 4900 40404
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 2156 38780 2212 38836
rect 5180 38834 5236 38836
rect 5180 38782 5182 38834
rect 5182 38782 5234 38834
rect 5234 38782 5236 38834
rect 5180 38780 5236 38782
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 2604 37938 2660 37940
rect 2604 37886 2606 37938
rect 2606 37886 2658 37938
rect 2658 37886 2660 37938
rect 2604 37884 2660 37886
rect 4172 37100 4228 37156
rect 4284 37436 4340 37492
rect 2828 36370 2884 36372
rect 2828 36318 2830 36370
rect 2830 36318 2882 36370
rect 2882 36318 2884 36370
rect 2828 36316 2884 36318
rect 3836 34860 3892 34916
rect 2716 34130 2772 34132
rect 2716 34078 2718 34130
rect 2718 34078 2770 34130
rect 2770 34078 2772 34130
rect 2716 34076 2772 34078
rect 4172 34130 4228 34132
rect 4172 34078 4174 34130
rect 4174 34078 4226 34130
rect 4226 34078 4228 34130
rect 4172 34076 4228 34078
rect 4956 38108 5012 38164
rect 4844 38050 4900 38052
rect 4844 37998 4846 38050
rect 4846 37998 4898 38050
rect 4898 37998 4900 38050
rect 4844 37996 4900 37998
rect 4732 37436 4788 37492
rect 5740 40348 5796 40404
rect 7084 39842 7140 39844
rect 7084 39790 7086 39842
rect 7086 39790 7138 39842
rect 7138 39790 7140 39842
rect 7084 39788 7140 39790
rect 5740 39676 5796 39732
rect 7644 41692 7700 41748
rect 8988 40514 9044 40516
rect 8988 40462 8990 40514
rect 8990 40462 9042 40514
rect 9042 40462 9044 40514
rect 8988 40460 9044 40462
rect 7644 40348 7700 40404
rect 9212 40124 9268 40180
rect 9324 39676 9380 39732
rect 5740 38780 5796 38836
rect 6636 38220 6692 38276
rect 7420 38220 7476 38276
rect 5516 38108 5572 38164
rect 6076 38162 6132 38164
rect 6076 38110 6078 38162
rect 6078 38110 6130 38162
rect 6130 38110 6132 38162
rect 6076 38108 6132 38110
rect 5292 37996 5348 38052
rect 4732 37154 4788 37156
rect 4732 37102 4734 37154
rect 4734 37102 4786 37154
rect 4786 37102 4788 37154
rect 4732 37100 4788 37102
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4732 34914 4788 34916
rect 4732 34862 4734 34914
rect 4734 34862 4786 34914
rect 4786 34862 4788 34914
rect 4732 34860 4788 34862
rect 5068 34860 5124 34916
rect 6300 37996 6356 38052
rect 5740 37938 5796 37940
rect 5740 37886 5742 37938
rect 5742 37886 5794 37938
rect 5794 37886 5796 37938
rect 5740 37884 5796 37886
rect 5740 36370 5796 36372
rect 5740 36318 5742 36370
rect 5742 36318 5794 36370
rect 5794 36318 5796 36370
rect 5740 36316 5796 36318
rect 5292 34188 5348 34244
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5740 34242 5796 34244
rect 5740 34190 5742 34242
rect 5742 34190 5794 34242
rect 5794 34190 5796 34242
rect 5740 34188 5796 34190
rect 6860 37436 6916 37492
rect 6860 37100 6916 37156
rect 8540 35922 8596 35924
rect 8540 35870 8542 35922
rect 8542 35870 8594 35922
rect 8594 35870 8596 35922
rect 8540 35868 8596 35870
rect 8428 35644 8484 35700
rect 6748 34802 6804 34804
rect 6748 34750 6750 34802
rect 6750 34750 6802 34802
rect 6802 34750 6804 34802
rect 6748 34748 6804 34750
rect 7980 34802 8036 34804
rect 7980 34750 7982 34802
rect 7982 34750 8034 34802
rect 8034 34750 8036 34802
rect 7980 34748 8036 34750
rect 8316 34636 8372 34692
rect 6076 33516 6132 33572
rect 4396 33180 4452 33236
rect 2492 33068 2548 33124
rect 1820 31948 1876 32004
rect 3500 33122 3556 33124
rect 3500 33070 3502 33122
rect 3502 33070 3554 33122
rect 3554 33070 3556 33122
rect 3500 33068 3556 33070
rect 3948 32732 4004 32788
rect 5068 33180 5124 33236
rect 4732 32786 4788 32788
rect 4732 32734 4734 32786
rect 4734 32734 4786 32786
rect 4786 32734 4788 32786
rect 4732 32732 4788 32734
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 2492 31500 2548 31556
rect 3612 31554 3668 31556
rect 3612 31502 3614 31554
rect 3614 31502 3666 31554
rect 3666 31502 3668 31554
rect 3612 31500 3668 31502
rect 6076 31948 6132 32004
rect 5740 31836 5796 31892
rect 3948 30940 4004 30996
rect 5404 31612 5460 31668
rect 4844 31106 4900 31108
rect 4844 31054 4846 31106
rect 4846 31054 4898 31106
rect 4898 31054 4900 31106
rect 4844 31052 4900 31054
rect 5740 31052 5796 31108
rect 5068 30994 5124 30996
rect 5068 30942 5070 30994
rect 5070 30942 5122 30994
rect 5122 30942 5124 30994
rect 5068 30940 5124 30942
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 2828 27858 2884 27860
rect 2828 27806 2830 27858
rect 2830 27806 2882 27858
rect 2882 27806 2884 27858
rect 2828 27804 2884 27806
rect 4060 27858 4116 27860
rect 4060 27806 4062 27858
rect 4062 27806 4114 27858
rect 4114 27806 4116 27858
rect 4060 27804 4116 27806
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 6076 30940 6132 30996
rect 5180 28028 5236 28084
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4172 27074 4228 27076
rect 4172 27022 4174 27074
rect 4174 27022 4226 27074
rect 4226 27022 4228 27074
rect 4172 27020 4228 27022
rect 2604 26962 2660 26964
rect 2604 26910 2606 26962
rect 2606 26910 2658 26962
rect 2658 26910 2660 26962
rect 2604 26908 2660 26910
rect 8092 32620 8148 32676
rect 5628 27074 5684 27076
rect 5628 27022 5630 27074
rect 5630 27022 5682 27074
rect 5682 27022 5684 27074
rect 5628 27020 5684 27022
rect 3836 26962 3892 26964
rect 3836 26910 3838 26962
rect 3838 26910 3890 26962
rect 3890 26910 3892 26962
rect 3836 26908 3892 26910
rect 5180 26290 5236 26292
rect 5180 26238 5182 26290
rect 5182 26238 5234 26290
rect 5234 26238 5236 26290
rect 5180 26236 5236 26238
rect 5740 26236 5796 26292
rect 1932 22428 1988 22484
rect 2044 26012 2100 26068
rect 1708 13692 1764 13748
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4172 23938 4228 23940
rect 4172 23886 4174 23938
rect 4174 23886 4226 23938
rect 4226 23886 4228 23938
rect 4172 23884 4228 23886
rect 2940 23826 2996 23828
rect 2940 23774 2942 23826
rect 2942 23774 2994 23826
rect 2994 23774 2996 23826
rect 2940 23772 2996 23774
rect 3836 23826 3892 23828
rect 3836 23774 3838 23826
rect 3838 23774 3890 23826
rect 3890 23774 3892 23826
rect 3836 23772 3892 23774
rect 5628 24556 5684 24612
rect 4844 23826 4900 23828
rect 4844 23774 4846 23826
rect 4846 23774 4898 23826
rect 4898 23774 4900 23826
rect 4844 23772 4900 23774
rect 4956 23212 5012 23268
rect 4732 23154 4788 23156
rect 4732 23102 4734 23154
rect 4734 23102 4786 23154
rect 4786 23102 4788 23154
rect 4732 23100 4788 23102
rect 5516 23100 5572 23156
rect 2604 22876 2660 22932
rect 5292 22930 5348 22932
rect 5292 22878 5294 22930
rect 5294 22878 5346 22930
rect 5346 22878 5348 22930
rect 5292 22876 5348 22878
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4956 22370 5012 22372
rect 4956 22318 4958 22370
rect 4958 22318 5010 22370
rect 5010 22318 5012 22370
rect 4956 22316 5012 22318
rect 4844 21586 4900 21588
rect 4844 21534 4846 21586
rect 4846 21534 4898 21586
rect 4898 21534 4900 21586
rect 4844 21532 4900 21534
rect 2940 21308 2996 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5852 23266 5908 23268
rect 5852 23214 5854 23266
rect 5854 23214 5906 23266
rect 5906 23214 5908 23266
rect 5852 23212 5908 23214
rect 5740 22316 5796 22372
rect 5740 22146 5796 22148
rect 5740 22094 5742 22146
rect 5742 22094 5794 22146
rect 5794 22094 5796 22146
rect 5740 22092 5796 22094
rect 8428 31836 8484 31892
rect 9660 38834 9716 38836
rect 9660 38782 9662 38834
rect 9662 38782 9714 38834
rect 9714 38782 9716 38834
rect 9660 38780 9716 38782
rect 9996 40178 10052 40180
rect 9996 40126 9998 40178
rect 9998 40126 10050 40178
rect 10050 40126 10052 40178
rect 9996 40124 10052 40126
rect 9660 38162 9716 38164
rect 9660 38110 9662 38162
rect 9662 38110 9714 38162
rect 9714 38110 9716 38162
rect 9660 38108 9716 38110
rect 9436 37938 9492 37940
rect 9436 37886 9438 37938
rect 9438 37886 9490 37938
rect 9490 37886 9492 37938
rect 9436 37884 9492 37886
rect 9100 37266 9156 37268
rect 9100 37214 9102 37266
rect 9102 37214 9154 37266
rect 9154 37214 9156 37266
rect 9100 37212 9156 37214
rect 8876 35868 8932 35924
rect 8876 35532 8932 35588
rect 10108 38556 10164 38612
rect 9996 37324 10052 37380
rect 10892 43708 10948 43764
rect 10892 43372 10948 43428
rect 10444 42140 10500 42196
rect 10332 37938 10388 37940
rect 10332 37886 10334 37938
rect 10334 37886 10386 37938
rect 10386 37886 10388 37938
rect 10332 37884 10388 37886
rect 10108 37212 10164 37268
rect 9884 35420 9940 35476
rect 8428 30322 8484 30324
rect 8428 30270 8430 30322
rect 8430 30270 8482 30322
rect 8482 30270 8484 30322
rect 8428 30268 8484 30270
rect 8316 28700 8372 28756
rect 6636 28588 6692 28644
rect 8204 28642 8260 28644
rect 8204 28590 8206 28642
rect 8206 28590 8258 28642
rect 8258 28590 8260 28642
rect 8204 28588 8260 28590
rect 8652 33516 8708 33572
rect 8988 33516 9044 33572
rect 8876 32620 8932 32676
rect 8764 30098 8820 30100
rect 8764 30046 8766 30098
rect 8766 30046 8818 30098
rect 8818 30046 8820 30098
rect 8764 30044 8820 30046
rect 8652 28476 8708 28532
rect 7868 27468 7924 27524
rect 7644 27132 7700 27188
rect 7756 24050 7812 24052
rect 7756 23998 7758 24050
rect 7758 23998 7810 24050
rect 7810 23998 7812 24050
rect 7756 23996 7812 23998
rect 8988 28588 9044 28644
rect 9660 34690 9716 34692
rect 9660 34638 9662 34690
rect 9662 34638 9714 34690
rect 9714 34638 9716 34690
rect 9660 34636 9716 34638
rect 11116 42754 11172 42756
rect 11116 42702 11118 42754
rect 11118 42702 11170 42754
rect 11170 42702 11172 42754
rect 11116 42700 11172 42702
rect 10668 42588 10724 42644
rect 12684 45724 12740 45780
rect 12908 46898 12964 46900
rect 12908 46846 12910 46898
rect 12910 46846 12962 46898
rect 12962 46846 12964 46898
rect 12908 46844 12964 46846
rect 12012 45612 12068 45668
rect 12012 43538 12068 43540
rect 12012 43486 12014 43538
rect 12014 43486 12066 43538
rect 12066 43486 12068 43538
rect 12012 43484 12068 43486
rect 11564 43426 11620 43428
rect 11564 43374 11566 43426
rect 11566 43374 11618 43426
rect 11618 43374 11620 43426
rect 11564 43372 11620 43374
rect 12348 43708 12404 43764
rect 12236 43650 12292 43652
rect 12236 43598 12238 43650
rect 12238 43598 12290 43650
rect 12290 43598 12292 43650
rect 12236 43596 12292 43598
rect 12124 43372 12180 43428
rect 12012 42754 12068 42756
rect 12012 42702 12014 42754
rect 12014 42702 12066 42754
rect 12066 42702 12068 42754
rect 12012 42700 12068 42702
rect 11452 42252 11508 42308
rect 11564 40908 11620 40964
rect 10556 39788 10612 39844
rect 11564 39788 11620 39844
rect 10556 39340 10612 39396
rect 10780 38834 10836 38836
rect 10780 38782 10782 38834
rect 10782 38782 10834 38834
rect 10834 38782 10836 38834
rect 10780 38780 10836 38782
rect 11788 39228 11844 39284
rect 11676 38668 11732 38724
rect 12460 40962 12516 40964
rect 12460 40910 12462 40962
rect 12462 40910 12514 40962
rect 12514 40910 12516 40962
rect 12460 40908 12516 40910
rect 13132 43596 13188 43652
rect 13580 43484 13636 43540
rect 13916 42754 13972 42756
rect 13916 42702 13918 42754
rect 13918 42702 13970 42754
rect 13970 42702 13972 42754
rect 13916 42700 13972 42702
rect 14364 45778 14420 45780
rect 14364 45726 14366 45778
rect 14366 45726 14418 45778
rect 14418 45726 14420 45778
rect 14364 45724 14420 45726
rect 14812 45778 14868 45780
rect 14812 45726 14814 45778
rect 14814 45726 14866 45778
rect 14866 45726 14868 45778
rect 14812 45724 14868 45726
rect 15708 45724 15764 45780
rect 14028 42252 14084 42308
rect 14700 42252 14756 42308
rect 15596 42028 15652 42084
rect 15484 41916 15540 41972
rect 12796 40572 12852 40628
rect 12236 40460 12292 40516
rect 12124 40402 12180 40404
rect 12124 40350 12126 40402
rect 12126 40350 12178 40402
rect 12178 40350 12180 40402
rect 12124 40348 12180 40350
rect 12908 40348 12964 40404
rect 12460 39506 12516 39508
rect 12460 39454 12462 39506
rect 12462 39454 12514 39506
rect 12514 39454 12516 39506
rect 12460 39452 12516 39454
rect 14588 40684 14644 40740
rect 14476 40572 14532 40628
rect 15036 40572 15092 40628
rect 15372 40962 15428 40964
rect 15372 40910 15374 40962
rect 15374 40910 15426 40962
rect 15426 40910 15428 40962
rect 15372 40908 15428 40910
rect 15484 40626 15540 40628
rect 15484 40574 15486 40626
rect 15486 40574 15538 40626
rect 15538 40574 15540 40626
rect 15484 40572 15540 40574
rect 17612 49026 17668 49028
rect 17612 48974 17614 49026
rect 17614 48974 17666 49026
rect 17666 48974 17668 49026
rect 17612 48972 17668 48974
rect 17276 48188 17332 48244
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 18396 48300 18452 48356
rect 17388 47292 17444 47348
rect 16828 46060 16884 46116
rect 16156 45724 16212 45780
rect 18172 47346 18228 47348
rect 18172 47294 18174 47346
rect 18174 47294 18226 47346
rect 18226 47294 18228 47346
rect 18172 47292 18228 47294
rect 17724 45388 17780 45444
rect 18620 47292 18676 47348
rect 18508 45388 18564 45444
rect 17836 44882 17892 44884
rect 17836 44830 17838 44882
rect 17838 44830 17890 44882
rect 17890 44830 17892 44882
rect 17836 44828 17892 44830
rect 17948 43372 18004 43428
rect 16268 41916 16324 41972
rect 15708 40514 15764 40516
rect 15708 40462 15710 40514
rect 15710 40462 15762 40514
rect 15762 40462 15764 40514
rect 15708 40460 15764 40462
rect 13132 39340 13188 39396
rect 13244 39452 13300 39508
rect 12908 39228 12964 39284
rect 12124 38780 12180 38836
rect 12684 38834 12740 38836
rect 12684 38782 12686 38834
rect 12686 38782 12738 38834
rect 12738 38782 12740 38834
rect 12684 38780 12740 38782
rect 12236 38668 12292 38724
rect 10444 37266 10500 37268
rect 10444 37214 10446 37266
rect 10446 37214 10498 37266
rect 10498 37214 10500 37266
rect 10444 37212 10500 37214
rect 10668 37100 10724 37156
rect 10780 36988 10836 37044
rect 10668 36092 10724 36148
rect 10220 35644 10276 35700
rect 10444 35586 10500 35588
rect 10444 35534 10446 35586
rect 10446 35534 10498 35586
rect 10498 35534 10500 35586
rect 10444 35532 10500 35534
rect 10332 35026 10388 35028
rect 10332 34974 10334 35026
rect 10334 34974 10386 35026
rect 10386 34974 10388 35026
rect 10332 34972 10388 34974
rect 10668 35420 10724 35476
rect 11004 37378 11060 37380
rect 11004 37326 11006 37378
rect 11006 37326 11058 37378
rect 11058 37326 11060 37378
rect 11004 37324 11060 37326
rect 10892 35084 10948 35140
rect 11228 37324 11284 37380
rect 10780 34914 10836 34916
rect 10780 34862 10782 34914
rect 10782 34862 10834 34914
rect 10834 34862 10836 34914
rect 10780 34860 10836 34862
rect 11228 35420 11284 35476
rect 11564 37884 11620 37940
rect 11340 35308 11396 35364
rect 12124 37884 12180 37940
rect 11676 37436 11732 37492
rect 12012 37378 12068 37380
rect 12012 37326 12014 37378
rect 12014 37326 12066 37378
rect 12066 37326 12068 37378
rect 12012 37324 12068 37326
rect 11788 37266 11844 37268
rect 11788 37214 11790 37266
rect 11790 37214 11842 37266
rect 11842 37214 11844 37266
rect 11788 37212 11844 37214
rect 11900 36204 11956 36260
rect 11116 34860 11172 34916
rect 11900 35644 11956 35700
rect 9660 33964 9716 34020
rect 9660 32786 9716 32788
rect 9660 32734 9662 32786
rect 9662 32734 9714 32786
rect 9714 32734 9716 32786
rect 9660 32732 9716 32734
rect 9660 30994 9716 30996
rect 9660 30942 9662 30994
rect 9662 30942 9714 30994
rect 9714 30942 9716 30994
rect 9660 30940 9716 30942
rect 10332 33516 10388 33572
rect 10220 33234 10276 33236
rect 10220 33182 10222 33234
rect 10222 33182 10274 33234
rect 10274 33182 10276 33234
rect 10220 33180 10276 33182
rect 10668 33234 10724 33236
rect 10668 33182 10670 33234
rect 10670 33182 10722 33234
rect 10722 33182 10724 33234
rect 10668 33180 10724 33182
rect 10892 32844 10948 32900
rect 9996 32732 10052 32788
rect 10108 32674 10164 32676
rect 10108 32622 10110 32674
rect 10110 32622 10162 32674
rect 10162 32622 10164 32674
rect 10108 32620 10164 32622
rect 11676 35084 11732 35140
rect 11788 34860 11844 34916
rect 12348 37548 12404 37604
rect 12348 37324 12404 37380
rect 12012 34972 12068 35028
rect 12124 35084 12180 35140
rect 12236 35026 12292 35028
rect 12236 34974 12238 35026
rect 12238 34974 12290 35026
rect 12290 34974 12292 35026
rect 12236 34972 12292 34974
rect 12124 34748 12180 34804
rect 14028 39506 14084 39508
rect 14028 39454 14030 39506
rect 14030 39454 14082 39506
rect 14082 39454 14084 39506
rect 14028 39452 14084 39454
rect 13692 39228 13748 39284
rect 13020 37548 13076 37604
rect 12908 37100 12964 37156
rect 12796 36482 12852 36484
rect 12796 36430 12798 36482
rect 12798 36430 12850 36482
rect 12850 36430 12852 36482
rect 12796 36428 12852 36430
rect 13244 38444 13300 38500
rect 13356 38108 13412 38164
rect 13580 38668 13636 38724
rect 13580 38332 13636 38388
rect 13468 36988 13524 37044
rect 14140 38444 14196 38500
rect 13692 38050 13748 38052
rect 13692 37998 13694 38050
rect 13694 37998 13746 38050
rect 13746 37998 13748 38050
rect 13692 37996 13748 37998
rect 14588 39394 14644 39396
rect 14588 39342 14590 39394
rect 14590 39342 14642 39394
rect 14642 39342 14644 39394
rect 14588 39340 14644 39342
rect 14700 39004 14756 39060
rect 16268 40402 16324 40404
rect 16268 40350 16270 40402
rect 16270 40350 16322 40402
rect 16322 40350 16324 40402
rect 16268 40348 16324 40350
rect 15820 39004 15876 39060
rect 14924 38780 14980 38836
rect 14812 38162 14868 38164
rect 14812 38110 14814 38162
rect 14814 38110 14866 38162
rect 14866 38110 14868 38162
rect 14812 38108 14868 38110
rect 14700 37826 14756 37828
rect 14700 37774 14702 37826
rect 14702 37774 14754 37826
rect 14754 37774 14756 37826
rect 14700 37772 14756 37774
rect 13692 37324 13748 37380
rect 13916 37378 13972 37380
rect 13916 37326 13918 37378
rect 13918 37326 13970 37378
rect 13970 37326 13972 37378
rect 13916 37324 13972 37326
rect 14140 37266 14196 37268
rect 14140 37214 14142 37266
rect 14142 37214 14194 37266
rect 14194 37214 14196 37266
rect 14140 37212 14196 37214
rect 13692 37154 13748 37156
rect 13692 37102 13694 37154
rect 13694 37102 13746 37154
rect 13746 37102 13748 37154
rect 13692 37100 13748 37102
rect 14028 36482 14084 36484
rect 14028 36430 14030 36482
rect 14030 36430 14082 36482
rect 14082 36430 14084 36482
rect 14028 36428 14084 36430
rect 13356 36316 13412 36372
rect 13692 36258 13748 36260
rect 13692 36206 13694 36258
rect 13694 36206 13746 36258
rect 13746 36206 13748 36258
rect 13692 36204 13748 36206
rect 13916 35868 13972 35924
rect 14364 36540 14420 36596
rect 14252 36370 14308 36372
rect 14252 36318 14254 36370
rect 14254 36318 14306 36370
rect 14306 36318 14308 36370
rect 14252 36316 14308 36318
rect 13468 35308 13524 35364
rect 13356 34972 13412 35028
rect 12012 32732 12068 32788
rect 12460 32956 12516 33012
rect 12460 32620 12516 32676
rect 11564 32562 11620 32564
rect 11564 32510 11566 32562
rect 11566 32510 11618 32562
rect 11618 32510 11620 32562
rect 11564 32508 11620 32510
rect 12684 32620 12740 32676
rect 12908 32956 12964 33012
rect 11564 31666 11620 31668
rect 11564 31614 11566 31666
rect 11566 31614 11618 31666
rect 11618 31614 11620 31666
rect 11564 31612 11620 31614
rect 11900 31666 11956 31668
rect 11900 31614 11902 31666
rect 11902 31614 11954 31666
rect 11954 31614 11956 31666
rect 11900 31612 11956 31614
rect 11116 30940 11172 30996
rect 10668 30210 10724 30212
rect 10668 30158 10670 30210
rect 10670 30158 10722 30210
rect 10722 30158 10724 30210
rect 10668 30156 10724 30158
rect 9884 28754 9940 28756
rect 9884 28702 9886 28754
rect 9886 28702 9938 28754
rect 9938 28702 9940 28754
rect 9884 28700 9940 28702
rect 9772 28642 9828 28644
rect 9772 28590 9774 28642
rect 9774 28590 9826 28642
rect 9826 28590 9828 28642
rect 9772 28588 9828 28590
rect 9660 28082 9716 28084
rect 9660 28030 9662 28082
rect 9662 28030 9714 28082
rect 9714 28030 9716 28082
rect 9660 28028 9716 28030
rect 10332 28476 10388 28532
rect 8204 27132 8260 27188
rect 9212 27468 9268 27524
rect 8092 27074 8148 27076
rect 8092 27022 8094 27074
rect 8094 27022 8146 27074
rect 8146 27022 8148 27074
rect 8092 27020 8148 27022
rect 8876 26908 8932 26964
rect 8764 26236 8820 26292
rect 8652 25228 8708 25284
rect 8316 24556 8372 24612
rect 6188 22092 6244 22148
rect 6300 23212 6356 23268
rect 6412 23100 6468 23156
rect 8540 24722 8596 24724
rect 8540 24670 8542 24722
rect 8542 24670 8594 24722
rect 8594 24670 8596 24722
rect 8540 24668 8596 24670
rect 9324 27356 9380 27412
rect 10108 27468 10164 27524
rect 10108 27244 10164 27300
rect 9436 27074 9492 27076
rect 9436 27022 9438 27074
rect 9438 27022 9490 27074
rect 9490 27022 9492 27074
rect 9436 27020 9492 27022
rect 9548 26348 9604 26404
rect 9212 25506 9268 25508
rect 9212 25454 9214 25506
rect 9214 25454 9266 25506
rect 9266 25454 9268 25506
rect 9212 25452 9268 25454
rect 9100 24780 9156 24836
rect 8988 24722 9044 24724
rect 8988 24670 8990 24722
rect 8990 24670 9042 24722
rect 9042 24670 9044 24722
rect 8988 24668 9044 24670
rect 6524 22370 6580 22372
rect 6524 22318 6526 22370
rect 6526 22318 6578 22370
rect 6578 22318 6580 22370
rect 6524 22316 6580 22318
rect 8204 22540 8260 22596
rect 6972 22092 7028 22148
rect 5292 21362 5348 21364
rect 5292 21310 5294 21362
rect 5294 21310 5346 21362
rect 5346 21310 5348 21362
rect 5292 21308 5348 21310
rect 6412 21532 6468 21588
rect 9996 26908 10052 26964
rect 10780 28028 10836 28084
rect 11676 30210 11732 30212
rect 11676 30158 11678 30210
rect 11678 30158 11730 30210
rect 11730 30158 11732 30210
rect 11676 30156 11732 30158
rect 10780 27356 10836 27412
rect 11116 26908 11172 26964
rect 10108 26402 10164 26404
rect 10108 26350 10110 26402
rect 10110 26350 10162 26402
rect 10162 26350 10164 26402
rect 10108 26348 10164 26350
rect 10668 26402 10724 26404
rect 10668 26350 10670 26402
rect 10670 26350 10722 26402
rect 10722 26350 10724 26402
rect 10668 26348 10724 26350
rect 9884 26124 9940 26180
rect 9660 25900 9716 25956
rect 9884 25004 9940 25060
rect 9884 24834 9940 24836
rect 9884 24782 9886 24834
rect 9886 24782 9938 24834
rect 9938 24782 9940 24834
rect 9884 24780 9940 24782
rect 9660 24668 9716 24724
rect 9436 24444 9492 24500
rect 8988 23826 9044 23828
rect 8988 23774 8990 23826
rect 8990 23774 9042 23826
rect 9042 23774 9044 23826
rect 8988 23772 9044 23774
rect 9324 23772 9380 23828
rect 12012 30434 12068 30436
rect 12012 30382 12014 30434
rect 12014 30382 12066 30434
rect 12066 30382 12068 30434
rect 12012 30380 12068 30382
rect 12012 29148 12068 29204
rect 12012 27074 12068 27076
rect 12012 27022 12014 27074
rect 12014 27022 12066 27074
rect 12066 27022 12068 27074
rect 12012 27020 12068 27022
rect 11116 25900 11172 25956
rect 9212 23548 9268 23604
rect 9100 23378 9156 23380
rect 9100 23326 9102 23378
rect 9102 23326 9154 23378
rect 9154 23326 9156 23378
rect 9100 23324 9156 23326
rect 9548 23324 9604 23380
rect 9772 24220 9828 24276
rect 9212 22540 9268 22596
rect 9996 23938 10052 23940
rect 9996 23886 9998 23938
rect 9998 23886 10050 23938
rect 10050 23886 10052 23938
rect 9996 23884 10052 23886
rect 11004 24892 11060 24948
rect 10556 24780 10612 24836
rect 10444 24220 10500 24276
rect 9772 23212 9828 23268
rect 10220 23436 10276 23492
rect 10108 23154 10164 23156
rect 10108 23102 10110 23154
rect 10110 23102 10162 23154
rect 10162 23102 10164 23154
rect 10108 23100 10164 23102
rect 9660 22258 9716 22260
rect 9660 22206 9662 22258
rect 9662 22206 9714 22258
rect 9714 22206 9716 22258
rect 9660 22204 9716 22206
rect 9996 22594 10052 22596
rect 9996 22542 9998 22594
rect 9998 22542 10050 22594
rect 10050 22542 10052 22594
rect 9996 22540 10052 22542
rect 10220 22428 10276 22484
rect 10108 22258 10164 22260
rect 10108 22206 10110 22258
rect 10110 22206 10162 22258
rect 10162 22206 10164 22258
rect 10108 22204 10164 22206
rect 9884 21868 9940 21924
rect 6972 21474 7028 21476
rect 6972 21422 6974 21474
rect 6974 21422 7026 21474
rect 7026 21422 7028 21474
rect 6972 21420 7028 21422
rect 7308 21420 7364 21476
rect 5068 20076 5124 20132
rect 5852 20076 5908 20132
rect 6972 20076 7028 20132
rect 5628 19964 5684 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4396 19404 4452 19460
rect 4172 18956 4228 19012
rect 2604 18450 2660 18452
rect 2604 18398 2606 18450
rect 2606 18398 2658 18450
rect 2658 18398 2660 18450
rect 2604 18396 2660 18398
rect 4060 18450 4116 18452
rect 4060 18398 4062 18450
rect 4062 18398 4114 18450
rect 4114 18398 4116 18450
rect 4060 18396 4116 18398
rect 6524 20018 6580 20020
rect 6524 19966 6526 20018
rect 6526 19966 6578 20018
rect 6578 19966 6580 20018
rect 6524 19964 6580 19966
rect 6972 19404 7028 19460
rect 8988 20914 9044 20916
rect 8988 20862 8990 20914
rect 8990 20862 9042 20914
rect 9042 20862 9044 20914
rect 8988 20860 9044 20862
rect 9772 21586 9828 21588
rect 9772 21534 9774 21586
rect 9774 21534 9826 21586
rect 9826 21534 9828 21586
rect 9772 21532 9828 21534
rect 8204 20748 8260 20804
rect 4732 19010 4788 19012
rect 4732 18958 4734 19010
rect 4734 18958 4786 19010
rect 4786 18958 4788 19010
rect 4732 18956 4788 18958
rect 5180 18956 5236 19012
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4956 17612 5012 17668
rect 2492 17554 2548 17556
rect 2492 17502 2494 17554
rect 2494 17502 2546 17554
rect 2546 17502 2548 17554
rect 2492 17500 2548 17502
rect 3836 17554 3892 17556
rect 3836 17502 3838 17554
rect 3838 17502 3890 17554
rect 3890 17502 3892 17554
rect 3836 17500 3892 17502
rect 4620 17500 4676 17556
rect 4172 16940 4228 16996
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4956 16828 5012 16884
rect 7532 20524 7588 20580
rect 6524 17666 6580 17668
rect 6524 17614 6526 17666
rect 6526 17614 6578 17666
rect 6578 17614 6580 17666
rect 6524 17612 6580 17614
rect 6076 17500 6132 17556
rect 2492 15820 2548 15876
rect 3836 15874 3892 15876
rect 3836 15822 3838 15874
rect 3838 15822 3890 15874
rect 3890 15822 3892 15874
rect 3836 15820 3892 15822
rect 3612 14252 3668 14308
rect 3612 13746 3668 13748
rect 3612 13694 3614 13746
rect 3614 13694 3666 13746
rect 3666 13694 3668 13746
rect 3612 13692 3668 13694
rect 4620 15036 4676 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5740 15036 5796 15092
rect 5068 14252 5124 14308
rect 5180 14700 5236 14756
rect 6748 17554 6804 17556
rect 6748 17502 6750 17554
rect 6750 17502 6802 17554
rect 6802 17502 6804 17554
rect 6748 17500 6804 17502
rect 7084 16940 7140 16996
rect 6076 15036 6132 15092
rect 7084 16044 7140 16100
rect 6076 14754 6132 14756
rect 6076 14702 6078 14754
rect 6078 14702 6130 14754
rect 6130 14702 6132 14754
rect 6076 14700 6132 14702
rect 5964 14252 6020 14308
rect 2604 12850 2660 12852
rect 2604 12798 2606 12850
rect 2606 12798 2658 12850
rect 2658 12798 2660 12850
rect 2604 12796 2660 12798
rect 3836 12850 3892 12852
rect 3836 12798 3838 12850
rect 3838 12798 3890 12850
rect 3890 12798 3892 12850
rect 3836 12796 3892 12798
rect 3612 12348 3668 12404
rect 2492 9714 2548 9716
rect 2492 9662 2494 9714
rect 2494 9662 2546 9714
rect 2546 9662 2548 9714
rect 2492 9660 2548 9662
rect 3500 9714 3556 9716
rect 3500 9662 3502 9714
rect 3502 9662 3554 9714
rect 3554 9662 3556 9714
rect 3500 9660 3556 9662
rect 1708 7644 1764 7700
rect 2492 8764 2548 8820
rect 3388 8818 3444 8820
rect 3388 8766 3390 8818
rect 3390 8766 3442 8818
rect 3442 8766 3444 8818
rect 3388 8764 3444 8766
rect 4172 12348 4228 12404
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4956 13356 5012 13412
rect 5740 13356 5796 13412
rect 4956 12962 5012 12964
rect 4956 12910 4958 12962
rect 4958 12910 5010 12962
rect 5010 12910 5012 12962
rect 4956 12908 5012 12910
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5292 12402 5348 12404
rect 5292 12350 5294 12402
rect 5294 12350 5346 12402
rect 5346 12350 5348 12402
rect 5292 12348 5348 12350
rect 4956 11170 5012 11172
rect 4956 11118 4958 11170
rect 4958 11118 5010 11170
rect 5010 11118 5012 11170
rect 4956 11116 5012 11118
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4396 9154 4452 9156
rect 4396 9102 4398 9154
rect 4398 9102 4450 9154
rect 4450 9102 4452 9154
rect 4396 9100 4452 9102
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4284 7698 4340 7700
rect 4284 7646 4286 7698
rect 4286 7646 4338 7698
rect 4338 7646 4340 7698
rect 4284 7644 4340 7646
rect 1932 5068 1988 5124
rect 2492 6412 2548 6468
rect 2716 4956 2772 5012
rect 3052 5628 3108 5684
rect 3612 6466 3668 6468
rect 3612 6414 3614 6466
rect 3614 6414 3666 6466
rect 3666 6414 3668 6466
rect 3612 6412 3668 6414
rect 4732 7362 4788 7364
rect 4732 7310 4734 7362
rect 4734 7310 4786 7362
rect 4786 7310 4788 7362
rect 4732 7308 4788 7310
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 6300 13804 6356 13860
rect 6972 14252 7028 14308
rect 6860 13692 6916 13748
rect 6748 13356 6804 13412
rect 6188 12908 6244 12964
rect 6412 9714 6468 9716
rect 6412 9662 6414 9714
rect 6414 9662 6466 9714
rect 6466 9662 6468 9714
rect 6412 9660 6468 9662
rect 5180 7308 5236 7364
rect 7420 14812 7476 14868
rect 7308 12348 7364 12404
rect 7084 9100 7140 9156
rect 6636 9042 6692 9044
rect 6636 8990 6638 9042
rect 6638 8990 6690 9042
rect 6690 8990 6692 9042
rect 6636 8988 6692 8990
rect 7420 9042 7476 9044
rect 7420 8990 7422 9042
rect 7422 8990 7474 9042
rect 7474 8990 7476 9042
rect 7420 8988 7476 8990
rect 7420 7756 7476 7812
rect 6076 7308 6132 7364
rect 3724 5628 3780 5684
rect 3724 5292 3780 5348
rect 4732 6130 4788 6132
rect 4732 6078 4734 6130
rect 4734 6078 4786 6130
rect 4786 6078 4788 6130
rect 4732 6076 4788 6078
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4732 5292 4788 5348
rect 3500 5234 3556 5236
rect 3500 5182 3502 5234
rect 3502 5182 3554 5234
rect 3554 5182 3556 5234
rect 3500 5180 3556 5182
rect 3836 5122 3892 5124
rect 3836 5070 3838 5122
rect 3838 5070 3890 5122
rect 3890 5070 3892 5122
rect 3836 5068 3892 5070
rect 5180 6130 5236 6132
rect 5180 6078 5182 6130
rect 5182 6078 5234 6130
rect 5234 6078 5236 6130
rect 5180 6076 5236 6078
rect 5740 4562 5796 4564
rect 5740 4510 5742 4562
rect 5742 4510 5794 4562
rect 5794 4510 5796 4562
rect 5740 4508 5796 4510
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 7196 7362 7252 7364
rect 7196 7310 7198 7362
rect 7198 7310 7250 7362
rect 7250 7310 7252 7362
rect 7196 7308 7252 7310
rect 6748 6578 6804 6580
rect 6748 6526 6750 6578
rect 6750 6526 6802 6578
rect 6802 6526 6804 6578
rect 6748 6524 6804 6526
rect 5516 3836 5572 3892
rect 3276 3724 3332 3780
rect 3724 3724 3780 3780
rect 3164 3612 3220 3668
rect 3388 3500 3444 3556
rect 5628 3724 5684 3780
rect 4284 3612 4340 3668
rect 4060 3442 4116 3444
rect 4060 3390 4062 3442
rect 4062 3390 4114 3442
rect 4114 3390 4116 3442
rect 4060 3388 4116 3390
rect 4396 3276 4452 3332
rect 5964 3554 6020 3556
rect 5964 3502 5966 3554
rect 5966 3502 6018 3554
rect 6018 3502 6020 3554
rect 5964 3500 6020 3502
rect 6188 3442 6244 3444
rect 6188 3390 6190 3442
rect 6190 3390 6242 3442
rect 6242 3390 6244 3442
rect 6188 3388 6244 3390
rect 7084 6412 7140 6468
rect 8540 20636 8596 20692
rect 7868 17388 7924 17444
rect 7756 15036 7812 15092
rect 7644 14476 7700 14532
rect 8428 20578 8484 20580
rect 8428 20526 8430 20578
rect 8430 20526 8482 20578
rect 8482 20526 8484 20578
rect 8428 20524 8484 20526
rect 8428 19346 8484 19348
rect 8428 19294 8430 19346
rect 8430 19294 8482 19346
rect 8482 19294 8484 19346
rect 8428 19292 8484 19294
rect 9660 20690 9716 20692
rect 9660 20638 9662 20690
rect 9662 20638 9714 20690
rect 9714 20638 9716 20690
rect 9660 20636 9716 20638
rect 10668 23436 10724 23492
rect 10892 23212 10948 23268
rect 10332 21698 10388 21700
rect 10332 21646 10334 21698
rect 10334 21646 10386 21698
rect 10386 21646 10388 21698
rect 10332 21644 10388 21646
rect 9996 20860 10052 20916
rect 10556 20524 10612 20580
rect 8988 20130 9044 20132
rect 8988 20078 8990 20130
rect 8990 20078 9042 20130
rect 9042 20078 9044 20130
rect 8988 20076 9044 20078
rect 9884 19292 9940 19348
rect 9212 19010 9268 19012
rect 9212 18958 9214 19010
rect 9214 18958 9266 19010
rect 9266 18958 9268 19010
rect 9212 18956 9268 18958
rect 8876 18844 8932 18900
rect 8764 17666 8820 17668
rect 8764 17614 8766 17666
rect 8766 17614 8818 17666
rect 8818 17614 8820 17666
rect 8764 17612 8820 17614
rect 9324 18396 9380 18452
rect 9660 18284 9716 18340
rect 8988 16994 9044 16996
rect 8988 16942 8990 16994
rect 8990 16942 9042 16994
rect 9042 16942 9044 16994
rect 8988 16940 9044 16942
rect 9772 18060 9828 18116
rect 9996 18956 10052 19012
rect 9884 17666 9940 17668
rect 9884 17614 9886 17666
rect 9886 17614 9938 17666
rect 9938 17614 9940 17666
rect 9884 17612 9940 17614
rect 10444 20018 10500 20020
rect 10444 19966 10446 20018
rect 10446 19966 10498 20018
rect 10498 19966 10500 20018
rect 10444 19964 10500 19966
rect 10556 19346 10612 19348
rect 10556 19294 10558 19346
rect 10558 19294 10610 19346
rect 10610 19294 10612 19346
rect 10556 19292 10612 19294
rect 10108 18284 10164 18340
rect 11340 24892 11396 24948
rect 11564 25394 11620 25396
rect 11564 25342 11566 25394
rect 11566 25342 11618 25394
rect 11618 25342 11620 25394
rect 11564 25340 11620 25342
rect 11340 24722 11396 24724
rect 11340 24670 11342 24722
rect 11342 24670 11394 24722
rect 11394 24670 11396 24722
rect 11340 24668 11396 24670
rect 11228 23884 11284 23940
rect 12012 25618 12068 25620
rect 12012 25566 12014 25618
rect 12014 25566 12066 25618
rect 12066 25566 12068 25618
rect 12012 25564 12068 25566
rect 13804 35084 13860 35140
rect 14140 34972 14196 35028
rect 13468 32844 13524 32900
rect 13132 32620 13188 32676
rect 13468 32562 13524 32564
rect 13468 32510 13470 32562
rect 13470 32510 13522 32562
rect 13522 32510 13524 32562
rect 13468 32508 13524 32510
rect 13356 32450 13412 32452
rect 13356 32398 13358 32450
rect 13358 32398 13410 32450
rect 13410 32398 13412 32450
rect 13356 32396 13412 32398
rect 14588 35084 14644 35140
rect 15036 37378 15092 37380
rect 15036 37326 15038 37378
rect 15038 37326 15090 37378
rect 15090 37326 15092 37378
rect 15036 37324 15092 37326
rect 16268 37938 16324 37940
rect 16268 37886 16270 37938
rect 16270 37886 16322 37938
rect 16322 37886 16324 37938
rect 16268 37884 16324 37886
rect 16156 37772 16212 37828
rect 15484 37490 15540 37492
rect 15484 37438 15486 37490
rect 15486 37438 15538 37490
rect 15538 37438 15540 37490
rect 15484 37436 15540 37438
rect 15372 37212 15428 37268
rect 15148 36540 15204 36596
rect 14700 36204 14756 36260
rect 17052 40908 17108 40964
rect 16940 39618 16996 39620
rect 16940 39566 16942 39618
rect 16942 39566 16994 39618
rect 16994 39566 16996 39618
rect 16940 39564 16996 39566
rect 17612 40514 17668 40516
rect 17612 40462 17614 40514
rect 17614 40462 17666 40514
rect 17666 40462 17668 40514
rect 17612 40460 17668 40462
rect 17500 40402 17556 40404
rect 17500 40350 17502 40402
rect 17502 40350 17554 40402
rect 17554 40350 17556 40402
rect 17500 40348 17556 40350
rect 15708 37042 15764 37044
rect 15708 36990 15710 37042
rect 15710 36990 15762 37042
rect 15762 36990 15764 37042
rect 15708 36988 15764 36990
rect 15372 36540 15428 36596
rect 15260 35756 15316 35812
rect 15820 35922 15876 35924
rect 15820 35870 15822 35922
rect 15822 35870 15874 35922
rect 15874 35870 15876 35922
rect 15820 35868 15876 35870
rect 15596 35532 15652 35588
rect 14476 34412 14532 34468
rect 14028 33180 14084 33236
rect 15036 34300 15092 34356
rect 14476 33404 14532 33460
rect 14364 32844 14420 32900
rect 15372 34690 15428 34692
rect 15372 34638 15374 34690
rect 15374 34638 15426 34690
rect 15426 34638 15428 34690
rect 15372 34636 15428 34638
rect 15372 34412 15428 34468
rect 15372 34188 15428 34244
rect 15596 33458 15652 33460
rect 15596 33406 15598 33458
rect 15598 33406 15650 33458
rect 15650 33406 15652 33458
rect 15596 33404 15652 33406
rect 16156 36204 16212 36260
rect 16380 36204 16436 36260
rect 16492 36988 16548 37044
rect 15820 33346 15876 33348
rect 15820 33294 15822 33346
rect 15822 33294 15874 33346
rect 15874 33294 15876 33346
rect 15820 33292 15876 33294
rect 17612 38946 17668 38948
rect 17612 38894 17614 38946
rect 17614 38894 17666 38946
rect 17666 38894 17668 38946
rect 17612 38892 17668 38894
rect 17388 38834 17444 38836
rect 17388 38782 17390 38834
rect 17390 38782 17442 38834
rect 17442 38782 17444 38834
rect 17388 38780 17444 38782
rect 16940 36876 16996 36932
rect 18396 42754 18452 42756
rect 18396 42702 18398 42754
rect 18398 42702 18450 42754
rect 18450 42702 18452 42754
rect 18396 42700 18452 42702
rect 17948 39004 18004 39060
rect 16940 34972 16996 35028
rect 12684 30940 12740 30996
rect 13580 31612 13636 31668
rect 12572 30882 12628 30884
rect 12572 30830 12574 30882
rect 12574 30830 12626 30882
rect 12626 30830 12628 30882
rect 12572 30828 12628 30830
rect 12572 30268 12628 30324
rect 12236 30098 12292 30100
rect 12236 30046 12238 30098
rect 12238 30046 12290 30098
rect 12290 30046 12292 30098
rect 12236 30044 12292 30046
rect 12348 27244 12404 27300
rect 12572 27244 12628 27300
rect 12572 27020 12628 27076
rect 12684 26962 12740 26964
rect 12684 26910 12686 26962
rect 12686 26910 12738 26962
rect 12738 26910 12740 26962
rect 12684 26908 12740 26910
rect 12348 26236 12404 26292
rect 11900 24892 11956 24948
rect 12124 24162 12180 24164
rect 12124 24110 12126 24162
rect 12126 24110 12178 24162
rect 12178 24110 12180 24162
rect 12124 24108 12180 24110
rect 12124 23938 12180 23940
rect 12124 23886 12126 23938
rect 12126 23886 12178 23938
rect 12178 23886 12180 23938
rect 12124 23884 12180 23886
rect 11676 23100 11732 23156
rect 11340 22988 11396 23044
rect 11116 21644 11172 21700
rect 10892 20188 10948 20244
rect 10892 18450 10948 18452
rect 10892 18398 10894 18450
rect 10894 18398 10946 18450
rect 10946 18398 10948 18450
rect 10892 18396 10948 18398
rect 10780 18172 10836 18228
rect 10444 18060 10500 18116
rect 10108 17276 10164 17332
rect 9324 16828 9380 16884
rect 9884 16828 9940 16884
rect 8876 16716 8932 16772
rect 9660 16716 9716 16772
rect 8764 16604 8820 16660
rect 8540 16098 8596 16100
rect 8540 16046 8542 16098
rect 8542 16046 8594 16098
rect 8594 16046 8596 16098
rect 8540 16044 8596 16046
rect 8428 15372 8484 15428
rect 9660 16044 9716 16100
rect 8204 14812 8260 14868
rect 8428 14588 8484 14644
rect 8540 14530 8596 14532
rect 8540 14478 8542 14530
rect 8542 14478 8594 14530
rect 8594 14478 8596 14530
rect 8540 14476 8596 14478
rect 7756 13746 7812 13748
rect 7756 13694 7758 13746
rect 7758 13694 7810 13746
rect 7810 13694 7812 13746
rect 7756 13692 7812 13694
rect 7980 13858 8036 13860
rect 7980 13806 7982 13858
rect 7982 13806 8034 13858
rect 8034 13806 8036 13858
rect 7980 13804 8036 13806
rect 7980 11676 8036 11732
rect 7868 11116 7924 11172
rect 9436 15874 9492 15876
rect 9436 15822 9438 15874
rect 9438 15822 9490 15874
rect 9490 15822 9492 15874
rect 9436 15820 9492 15822
rect 9660 15426 9716 15428
rect 9660 15374 9662 15426
rect 9662 15374 9714 15426
rect 9714 15374 9716 15426
rect 9660 15372 9716 15374
rect 10332 16940 10388 16996
rect 10892 17164 10948 17220
rect 10444 16828 10500 16884
rect 10780 16044 10836 16100
rect 10108 15036 10164 15092
rect 10556 15874 10612 15876
rect 10556 15822 10558 15874
rect 10558 15822 10610 15874
rect 10610 15822 10612 15874
rect 10556 15820 10612 15822
rect 11564 22428 11620 22484
rect 12124 23154 12180 23156
rect 12124 23102 12126 23154
rect 12126 23102 12178 23154
rect 12178 23102 12180 23154
rect 12124 23100 12180 23102
rect 11788 22988 11844 23044
rect 11340 20076 11396 20132
rect 11228 18060 11284 18116
rect 11340 18396 11396 18452
rect 11116 17836 11172 17892
rect 11116 17500 11172 17556
rect 10332 14700 10388 14756
rect 11004 14642 11060 14644
rect 11004 14590 11006 14642
rect 11006 14590 11058 14642
rect 11058 14590 11060 14642
rect 11004 14588 11060 14590
rect 11116 14252 11172 14308
rect 9884 13692 9940 13748
rect 9212 13468 9268 13524
rect 8764 12850 8820 12852
rect 8764 12798 8766 12850
rect 8766 12798 8818 12850
rect 8818 12798 8820 12850
rect 8764 12796 8820 12798
rect 11564 19964 11620 20020
rect 11340 17612 11396 17668
rect 11564 18284 11620 18340
rect 11788 17890 11844 17892
rect 11788 17838 11790 17890
rect 11790 17838 11842 17890
rect 11842 17838 11844 17890
rect 11788 17836 11844 17838
rect 11676 17612 11732 17668
rect 12124 20802 12180 20804
rect 12124 20750 12126 20802
rect 12126 20750 12178 20802
rect 12178 20750 12180 20802
rect 12124 20748 12180 20750
rect 12460 24892 12516 24948
rect 12460 24556 12516 24612
rect 12684 24332 12740 24388
rect 12684 23884 12740 23940
rect 12572 23042 12628 23044
rect 12572 22990 12574 23042
rect 12574 22990 12626 23042
rect 12626 22990 12628 23042
rect 12572 22988 12628 22990
rect 13468 30380 13524 30436
rect 13356 29202 13412 29204
rect 13356 29150 13358 29202
rect 13358 29150 13410 29202
rect 13410 29150 13412 29202
rect 13356 29148 13412 29150
rect 12908 25506 12964 25508
rect 12908 25454 12910 25506
rect 12910 25454 12962 25506
rect 12962 25454 12964 25506
rect 12908 25452 12964 25454
rect 15260 33180 15316 33236
rect 14588 30828 14644 30884
rect 13692 29202 13748 29204
rect 13692 29150 13694 29202
rect 13694 29150 13746 29202
rect 13746 29150 13748 29202
rect 13692 29148 13748 29150
rect 14812 30604 14868 30660
rect 14028 30380 14084 30436
rect 13916 30044 13972 30100
rect 13916 29538 13972 29540
rect 13916 29486 13918 29538
rect 13918 29486 13970 29538
rect 13970 29486 13972 29538
rect 13916 29484 13972 29486
rect 13580 27916 13636 27972
rect 13580 27132 13636 27188
rect 13804 26290 13860 26292
rect 13804 26238 13806 26290
rect 13806 26238 13858 26290
rect 13858 26238 13860 26290
rect 13804 26236 13860 26238
rect 14364 28588 14420 28644
rect 15260 31778 15316 31780
rect 15260 31726 15262 31778
rect 15262 31726 15314 31778
rect 15314 31726 15316 31778
rect 15260 31724 15316 31726
rect 16044 33234 16100 33236
rect 16044 33182 16046 33234
rect 16046 33182 16098 33234
rect 16098 33182 16100 33234
rect 16044 33180 16100 33182
rect 15372 31388 15428 31444
rect 15932 32396 15988 32452
rect 15820 31164 15876 31220
rect 15484 31052 15540 31108
rect 15372 30604 15428 30660
rect 15708 29596 15764 29652
rect 15260 29148 15316 29204
rect 14140 27970 14196 27972
rect 14140 27918 14142 27970
rect 14142 27918 14194 27970
rect 14194 27918 14196 27970
rect 14140 27916 14196 27918
rect 14476 27970 14532 27972
rect 14476 27918 14478 27970
rect 14478 27918 14530 27970
rect 14530 27918 14532 27970
rect 14476 27916 14532 27918
rect 14812 28252 14868 28308
rect 14924 28642 14980 28644
rect 14924 28590 14926 28642
rect 14926 28590 14978 28642
rect 14978 28590 14980 28642
rect 14924 28588 14980 28590
rect 14588 27468 14644 27524
rect 14476 27132 14532 27188
rect 14028 25900 14084 25956
rect 13580 25452 13636 25508
rect 13804 25228 13860 25284
rect 13468 24892 13524 24948
rect 13468 24556 13524 24612
rect 13356 24332 13412 24388
rect 12908 23660 12964 23716
rect 12460 22370 12516 22372
rect 12460 22318 12462 22370
rect 12462 22318 12514 22370
rect 12514 22318 12516 22370
rect 12460 22316 12516 22318
rect 12796 22540 12852 22596
rect 12684 20748 12740 20804
rect 12908 22482 12964 22484
rect 12908 22430 12910 22482
rect 12910 22430 12962 22482
rect 12962 22430 12964 22482
rect 12908 22428 12964 22430
rect 13020 21756 13076 21812
rect 13132 22764 13188 22820
rect 13580 24050 13636 24052
rect 13580 23998 13582 24050
rect 13582 23998 13634 24050
rect 13634 23998 13636 24050
rect 13580 23996 13636 23998
rect 13468 23100 13524 23156
rect 14252 24946 14308 24948
rect 14252 24894 14254 24946
rect 14254 24894 14306 24946
rect 14306 24894 14308 24946
rect 14252 24892 14308 24894
rect 14476 26290 14532 26292
rect 14476 26238 14478 26290
rect 14478 26238 14530 26290
rect 14530 26238 14532 26290
rect 14476 26236 14532 26238
rect 14364 24444 14420 24500
rect 14476 25900 14532 25956
rect 14140 23996 14196 24052
rect 13916 22764 13972 22820
rect 14028 22204 14084 22260
rect 13580 21756 13636 21812
rect 14028 21644 14084 21700
rect 13580 21084 13636 21140
rect 13804 20802 13860 20804
rect 13804 20750 13806 20802
rect 13806 20750 13858 20802
rect 13858 20750 13860 20802
rect 13804 20748 13860 20750
rect 12124 18396 12180 18452
rect 12348 18450 12404 18452
rect 12348 18398 12350 18450
rect 12350 18398 12402 18450
rect 12402 18398 12404 18450
rect 12348 18396 12404 18398
rect 12012 18060 12068 18116
rect 12460 17724 12516 17780
rect 12012 17164 12068 17220
rect 11900 16994 11956 16996
rect 11900 16942 11902 16994
rect 11902 16942 11954 16994
rect 11954 16942 11956 16994
rect 11900 16940 11956 16942
rect 12124 16658 12180 16660
rect 12124 16606 12126 16658
rect 12126 16606 12178 16658
rect 12178 16606 12180 16658
rect 12124 16604 12180 16606
rect 11564 15820 11620 15876
rect 11676 15314 11732 15316
rect 11676 15262 11678 15314
rect 11678 15262 11730 15314
rect 11730 15262 11732 15314
rect 11676 15260 11732 15262
rect 11564 15036 11620 15092
rect 12460 17500 12516 17556
rect 12796 20076 12852 20132
rect 13356 20076 13412 20132
rect 14924 27132 14980 27188
rect 15036 27468 15092 27524
rect 15036 27020 15092 27076
rect 14924 26290 14980 26292
rect 14924 26238 14926 26290
rect 14926 26238 14978 26290
rect 14978 26238 14980 26290
rect 14924 26236 14980 26238
rect 15372 26908 15428 26964
rect 14812 25228 14868 25284
rect 14924 25900 14980 25956
rect 16492 33234 16548 33236
rect 16492 33182 16494 33234
rect 16494 33182 16546 33234
rect 16546 33182 16548 33234
rect 16492 33180 16548 33182
rect 16380 31836 16436 31892
rect 16828 34130 16884 34132
rect 16828 34078 16830 34130
rect 16830 34078 16882 34130
rect 16882 34078 16884 34130
rect 16828 34076 16884 34078
rect 16604 31052 16660 31108
rect 16380 29596 16436 29652
rect 17724 38220 17780 38276
rect 17724 37938 17780 37940
rect 17724 37886 17726 37938
rect 17726 37886 17778 37938
rect 17778 37886 17780 37938
rect 17724 37884 17780 37886
rect 17500 36988 17556 37044
rect 17612 37772 17668 37828
rect 17388 34354 17444 34356
rect 17388 34302 17390 34354
rect 17390 34302 17442 34354
rect 17442 34302 17444 34354
rect 17388 34300 17444 34302
rect 17276 33964 17332 34020
rect 17052 29372 17108 29428
rect 16156 28476 16212 28532
rect 16604 29148 16660 29204
rect 17052 28700 17108 28756
rect 16940 28642 16996 28644
rect 16940 28590 16942 28642
rect 16942 28590 16994 28642
rect 16994 28590 16996 28642
rect 16940 28588 16996 28590
rect 17500 31218 17556 31220
rect 17500 31166 17502 31218
rect 17502 31166 17554 31218
rect 17554 31166 17556 31218
rect 17500 31164 17556 31166
rect 17388 31106 17444 31108
rect 17388 31054 17390 31106
rect 17390 31054 17442 31106
rect 17442 31054 17444 31106
rect 17388 31052 17444 31054
rect 17276 29484 17332 29540
rect 17388 28754 17444 28756
rect 17388 28702 17390 28754
rect 17390 28702 17442 28754
rect 17442 28702 17444 28754
rect 17388 28700 17444 28702
rect 16940 28364 16996 28420
rect 16828 27804 16884 27860
rect 16716 27580 16772 27636
rect 15372 25788 15428 25844
rect 14700 24722 14756 24724
rect 14700 24670 14702 24722
rect 14702 24670 14754 24722
rect 14754 24670 14756 24722
rect 14700 24668 14756 24670
rect 14700 24444 14756 24500
rect 14476 23660 14532 23716
rect 14700 23660 14756 23716
rect 14364 21756 14420 21812
rect 15036 23996 15092 24052
rect 16156 25228 16212 25284
rect 15484 23826 15540 23828
rect 15484 23774 15486 23826
rect 15486 23774 15538 23826
rect 15538 23774 15540 23826
rect 15484 23772 15540 23774
rect 14812 21308 14868 21364
rect 14476 21196 14532 21252
rect 14140 20690 14196 20692
rect 14140 20638 14142 20690
rect 14142 20638 14194 20690
rect 14194 20638 14196 20690
rect 14140 20636 14196 20638
rect 14364 20188 14420 20244
rect 13468 19010 13524 19012
rect 13468 18958 13470 19010
rect 13470 18958 13522 19010
rect 13522 18958 13524 19010
rect 13468 18956 13524 18958
rect 14364 19068 14420 19124
rect 13916 18956 13972 19012
rect 13804 18338 13860 18340
rect 13804 18286 13806 18338
rect 13806 18286 13858 18338
rect 13858 18286 13860 18338
rect 13804 18284 13860 18286
rect 13020 18060 13076 18116
rect 12684 16940 12740 16996
rect 12796 15372 12852 15428
rect 12236 14588 12292 14644
rect 11228 12796 11284 12852
rect 8764 11676 8820 11732
rect 8876 12684 8932 12740
rect 7644 9714 7700 9716
rect 7644 9662 7646 9714
rect 7646 9662 7698 9714
rect 7698 9662 7700 9714
rect 7644 9660 7700 9662
rect 8204 9660 8260 9716
rect 8316 9042 8372 9044
rect 8316 8990 8318 9042
rect 8318 8990 8370 9042
rect 8370 8990 8372 9042
rect 8316 8988 8372 8990
rect 7532 7644 7588 7700
rect 8652 10610 8708 10612
rect 8652 10558 8654 10610
rect 8654 10558 8706 10610
rect 8706 10558 8708 10610
rect 8652 10556 8708 10558
rect 8540 9714 8596 9716
rect 8540 9662 8542 9714
rect 8542 9662 8594 9714
rect 8594 9662 8596 9714
rect 8540 9660 8596 9662
rect 7532 6578 7588 6580
rect 7532 6526 7534 6578
rect 7534 6526 7586 6578
rect 7586 6526 7588 6578
rect 7532 6524 7588 6526
rect 8204 7698 8260 7700
rect 8204 7646 8206 7698
rect 8206 7646 8258 7698
rect 8258 7646 8260 7698
rect 8204 7644 8260 7646
rect 8540 7362 8596 7364
rect 8540 7310 8542 7362
rect 8542 7310 8594 7362
rect 8594 7310 8596 7362
rect 8540 7308 8596 7310
rect 11340 14252 11396 14308
rect 12012 13916 12068 13972
rect 12124 12738 12180 12740
rect 12124 12686 12126 12738
rect 12126 12686 12178 12738
rect 12178 12686 12180 12738
rect 12124 12684 12180 12686
rect 12348 12124 12404 12180
rect 9324 10892 9380 10948
rect 9660 10610 9716 10612
rect 9660 10558 9662 10610
rect 9662 10558 9714 10610
rect 9714 10558 9716 10610
rect 9660 10556 9716 10558
rect 11452 10556 11508 10612
rect 10892 10332 10948 10388
rect 12460 10498 12516 10500
rect 12460 10446 12462 10498
rect 12462 10446 12514 10498
rect 12514 10446 12516 10498
rect 12460 10444 12516 10446
rect 11452 9884 11508 9940
rect 11004 9548 11060 9604
rect 9436 8988 9492 9044
rect 9660 8652 9716 8708
rect 9324 7644 9380 7700
rect 10780 8092 10836 8148
rect 10444 7474 10500 7476
rect 10444 7422 10446 7474
rect 10446 7422 10498 7474
rect 10498 7422 10500 7474
rect 10444 7420 10500 7422
rect 8988 7308 9044 7364
rect 8204 6748 8260 6804
rect 8988 6972 9044 7028
rect 7532 5122 7588 5124
rect 7532 5070 7534 5122
rect 7534 5070 7586 5122
rect 7586 5070 7588 5122
rect 7532 5068 7588 5070
rect 7420 4956 7476 5012
rect 7644 4844 7700 4900
rect 7196 3948 7252 4004
rect 6972 3724 7028 3780
rect 8204 4284 8260 4340
rect 8540 6748 8596 6804
rect 9772 7362 9828 7364
rect 9772 7310 9774 7362
rect 9774 7310 9826 7362
rect 9826 7310 9828 7362
rect 9772 7308 9828 7310
rect 8764 6188 8820 6244
rect 8316 3612 8372 3668
rect 8988 6076 9044 6132
rect 8876 5852 8932 5908
rect 9212 6188 9268 6244
rect 9660 6524 9716 6580
rect 10220 6860 10276 6916
rect 9884 6690 9940 6692
rect 9884 6638 9886 6690
rect 9886 6638 9938 6690
rect 9938 6638 9940 6690
rect 9884 6636 9940 6638
rect 10668 6690 10724 6692
rect 10668 6638 10670 6690
rect 10670 6638 10722 6690
rect 10722 6638 10724 6690
rect 10668 6636 10724 6638
rect 9996 6300 10052 6356
rect 9884 5852 9940 5908
rect 9324 3666 9380 3668
rect 9324 3614 9326 3666
rect 9326 3614 9378 3666
rect 9378 3614 9380 3666
rect 9324 3612 9380 3614
rect 7868 3442 7924 3444
rect 7868 3390 7870 3442
rect 7870 3390 7922 3442
rect 7922 3390 7924 3442
rect 7868 3388 7924 3390
rect 9772 5516 9828 5572
rect 10668 5404 10724 5460
rect 10444 5292 10500 5348
rect 10444 5068 10500 5124
rect 10220 4338 10276 4340
rect 10220 4286 10222 4338
rect 10222 4286 10274 4338
rect 10274 4286 10276 4338
rect 10220 4284 10276 4286
rect 10556 4450 10612 4452
rect 10556 4398 10558 4450
rect 10558 4398 10610 4450
rect 10610 4398 10612 4450
rect 10556 4396 10612 4398
rect 12348 9602 12404 9604
rect 12348 9550 12350 9602
rect 12350 9550 12402 9602
rect 12402 9550 12404 9602
rect 12348 9548 12404 9550
rect 11900 8540 11956 8596
rect 11004 6076 11060 6132
rect 11004 5906 11060 5908
rect 11004 5854 11006 5906
rect 11006 5854 11058 5906
rect 11058 5854 11060 5906
rect 11004 5852 11060 5854
rect 11340 6636 11396 6692
rect 11564 7196 11620 7252
rect 11788 7474 11844 7476
rect 11788 7422 11790 7474
rect 11790 7422 11842 7474
rect 11842 7422 11844 7474
rect 11788 7420 11844 7422
rect 11788 6748 11844 6804
rect 11788 5628 11844 5684
rect 11788 4508 11844 4564
rect 13804 17948 13860 18004
rect 13580 17778 13636 17780
rect 13580 17726 13582 17778
rect 13582 17726 13634 17778
rect 13634 17726 13636 17778
rect 13580 17724 13636 17726
rect 13804 17554 13860 17556
rect 13804 17502 13806 17554
rect 13806 17502 13858 17554
rect 13858 17502 13860 17554
rect 13804 17500 13860 17502
rect 14252 18450 14308 18452
rect 14252 18398 14254 18450
rect 14254 18398 14306 18450
rect 14306 18398 14308 18450
rect 14252 18396 14308 18398
rect 14028 18226 14084 18228
rect 14028 18174 14030 18226
rect 14030 18174 14082 18226
rect 14082 18174 14084 18226
rect 14028 18172 14084 18174
rect 14252 17724 14308 17780
rect 13468 17442 13524 17444
rect 13468 17390 13470 17442
rect 13470 17390 13522 17442
rect 13522 17390 13524 17442
rect 13468 17388 13524 17390
rect 13468 17164 13524 17220
rect 14924 22428 14980 22484
rect 14924 21868 14980 21924
rect 14812 20802 14868 20804
rect 14812 20750 14814 20802
rect 14814 20750 14866 20802
rect 14866 20750 14868 20802
rect 14812 20748 14868 20750
rect 14700 20018 14756 20020
rect 14700 19966 14702 20018
rect 14702 19966 14754 20018
rect 14754 19966 14756 20018
rect 14700 19964 14756 19966
rect 15148 21084 15204 21140
rect 15148 20130 15204 20132
rect 15148 20078 15150 20130
rect 15150 20078 15202 20130
rect 15202 20078 15204 20130
rect 15148 20076 15204 20078
rect 15820 19628 15876 19684
rect 14700 18450 14756 18452
rect 14700 18398 14702 18450
rect 14702 18398 14754 18450
rect 14754 18398 14756 18450
rect 14700 18396 14756 18398
rect 14700 17948 14756 18004
rect 14588 17164 14644 17220
rect 14812 17612 14868 17668
rect 14588 16994 14644 16996
rect 14588 16942 14590 16994
rect 14590 16942 14642 16994
rect 14642 16942 14644 16994
rect 14588 16940 14644 16942
rect 15708 18450 15764 18452
rect 15708 18398 15710 18450
rect 15710 18398 15762 18450
rect 15762 18398 15764 18450
rect 15708 18396 15764 18398
rect 16380 24108 16436 24164
rect 17164 26962 17220 26964
rect 17164 26910 17166 26962
rect 17166 26910 17218 26962
rect 17218 26910 17220 26962
rect 17164 26908 17220 26910
rect 17836 36988 17892 37044
rect 18060 38834 18116 38836
rect 18060 38782 18062 38834
rect 18062 38782 18114 38834
rect 18114 38782 18116 38834
rect 18060 38780 18116 38782
rect 18284 42028 18340 42084
rect 18396 41916 18452 41972
rect 20076 48300 20132 48356
rect 19852 47964 19908 48020
rect 20748 47964 20804 48020
rect 21308 48018 21364 48020
rect 21308 47966 21310 48018
rect 21310 47966 21362 48018
rect 21362 47966 21364 48018
rect 21308 47964 21364 47966
rect 19292 47292 19348 47348
rect 21532 48354 21588 48356
rect 21532 48302 21534 48354
rect 21534 48302 21586 48354
rect 21586 48302 21588 48354
rect 21532 48300 21588 48302
rect 21980 48354 22036 48356
rect 21980 48302 21982 48354
rect 21982 48302 22034 48354
rect 22034 48302 22036 48354
rect 21980 48300 22036 48302
rect 22652 48354 22708 48356
rect 22652 48302 22654 48354
rect 22654 48302 22706 48354
rect 22706 48302 22708 48354
rect 22652 48300 22708 48302
rect 21980 47964 22036 48020
rect 21420 47180 21476 47236
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 18732 46060 18788 46116
rect 19628 46060 19684 46116
rect 21196 46060 21252 46116
rect 19292 45388 19348 45444
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19180 44828 19236 44884
rect 20748 45836 20804 45892
rect 21868 45890 21924 45892
rect 21868 45838 21870 45890
rect 21870 45838 21922 45890
rect 21922 45838 21924 45890
rect 21868 45836 21924 45838
rect 20972 44268 21028 44324
rect 19404 43596 19460 43652
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20188 42924 20244 42980
rect 20412 43596 20468 43652
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 18508 39004 18564 39060
rect 18172 37436 18228 37492
rect 18620 38668 18676 38724
rect 18844 38834 18900 38836
rect 18844 38782 18846 38834
rect 18846 38782 18898 38834
rect 18898 38782 18900 38834
rect 18844 38780 18900 38782
rect 18284 36204 18340 36260
rect 17948 34972 18004 35028
rect 18172 35586 18228 35588
rect 18172 35534 18174 35586
rect 18174 35534 18226 35586
rect 18226 35534 18228 35586
rect 18172 35532 18228 35534
rect 18060 34914 18116 34916
rect 18060 34862 18062 34914
rect 18062 34862 18114 34914
rect 18114 34862 18116 34914
rect 18060 34860 18116 34862
rect 18732 37100 18788 37156
rect 18508 36370 18564 36372
rect 18508 36318 18510 36370
rect 18510 36318 18562 36370
rect 18562 36318 18564 36370
rect 18508 36316 18564 36318
rect 19180 41970 19236 41972
rect 19180 41918 19182 41970
rect 19182 41918 19234 41970
rect 19234 41918 19236 41970
rect 19180 41916 19236 41918
rect 19180 41298 19236 41300
rect 19180 41246 19182 41298
rect 19182 41246 19234 41298
rect 19234 41246 19236 41298
rect 19180 41244 19236 41246
rect 19628 41916 19684 41972
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19180 40402 19236 40404
rect 19180 40350 19182 40402
rect 19182 40350 19234 40402
rect 19234 40350 19236 40402
rect 19180 40348 19236 40350
rect 20188 40402 20244 40404
rect 20188 40350 20190 40402
rect 20190 40350 20242 40402
rect 20242 40350 20244 40402
rect 20188 40348 20244 40350
rect 19068 38556 19124 38612
rect 19068 38220 19124 38276
rect 20188 39564 20244 39620
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19516 38834 19572 38836
rect 19516 38782 19518 38834
rect 19518 38782 19570 38834
rect 19570 38782 19572 38834
rect 19516 38780 19572 38782
rect 19292 38556 19348 38612
rect 20076 38556 20132 38612
rect 19180 38050 19236 38052
rect 19180 37998 19182 38050
rect 19182 37998 19234 38050
rect 19234 37998 19236 38050
rect 19180 37996 19236 37998
rect 19628 37884 19684 37940
rect 19404 37826 19460 37828
rect 19404 37774 19406 37826
rect 19406 37774 19458 37826
rect 19458 37774 19460 37826
rect 19404 37772 19460 37774
rect 19404 36876 19460 36932
rect 18844 36764 18900 36820
rect 19292 36764 19348 36820
rect 19068 36652 19124 36708
rect 18956 36370 19012 36372
rect 18956 36318 18958 36370
rect 18958 36318 19010 36370
rect 19010 36318 19012 36370
rect 18956 36316 19012 36318
rect 18844 36258 18900 36260
rect 18844 36206 18846 36258
rect 18846 36206 18898 36258
rect 18898 36206 18900 36258
rect 18844 36204 18900 36206
rect 18732 35868 18788 35924
rect 18396 35420 18452 35476
rect 18620 35644 18676 35700
rect 18956 36092 19012 36148
rect 18844 35196 18900 35252
rect 18620 34914 18676 34916
rect 18620 34862 18622 34914
rect 18622 34862 18674 34914
rect 18674 34862 18676 34914
rect 18620 34860 18676 34862
rect 18956 34914 19012 34916
rect 18956 34862 18958 34914
rect 18958 34862 19010 34914
rect 19010 34862 19012 34914
rect 18956 34860 19012 34862
rect 19852 37826 19908 37828
rect 19852 37774 19854 37826
rect 19854 37774 19906 37826
rect 19906 37774 19908 37826
rect 19852 37772 19908 37774
rect 20076 37772 20132 37828
rect 19628 37660 19684 37716
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20076 37100 20132 37156
rect 19516 36428 19572 36484
rect 19628 36540 19684 36596
rect 19964 36204 20020 36260
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19628 35644 19684 35700
rect 21420 42978 21476 42980
rect 21420 42926 21422 42978
rect 21422 42926 21474 42978
rect 21474 42926 21476 42978
rect 21420 42924 21476 42926
rect 21756 41804 21812 41860
rect 21756 40908 21812 40964
rect 20636 39452 20692 39508
rect 20412 37938 20468 37940
rect 20412 37886 20414 37938
rect 20414 37886 20466 37938
rect 20466 37886 20468 37938
rect 20412 37884 20468 37886
rect 20972 38556 21028 38612
rect 20972 37884 21028 37940
rect 20188 35586 20244 35588
rect 20188 35534 20190 35586
rect 20190 35534 20242 35586
rect 20242 35534 20244 35586
rect 20188 35532 20244 35534
rect 20300 37660 20356 37716
rect 19516 35084 19572 35140
rect 20188 35138 20244 35140
rect 20188 35086 20190 35138
rect 20190 35086 20242 35138
rect 20242 35086 20244 35138
rect 20188 35084 20244 35086
rect 18620 34300 18676 34356
rect 17724 32620 17780 32676
rect 17836 33068 17892 33124
rect 17724 31612 17780 31668
rect 17948 32396 18004 32452
rect 18956 34130 19012 34132
rect 18956 34078 18958 34130
rect 18958 34078 19010 34130
rect 19010 34078 19012 34130
rect 18956 34076 19012 34078
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19964 34018 20020 34020
rect 19964 33966 19966 34018
rect 19966 33966 20018 34018
rect 20018 33966 20020 34018
rect 19964 33964 20020 33966
rect 19516 33516 19572 33572
rect 19516 33346 19572 33348
rect 19516 33294 19518 33346
rect 19518 33294 19570 33346
rect 19570 33294 19572 33346
rect 19516 33292 19572 33294
rect 18060 31724 18116 31780
rect 17948 31500 18004 31556
rect 18284 31724 18340 31780
rect 18508 31890 18564 31892
rect 18508 31838 18510 31890
rect 18510 31838 18562 31890
rect 18562 31838 18564 31890
rect 18508 31836 18564 31838
rect 18060 30828 18116 30884
rect 17724 30492 17780 30548
rect 18172 29484 18228 29540
rect 17836 29314 17892 29316
rect 17836 29262 17838 29314
rect 17838 29262 17890 29314
rect 17890 29262 17892 29314
rect 17836 29260 17892 29262
rect 17724 28028 17780 28084
rect 17724 27580 17780 27636
rect 17612 27132 17668 27188
rect 17500 26908 17556 26964
rect 17388 26178 17444 26180
rect 17388 26126 17390 26178
rect 17390 26126 17442 26178
rect 17442 26126 17444 26178
rect 17388 26124 17444 26126
rect 17388 25228 17444 25284
rect 17724 27074 17780 27076
rect 17724 27022 17726 27074
rect 17726 27022 17778 27074
rect 17778 27022 17780 27074
rect 17724 27020 17780 27022
rect 19292 33122 19348 33124
rect 19292 33070 19294 33122
rect 19294 33070 19346 33122
rect 19346 33070 19348 33122
rect 19292 33068 19348 33070
rect 20636 36540 20692 36596
rect 21756 39506 21812 39508
rect 21756 39454 21758 39506
rect 21758 39454 21810 39506
rect 21810 39454 21812 39506
rect 21756 39452 21812 39454
rect 21644 39228 21700 39284
rect 22092 43426 22148 43428
rect 22092 43374 22094 43426
rect 22094 43374 22146 43426
rect 22146 43374 22148 43426
rect 22092 43372 22148 43374
rect 22540 43372 22596 43428
rect 22316 41858 22372 41860
rect 22316 41806 22318 41858
rect 22318 41806 22370 41858
rect 22370 41806 22372 41858
rect 22316 41804 22372 41806
rect 22092 39618 22148 39620
rect 22092 39566 22094 39618
rect 22094 39566 22146 39618
rect 22146 39566 22148 39618
rect 22092 39564 22148 39566
rect 22428 40796 22484 40852
rect 21644 38162 21700 38164
rect 21644 38110 21646 38162
rect 21646 38110 21698 38162
rect 21698 38110 21700 38162
rect 21644 38108 21700 38110
rect 21868 39004 21924 39060
rect 21756 37772 21812 37828
rect 21308 37154 21364 37156
rect 21308 37102 21310 37154
rect 21310 37102 21362 37154
rect 21362 37102 21364 37154
rect 21308 37100 21364 37102
rect 20972 36988 21028 37044
rect 20748 36428 20804 36484
rect 21420 36370 21476 36372
rect 21420 36318 21422 36370
rect 21422 36318 21474 36370
rect 21474 36318 21476 36370
rect 21420 36316 21476 36318
rect 20860 36258 20916 36260
rect 20860 36206 20862 36258
rect 20862 36206 20914 36258
rect 20914 36206 20916 36258
rect 20860 36204 20916 36206
rect 20636 34412 20692 34468
rect 20524 33404 20580 33460
rect 20300 33292 20356 33348
rect 19836 32954 19892 32956
rect 19180 32844 19236 32900
rect 19628 32844 19684 32900
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 18844 32450 18900 32452
rect 18844 32398 18846 32450
rect 18846 32398 18898 32450
rect 18898 32398 18900 32450
rect 18844 32396 18900 32398
rect 18732 31724 18788 31780
rect 18844 31500 18900 31556
rect 20188 32844 20244 32900
rect 20636 32172 20692 32228
rect 19964 31778 20020 31780
rect 19964 31726 19966 31778
rect 19966 31726 20018 31778
rect 20018 31726 20020 31778
rect 19964 31724 20020 31726
rect 19628 31612 19684 31668
rect 19404 31554 19460 31556
rect 19404 31502 19406 31554
rect 19406 31502 19458 31554
rect 19458 31502 19460 31554
rect 19404 31500 19460 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 18396 29036 18452 29092
rect 18620 29538 18676 29540
rect 18620 29486 18622 29538
rect 18622 29486 18674 29538
rect 18674 29486 18676 29538
rect 18620 29484 18676 29486
rect 18508 28364 18564 28420
rect 18620 28082 18676 28084
rect 18620 28030 18622 28082
rect 18622 28030 18674 28082
rect 18674 28030 18676 28082
rect 18620 28028 18676 28030
rect 18060 25564 18116 25620
rect 18508 27692 18564 27748
rect 18284 25900 18340 25956
rect 18396 25506 18452 25508
rect 18396 25454 18398 25506
rect 18398 25454 18450 25506
rect 18450 25454 18452 25506
rect 18396 25452 18452 25454
rect 20412 31666 20468 31668
rect 20412 31614 20414 31666
rect 20414 31614 20466 31666
rect 20466 31614 20468 31666
rect 20412 31612 20468 31614
rect 20636 31666 20692 31668
rect 20636 31614 20638 31666
rect 20638 31614 20690 31666
rect 20690 31614 20692 31666
rect 20636 31612 20692 31614
rect 19740 30828 19796 30884
rect 19068 30604 19124 30660
rect 19740 30268 19796 30324
rect 19404 30156 19460 30212
rect 18844 29932 18900 29988
rect 19180 29538 19236 29540
rect 19180 29486 19182 29538
rect 19182 29486 19234 29538
rect 19234 29486 19236 29538
rect 19180 29484 19236 29486
rect 18844 28028 18900 28084
rect 18956 28812 19012 28868
rect 18732 25564 18788 25620
rect 18844 25340 18900 25396
rect 16268 22092 16324 22148
rect 16716 23548 16772 23604
rect 17164 23714 17220 23716
rect 17164 23662 17166 23714
rect 17166 23662 17218 23714
rect 17218 23662 17220 23714
rect 17164 23660 17220 23662
rect 16940 23100 16996 23156
rect 16492 22316 16548 22372
rect 17052 20578 17108 20580
rect 17052 20526 17054 20578
rect 17054 20526 17106 20578
rect 17106 20526 17108 20578
rect 17052 20524 17108 20526
rect 16380 19964 16436 20020
rect 16156 18060 16212 18116
rect 15820 17836 15876 17892
rect 17388 23660 17444 23716
rect 17724 23772 17780 23828
rect 17612 23714 17668 23716
rect 17612 23662 17614 23714
rect 17614 23662 17666 23714
rect 17666 23662 17668 23714
rect 17612 23660 17668 23662
rect 17500 23324 17556 23380
rect 17388 23154 17444 23156
rect 17388 23102 17390 23154
rect 17390 23102 17442 23154
rect 17442 23102 17444 23154
rect 17388 23100 17444 23102
rect 17500 22764 17556 22820
rect 17388 22482 17444 22484
rect 17388 22430 17390 22482
rect 17390 22430 17442 22482
rect 17442 22430 17444 22482
rect 17388 22428 17444 22430
rect 18060 25004 18116 25060
rect 18172 24332 18228 24388
rect 17948 23436 18004 23492
rect 18172 23212 18228 23268
rect 19292 28588 19348 28644
rect 19068 28028 19124 28084
rect 19404 28028 19460 28084
rect 19516 28812 19572 28868
rect 20076 30210 20132 30212
rect 20076 30158 20078 30210
rect 20078 30158 20130 30210
rect 20130 30158 20132 30210
rect 20076 30156 20132 30158
rect 19852 29932 19908 29988
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19740 28642 19796 28644
rect 19740 28590 19742 28642
rect 19742 28590 19794 28642
rect 19794 28590 19796 28642
rect 19740 28588 19796 28590
rect 19516 27804 19572 27860
rect 19292 26178 19348 26180
rect 19292 26126 19294 26178
rect 19294 26126 19346 26178
rect 19346 26126 19348 26178
rect 19292 26124 19348 26126
rect 21084 35532 21140 35588
rect 21644 35922 21700 35924
rect 21644 35870 21646 35922
rect 21646 35870 21698 35922
rect 21698 35870 21700 35922
rect 21644 35868 21700 35870
rect 21532 34412 21588 34468
rect 21644 35644 21700 35700
rect 20860 32844 20916 32900
rect 21308 32844 21364 32900
rect 21308 32450 21364 32452
rect 21308 32398 21310 32450
rect 21310 32398 21362 32450
rect 21362 32398 21364 32450
rect 21308 32396 21364 32398
rect 20860 29986 20916 29988
rect 20860 29934 20862 29986
rect 20862 29934 20914 29986
rect 20914 29934 20916 29986
rect 20860 29932 20916 29934
rect 22204 37996 22260 38052
rect 21980 37826 22036 37828
rect 21980 37774 21982 37826
rect 21982 37774 22034 37826
rect 22034 37774 22036 37826
rect 21980 37772 22036 37774
rect 24332 48300 24388 48356
rect 29260 49026 29316 49028
rect 29260 48974 29262 49026
rect 29262 48974 29314 49026
rect 29314 48974 29316 49026
rect 29260 48972 29316 48974
rect 25676 48300 25732 48356
rect 22988 47234 23044 47236
rect 22988 47182 22990 47234
rect 22990 47182 23042 47234
rect 23042 47182 23044 47234
rect 22988 47180 23044 47182
rect 24444 46844 24500 46900
rect 25340 46898 25396 46900
rect 25340 46846 25342 46898
rect 25342 46846 25394 46898
rect 25394 46846 25396 46898
rect 25340 46844 25396 46846
rect 28252 48354 28308 48356
rect 28252 48302 28254 48354
rect 28254 48302 28306 48354
rect 28306 48302 28308 48354
rect 28252 48300 28308 48302
rect 26908 48076 26964 48132
rect 22764 45612 22820 45668
rect 24332 45666 24388 45668
rect 24332 45614 24334 45666
rect 24334 45614 24386 45666
rect 24386 45614 24388 45666
rect 24332 45612 24388 45614
rect 25788 44828 25844 44884
rect 23324 44322 23380 44324
rect 23324 44270 23326 44322
rect 23326 44270 23378 44322
rect 23378 44270 23380 44322
rect 23324 44268 23380 44270
rect 25676 44044 25732 44100
rect 24556 42754 24612 42756
rect 24556 42702 24558 42754
rect 24558 42702 24610 42754
rect 24610 42702 24612 42754
rect 24556 42700 24612 42702
rect 25228 42700 25284 42756
rect 25564 42028 25620 42084
rect 24444 41074 24500 41076
rect 24444 41022 24446 41074
rect 24446 41022 24498 41074
rect 24498 41022 24500 41074
rect 24444 41020 24500 41022
rect 25340 41020 25396 41076
rect 23100 40962 23156 40964
rect 23100 40910 23102 40962
rect 23102 40910 23154 40962
rect 23154 40910 23156 40962
rect 23100 40908 23156 40910
rect 22764 39564 22820 39620
rect 22652 39004 22708 39060
rect 22988 38162 23044 38164
rect 22988 38110 22990 38162
rect 22990 38110 23042 38162
rect 23042 38110 23044 38162
rect 22988 38108 23044 38110
rect 23324 38668 23380 38724
rect 23324 38108 23380 38164
rect 22204 36988 22260 37044
rect 22204 35810 22260 35812
rect 22204 35758 22206 35810
rect 22206 35758 22258 35810
rect 22258 35758 22260 35810
rect 22204 35756 22260 35758
rect 22540 36482 22596 36484
rect 22540 36430 22542 36482
rect 22542 36430 22594 36482
rect 22594 36430 22596 36482
rect 22540 36428 22596 36430
rect 21980 34972 22036 35028
rect 21756 32508 21812 32564
rect 22092 32620 22148 32676
rect 21644 29484 21700 29540
rect 20748 28530 20804 28532
rect 20748 28478 20750 28530
rect 20750 28478 20802 28530
rect 20802 28478 20804 28530
rect 20748 28476 20804 28478
rect 20636 28364 20692 28420
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19628 27132 19684 27188
rect 20860 27132 20916 27188
rect 19740 27074 19796 27076
rect 19740 27022 19742 27074
rect 19742 27022 19794 27074
rect 19794 27022 19796 27074
rect 19740 27020 19796 27022
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20188 26572 20244 26628
rect 19740 25564 19796 25620
rect 19292 25394 19348 25396
rect 19292 25342 19294 25394
rect 19294 25342 19346 25394
rect 19346 25342 19348 25394
rect 19292 25340 19348 25342
rect 19180 25282 19236 25284
rect 19180 25230 19182 25282
rect 19182 25230 19234 25282
rect 19234 25230 19236 25282
rect 19180 25228 19236 25230
rect 19964 25452 20020 25508
rect 19852 25228 19908 25284
rect 20748 26572 20804 26628
rect 20300 25564 20356 25620
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19068 24892 19124 24948
rect 20748 24946 20804 24948
rect 20748 24894 20750 24946
rect 20750 24894 20802 24946
rect 20802 24894 20804 24946
rect 20748 24892 20804 24894
rect 21756 31724 21812 31780
rect 21868 31612 21924 31668
rect 21756 29820 21812 29876
rect 21644 28476 21700 28532
rect 21980 28364 22036 28420
rect 22092 27244 22148 27300
rect 21756 27132 21812 27188
rect 21308 26908 21364 26964
rect 21532 26850 21588 26852
rect 21532 26798 21534 26850
rect 21534 26798 21586 26850
rect 21586 26798 21588 26850
rect 21532 26796 21588 26798
rect 21756 26684 21812 26740
rect 23100 36988 23156 37044
rect 22764 35868 22820 35924
rect 22764 35698 22820 35700
rect 22764 35646 22766 35698
rect 22766 35646 22818 35698
rect 22818 35646 22820 35698
rect 22764 35644 22820 35646
rect 23100 35644 23156 35700
rect 22652 35084 22708 35140
rect 22764 34972 22820 35028
rect 23324 36482 23380 36484
rect 23324 36430 23326 36482
rect 23326 36430 23378 36482
rect 23378 36430 23380 36482
rect 23324 36428 23380 36430
rect 23548 40402 23604 40404
rect 23548 40350 23550 40402
rect 23550 40350 23602 40402
rect 23602 40350 23604 40402
rect 23548 40348 23604 40350
rect 24556 40796 24612 40852
rect 24108 38722 24164 38724
rect 24108 38670 24110 38722
rect 24110 38670 24162 38722
rect 24162 38670 24164 38722
rect 24108 38668 24164 38670
rect 24332 39340 24388 39396
rect 24332 38834 24388 38836
rect 24332 38782 24334 38834
rect 24334 38782 24386 38834
rect 24386 38782 24388 38834
rect 24332 38780 24388 38782
rect 24220 38556 24276 38612
rect 23772 38108 23828 38164
rect 24108 38332 24164 38388
rect 24220 37996 24276 38052
rect 25116 40236 25172 40292
rect 24668 38780 24724 38836
rect 24780 39564 24836 39620
rect 24780 37996 24836 38052
rect 24668 37938 24724 37940
rect 24668 37886 24670 37938
rect 24670 37886 24722 37938
rect 24722 37886 24724 37938
rect 24668 37884 24724 37886
rect 24444 37772 24500 37828
rect 25004 38108 25060 38164
rect 23884 36988 23940 37044
rect 25004 36988 25060 37044
rect 24780 36876 24836 36932
rect 24892 36706 24948 36708
rect 24892 36654 24894 36706
rect 24894 36654 24946 36706
rect 24946 36654 24948 36706
rect 24892 36652 24948 36654
rect 24780 36540 24836 36596
rect 23772 36204 23828 36260
rect 23660 35868 23716 35924
rect 23436 35532 23492 35588
rect 23324 35474 23380 35476
rect 23324 35422 23326 35474
rect 23326 35422 23378 35474
rect 23378 35422 23380 35474
rect 23324 35420 23380 35422
rect 23548 35196 23604 35252
rect 22988 34748 23044 34804
rect 24332 36428 24388 36484
rect 25676 40348 25732 40404
rect 25452 38722 25508 38724
rect 25452 38670 25454 38722
rect 25454 38670 25506 38722
rect 25506 38670 25508 38722
rect 25452 38668 25508 38670
rect 25228 38444 25284 38500
rect 25340 38332 25396 38388
rect 25788 38722 25844 38724
rect 25788 38670 25790 38722
rect 25790 38670 25842 38722
rect 25842 38670 25844 38722
rect 25788 38668 25844 38670
rect 27692 48018 27748 48020
rect 27692 47966 27694 48018
rect 27694 47966 27746 48018
rect 27746 47966 27748 48018
rect 27692 47964 27748 47966
rect 26908 46060 26964 46116
rect 27020 45106 27076 45108
rect 27020 45054 27022 45106
rect 27022 45054 27074 45106
rect 27074 45054 27076 45106
rect 27020 45052 27076 45054
rect 27692 46114 27748 46116
rect 27692 46062 27694 46114
rect 27694 46062 27746 46114
rect 27746 46062 27748 46114
rect 27692 46060 27748 46062
rect 26348 44828 26404 44884
rect 27916 44940 27972 44996
rect 26236 44044 26292 44100
rect 26236 42082 26292 42084
rect 26236 42030 26238 42082
rect 26238 42030 26290 42082
rect 26290 42030 26292 42082
rect 26236 42028 26292 42030
rect 26908 42028 26964 42084
rect 32396 48972 32452 49028
rect 30828 48354 30884 48356
rect 30828 48302 30830 48354
rect 30830 48302 30882 48354
rect 30882 48302 30884 48354
rect 30828 48300 30884 48302
rect 30268 48242 30324 48244
rect 30268 48190 30270 48242
rect 30270 48190 30322 48242
rect 30322 48190 30324 48242
rect 30268 48188 30324 48190
rect 30716 48076 30772 48132
rect 28476 46956 28532 47012
rect 28476 45276 28532 45332
rect 29036 45276 29092 45332
rect 28364 44828 28420 44884
rect 28028 43538 28084 43540
rect 28028 43486 28030 43538
rect 28030 43486 28082 43538
rect 28082 43486 28084 43538
rect 28028 43484 28084 43486
rect 27356 41132 27412 41188
rect 26460 39394 26516 39396
rect 26460 39342 26462 39394
rect 26462 39342 26514 39394
rect 26514 39342 26516 39394
rect 26460 39340 26516 39342
rect 25676 38050 25732 38052
rect 25676 37998 25678 38050
rect 25678 37998 25730 38050
rect 25730 37998 25732 38050
rect 25676 37996 25732 37998
rect 25900 37826 25956 37828
rect 25900 37774 25902 37826
rect 25902 37774 25954 37826
rect 25954 37774 25956 37826
rect 25900 37772 25956 37774
rect 25228 37548 25284 37604
rect 25788 37660 25844 37716
rect 26348 37996 26404 38052
rect 26684 38220 26740 38276
rect 26348 37660 26404 37716
rect 26124 37548 26180 37604
rect 26460 37548 26516 37604
rect 25340 36652 25396 36708
rect 26012 36876 26068 36932
rect 26460 36428 26516 36484
rect 24108 35810 24164 35812
rect 24108 35758 24110 35810
rect 24110 35758 24162 35810
rect 24162 35758 24164 35810
rect 24108 35756 24164 35758
rect 23884 34860 23940 34916
rect 22652 31836 22708 31892
rect 22540 31778 22596 31780
rect 22540 31726 22542 31778
rect 22542 31726 22594 31778
rect 22594 31726 22596 31778
rect 22540 31724 22596 31726
rect 23212 34412 23268 34468
rect 24108 33346 24164 33348
rect 24108 33294 24110 33346
rect 24110 33294 24162 33346
rect 24162 33294 24164 33346
rect 24108 33292 24164 33294
rect 24556 35644 24612 35700
rect 25452 35756 25508 35812
rect 24892 35308 24948 35364
rect 24556 34690 24612 34692
rect 24556 34638 24558 34690
rect 24558 34638 24610 34690
rect 24610 34638 24612 34690
rect 24556 34636 24612 34638
rect 24332 33458 24388 33460
rect 24332 33406 24334 33458
rect 24334 33406 24386 33458
rect 24386 33406 24388 33458
rect 24332 33404 24388 33406
rect 23660 31890 23716 31892
rect 23660 31838 23662 31890
rect 23662 31838 23714 31890
rect 23714 31838 23716 31890
rect 23660 31836 23716 31838
rect 23212 31724 23268 31780
rect 23884 31500 23940 31556
rect 22204 26460 22260 26516
rect 21308 25394 21364 25396
rect 21308 25342 21310 25394
rect 21310 25342 21362 25394
rect 21362 25342 21364 25394
rect 21308 25340 21364 25342
rect 20188 23884 20244 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20188 23324 20244 23380
rect 18956 23100 19012 23156
rect 19740 23100 19796 23156
rect 18172 22204 18228 22260
rect 17724 21756 17780 21812
rect 18284 22316 18340 22372
rect 19516 22204 19572 22260
rect 18284 21196 18340 21252
rect 18396 22092 18452 22148
rect 18172 20860 18228 20916
rect 18060 20188 18116 20244
rect 16828 19292 16884 19348
rect 17052 19404 17108 19460
rect 17052 18396 17108 18452
rect 16044 17890 16100 17892
rect 16044 17838 16046 17890
rect 16046 17838 16098 17890
rect 16098 17838 16100 17890
rect 16044 17836 16100 17838
rect 16604 17948 16660 18004
rect 16604 17724 16660 17780
rect 16716 17836 16772 17892
rect 15484 17388 15540 17444
rect 15372 17106 15428 17108
rect 15372 17054 15374 17106
rect 15374 17054 15426 17106
rect 15426 17054 15428 17106
rect 15372 17052 15428 17054
rect 16156 17666 16212 17668
rect 16156 17614 16158 17666
rect 16158 17614 16210 17666
rect 16210 17614 16212 17666
rect 16156 17612 16212 17614
rect 17052 17724 17108 17780
rect 16156 17442 16212 17444
rect 16156 17390 16158 17442
rect 16158 17390 16210 17442
rect 16210 17390 16212 17442
rect 16156 17388 16212 17390
rect 16044 16994 16100 16996
rect 16044 16942 16046 16994
rect 16046 16942 16098 16994
rect 16098 16942 16100 16994
rect 16044 16940 16100 16942
rect 16716 16940 16772 16996
rect 16604 16828 16660 16884
rect 15372 16044 15428 16100
rect 14364 15260 14420 15316
rect 13132 15036 13188 15092
rect 14364 14306 14420 14308
rect 14364 14254 14366 14306
rect 14366 14254 14418 14306
rect 14418 14254 14420 14306
rect 14364 14252 14420 14254
rect 14924 15314 14980 15316
rect 14924 15262 14926 15314
rect 14926 15262 14978 15314
rect 14978 15262 14980 15314
rect 14924 15260 14980 15262
rect 15260 15484 15316 15540
rect 16156 16658 16212 16660
rect 16156 16606 16158 16658
rect 16158 16606 16210 16658
rect 16210 16606 16212 16658
rect 16156 16604 16212 16606
rect 16268 16156 16324 16212
rect 15596 15484 15652 15540
rect 15820 15708 15876 15764
rect 14700 14588 14756 14644
rect 15036 13634 15092 13636
rect 15036 13582 15038 13634
rect 15038 13582 15090 13634
rect 15090 13582 15092 13634
rect 15036 13580 15092 13582
rect 14252 13244 14308 13300
rect 14140 12684 14196 12740
rect 16044 15148 16100 15204
rect 16492 15484 16548 15540
rect 16716 16380 16772 16436
rect 15260 13858 15316 13860
rect 15260 13806 15262 13858
rect 15262 13806 15314 13858
rect 15314 13806 15316 13858
rect 15260 13804 15316 13806
rect 15260 13468 15316 13524
rect 14364 13074 14420 13076
rect 14364 13022 14366 13074
rect 14366 13022 14418 13074
rect 14418 13022 14420 13074
rect 14364 13020 14420 13022
rect 14812 13074 14868 13076
rect 14812 13022 14814 13074
rect 14814 13022 14866 13074
rect 14866 13022 14868 13074
rect 14812 13020 14868 13022
rect 14364 11900 14420 11956
rect 14140 11788 14196 11844
rect 14700 12012 14756 12068
rect 12908 11452 12964 11508
rect 13916 11506 13972 11508
rect 13916 11454 13918 11506
rect 13918 11454 13970 11506
rect 13970 11454 13972 11506
rect 13916 11452 13972 11454
rect 14252 11394 14308 11396
rect 14252 11342 14254 11394
rect 14254 11342 14306 11394
rect 14306 11342 14308 11394
rect 14252 11340 14308 11342
rect 14700 11506 14756 11508
rect 14700 11454 14702 11506
rect 14702 11454 14754 11506
rect 14754 11454 14756 11506
rect 14700 11452 14756 11454
rect 14140 10780 14196 10836
rect 13132 10444 13188 10500
rect 12908 10386 12964 10388
rect 12908 10334 12910 10386
rect 12910 10334 12962 10386
rect 12962 10334 12964 10386
rect 12908 10332 12964 10334
rect 13580 10332 13636 10388
rect 13132 10220 13188 10276
rect 12684 9938 12740 9940
rect 12684 9886 12686 9938
rect 12686 9886 12738 9938
rect 12738 9886 12740 9938
rect 12684 9884 12740 9886
rect 12572 9772 12628 9828
rect 12236 8092 12292 8148
rect 12572 8146 12628 8148
rect 12572 8094 12574 8146
rect 12574 8094 12626 8146
rect 12626 8094 12628 8146
rect 12572 8092 12628 8094
rect 12796 7868 12852 7924
rect 12908 8540 12964 8596
rect 12124 7196 12180 7252
rect 12460 6972 12516 7028
rect 12572 7196 12628 7252
rect 13580 9826 13636 9828
rect 13580 9774 13582 9826
rect 13582 9774 13634 9826
rect 13634 9774 13636 9826
rect 13580 9772 13636 9774
rect 13468 9548 13524 9604
rect 15036 12348 15092 12404
rect 15148 12572 15204 12628
rect 15036 11564 15092 11620
rect 14812 10780 14868 10836
rect 14924 11004 14980 11060
rect 13692 8370 13748 8372
rect 13692 8318 13694 8370
rect 13694 8318 13746 8370
rect 13746 8318 13748 8370
rect 13692 8316 13748 8318
rect 13580 7756 13636 7812
rect 12684 6972 12740 7028
rect 12236 6466 12292 6468
rect 12236 6414 12238 6466
rect 12238 6414 12290 6466
rect 12290 6414 12292 6466
rect 12236 6412 12292 6414
rect 12348 5346 12404 5348
rect 12348 5294 12350 5346
rect 12350 5294 12402 5346
rect 12402 5294 12404 5346
rect 12348 5292 12404 5294
rect 12908 5122 12964 5124
rect 12908 5070 12910 5122
rect 12910 5070 12962 5122
rect 12962 5070 12964 5122
rect 12908 5068 12964 5070
rect 11900 4956 11956 5012
rect 11228 4284 11284 4340
rect 11116 3836 11172 3892
rect 13468 4844 13524 4900
rect 13580 4956 13636 5012
rect 14812 8316 14868 8372
rect 15484 13634 15540 13636
rect 15484 13582 15486 13634
rect 15486 13582 15538 13634
rect 15538 13582 15540 13634
rect 15484 13580 15540 13582
rect 16044 14252 16100 14308
rect 15708 13970 15764 13972
rect 15708 13918 15710 13970
rect 15710 13918 15762 13970
rect 15762 13918 15764 13970
rect 15708 13916 15764 13918
rect 15708 13522 15764 13524
rect 15708 13470 15710 13522
rect 15710 13470 15762 13522
rect 15762 13470 15764 13522
rect 15708 13468 15764 13470
rect 16604 14306 16660 14308
rect 16604 14254 16606 14306
rect 16606 14254 16658 14306
rect 16658 14254 16660 14306
rect 16604 14252 16660 14254
rect 17276 19346 17332 19348
rect 17276 19294 17278 19346
rect 17278 19294 17330 19346
rect 17330 19294 17332 19346
rect 17276 19292 17332 19294
rect 19068 21698 19124 21700
rect 19068 21646 19070 21698
rect 19070 21646 19122 21698
rect 19122 21646 19124 21698
rect 19068 21644 19124 21646
rect 18508 21474 18564 21476
rect 18508 21422 18510 21474
rect 18510 21422 18562 21474
rect 18562 21422 18564 21474
rect 18508 21420 18564 21422
rect 20412 23548 20468 23604
rect 21532 25282 21588 25284
rect 21532 25230 21534 25282
rect 21534 25230 21586 25282
rect 21586 25230 21588 25282
rect 21532 25228 21588 25230
rect 20636 23212 20692 23268
rect 21532 25004 21588 25060
rect 20860 23884 20916 23940
rect 22204 25564 22260 25620
rect 22876 30268 22932 30324
rect 22428 29820 22484 29876
rect 22428 29596 22484 29652
rect 22652 28700 22708 28756
rect 22428 28082 22484 28084
rect 22428 28030 22430 28082
rect 22430 28030 22482 28082
rect 22482 28030 22484 28082
rect 22428 28028 22484 28030
rect 22540 27244 22596 27300
rect 22428 25506 22484 25508
rect 22428 25454 22430 25506
rect 22430 25454 22482 25506
rect 22482 25454 22484 25506
rect 22428 25452 22484 25454
rect 22204 25228 22260 25284
rect 21644 23884 21700 23940
rect 21756 25004 21812 25060
rect 20860 22204 20916 22260
rect 21308 22428 21364 22484
rect 20636 22092 20692 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20300 21644 20356 21700
rect 20524 21474 20580 21476
rect 20524 21422 20526 21474
rect 20526 21422 20578 21474
rect 20578 21422 20580 21474
rect 20524 21420 20580 21422
rect 21084 21698 21140 21700
rect 21084 21646 21086 21698
rect 21086 21646 21138 21698
rect 21138 21646 21140 21698
rect 21084 21644 21140 21646
rect 19516 20914 19572 20916
rect 19516 20862 19518 20914
rect 19518 20862 19570 20914
rect 19570 20862 19572 20914
rect 19516 20860 19572 20862
rect 18396 20748 18452 20804
rect 18396 20524 18452 20580
rect 18284 19292 18340 19348
rect 17836 19068 17892 19124
rect 17388 17666 17444 17668
rect 17388 17614 17390 17666
rect 17390 17614 17442 17666
rect 17442 17614 17444 17666
rect 17388 17612 17444 17614
rect 17500 17276 17556 17332
rect 17612 17164 17668 17220
rect 17612 16492 17668 16548
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20412 20188 20468 20244
rect 18396 18060 18452 18116
rect 18284 17612 18340 17668
rect 18060 16940 18116 16996
rect 17836 16882 17892 16884
rect 17836 16830 17838 16882
rect 17838 16830 17890 16882
rect 17890 16830 17892 16882
rect 17836 16828 17892 16830
rect 17724 16268 17780 16324
rect 17612 16098 17668 16100
rect 17612 16046 17614 16098
rect 17614 16046 17666 16098
rect 17666 16046 17668 16098
rect 17612 16044 17668 16046
rect 17948 15986 18004 15988
rect 17948 15934 17950 15986
rect 17950 15934 18002 15986
rect 18002 15934 18004 15986
rect 17948 15932 18004 15934
rect 18284 17106 18340 17108
rect 18284 17054 18286 17106
rect 18286 17054 18338 17106
rect 18338 17054 18340 17106
rect 18284 17052 18340 17054
rect 18284 16882 18340 16884
rect 18284 16830 18286 16882
rect 18286 16830 18338 16882
rect 18338 16830 18340 16882
rect 18284 16828 18340 16830
rect 18732 17276 18788 17332
rect 19964 19068 20020 19124
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 18956 17890 19012 17892
rect 18956 17838 18958 17890
rect 18958 17838 19010 17890
rect 19010 17838 19012 17890
rect 18956 17836 19012 17838
rect 19180 17778 19236 17780
rect 19180 17726 19182 17778
rect 19182 17726 19234 17778
rect 19234 17726 19236 17778
rect 19180 17724 19236 17726
rect 19628 18450 19684 18452
rect 19628 18398 19630 18450
rect 19630 18398 19682 18450
rect 19682 18398 19684 18450
rect 19628 18396 19684 18398
rect 21868 24892 21924 24948
rect 23548 30492 23604 30548
rect 24108 30492 24164 30548
rect 24556 33570 24612 33572
rect 24556 33518 24558 33570
rect 24558 33518 24610 33570
rect 24610 33518 24612 33570
rect 24556 33516 24612 33518
rect 25452 35196 25508 35252
rect 25004 34972 25060 35028
rect 25116 34914 25172 34916
rect 25116 34862 25118 34914
rect 25118 34862 25170 34914
rect 25170 34862 25172 34914
rect 25116 34860 25172 34862
rect 25676 34860 25732 34916
rect 25900 34972 25956 35028
rect 25452 34802 25508 34804
rect 25452 34750 25454 34802
rect 25454 34750 25506 34802
rect 25506 34750 25508 34802
rect 25452 34748 25508 34750
rect 25788 34690 25844 34692
rect 25788 34638 25790 34690
rect 25790 34638 25842 34690
rect 25842 34638 25844 34690
rect 25788 34636 25844 34638
rect 25452 34188 25508 34244
rect 24892 33068 24948 33124
rect 24668 31218 24724 31220
rect 24668 31166 24670 31218
rect 24670 31166 24722 31218
rect 24722 31166 24724 31218
rect 24668 31164 24724 31166
rect 23212 30156 23268 30212
rect 23212 29650 23268 29652
rect 23212 29598 23214 29650
rect 23214 29598 23266 29650
rect 23266 29598 23268 29650
rect 23212 29596 23268 29598
rect 23436 29036 23492 29092
rect 23548 28812 23604 28868
rect 23212 27244 23268 27300
rect 22540 23660 22596 23716
rect 22204 23324 22260 23380
rect 21980 22370 22036 22372
rect 21980 22318 21982 22370
rect 21982 22318 22034 22370
rect 22034 22318 22036 22370
rect 21980 22316 22036 22318
rect 22540 21980 22596 22036
rect 22204 21698 22260 21700
rect 22204 21646 22206 21698
rect 22206 21646 22258 21698
rect 22258 21646 22260 21698
rect 22204 21644 22260 21646
rect 23100 25618 23156 25620
rect 23100 25566 23102 25618
rect 23102 25566 23154 25618
rect 23154 25566 23156 25618
rect 23100 25564 23156 25566
rect 22988 25394 23044 25396
rect 22988 25342 22990 25394
rect 22990 25342 23042 25394
rect 23042 25342 23044 25394
rect 22988 25340 23044 25342
rect 23660 28642 23716 28644
rect 23660 28590 23662 28642
rect 23662 28590 23714 28642
rect 23714 28590 23716 28642
rect 23660 28588 23716 28590
rect 23884 29596 23940 29652
rect 23884 28364 23940 28420
rect 23660 28028 23716 28084
rect 24444 30716 24500 30772
rect 24892 30268 24948 30324
rect 25340 33346 25396 33348
rect 25340 33294 25342 33346
rect 25342 33294 25394 33346
rect 25394 33294 25396 33346
rect 25340 33292 25396 33294
rect 25004 30156 25060 30212
rect 25452 31554 25508 31556
rect 25452 31502 25454 31554
rect 25454 31502 25506 31554
rect 25506 31502 25508 31554
rect 25452 31500 25508 31502
rect 25228 31052 25284 31108
rect 25452 31164 25508 31220
rect 25900 34300 25956 34356
rect 25900 33964 25956 34020
rect 25116 30716 25172 30772
rect 24556 29932 24612 29988
rect 24220 29202 24276 29204
rect 24220 29150 24222 29202
rect 24222 29150 24274 29202
rect 24274 29150 24276 29202
rect 24220 29148 24276 29150
rect 24108 28530 24164 28532
rect 24108 28478 24110 28530
rect 24110 28478 24162 28530
rect 24162 28478 24164 28530
rect 24108 28476 24164 28478
rect 24108 28082 24164 28084
rect 24108 28030 24110 28082
rect 24110 28030 24162 28082
rect 24162 28030 24164 28082
rect 24108 28028 24164 28030
rect 25004 28642 25060 28644
rect 25004 28590 25006 28642
rect 25006 28590 25058 28642
rect 25058 28590 25060 28642
rect 25004 28588 25060 28590
rect 25676 30604 25732 30660
rect 25228 29426 25284 29428
rect 25228 29374 25230 29426
rect 25230 29374 25282 29426
rect 25282 29374 25284 29426
rect 25228 29372 25284 29374
rect 25228 29202 25284 29204
rect 25228 29150 25230 29202
rect 25230 29150 25282 29202
rect 25282 29150 25284 29202
rect 25228 29148 25284 29150
rect 25564 29202 25620 29204
rect 25564 29150 25566 29202
rect 25566 29150 25618 29202
rect 25618 29150 25620 29202
rect 25564 29148 25620 29150
rect 24332 28028 24388 28084
rect 24668 28364 24724 28420
rect 24444 27298 24500 27300
rect 24444 27246 24446 27298
rect 24446 27246 24498 27298
rect 24498 27246 24500 27298
rect 24444 27244 24500 27246
rect 23772 25452 23828 25508
rect 23996 25340 24052 25396
rect 24556 25676 24612 25732
rect 24444 25394 24500 25396
rect 24444 25342 24446 25394
rect 24446 25342 24498 25394
rect 24498 25342 24500 25394
rect 24444 25340 24500 25342
rect 24220 24834 24276 24836
rect 24220 24782 24222 24834
rect 24222 24782 24274 24834
rect 24274 24782 24276 24834
rect 24220 24780 24276 24782
rect 23100 23378 23156 23380
rect 23100 23326 23102 23378
rect 23102 23326 23154 23378
rect 23154 23326 23156 23378
rect 23100 23324 23156 23326
rect 22988 21980 23044 22036
rect 22876 21308 22932 21364
rect 23324 23938 23380 23940
rect 23324 23886 23326 23938
rect 23326 23886 23378 23938
rect 23378 23886 23380 23938
rect 23324 23884 23380 23886
rect 25564 28700 25620 28756
rect 25452 28476 25508 28532
rect 25676 27244 25732 27300
rect 25228 26012 25284 26068
rect 25564 25900 25620 25956
rect 26572 36370 26628 36372
rect 26572 36318 26574 36370
rect 26574 36318 26626 36370
rect 26626 36318 26628 36370
rect 26572 36316 26628 36318
rect 26460 35868 26516 35924
rect 27804 41132 27860 41188
rect 28700 43538 28756 43540
rect 28700 43486 28702 43538
rect 28702 43486 28754 43538
rect 28754 43486 28756 43538
rect 28700 43484 28756 43486
rect 29260 44828 29316 44884
rect 32172 48300 32228 48356
rect 30828 47964 30884 48020
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 32284 47404 32340 47460
rect 34076 48188 34132 48244
rect 35756 48188 35812 48244
rect 33740 48076 33796 48132
rect 30716 46956 30772 47012
rect 33068 47458 33124 47460
rect 33068 47406 33070 47458
rect 33070 47406 33122 47458
rect 33122 47406 33124 47458
rect 33068 47404 33124 47406
rect 32620 47180 32676 47236
rect 30156 46732 30212 46788
rect 31948 46786 32004 46788
rect 31948 46734 31950 46786
rect 31950 46734 32002 46786
rect 32002 46734 32004 46786
rect 31948 46732 32004 46734
rect 32396 46786 32452 46788
rect 32396 46734 32398 46786
rect 32398 46734 32450 46786
rect 32450 46734 32452 46786
rect 32396 46732 32452 46734
rect 33404 46732 33460 46788
rect 33516 47180 33572 47236
rect 29932 45330 29988 45332
rect 29932 45278 29934 45330
rect 29934 45278 29986 45330
rect 29986 45278 29988 45330
rect 29932 45276 29988 45278
rect 30268 45164 30324 45220
rect 30156 45052 30212 45108
rect 30604 45164 30660 45220
rect 30268 44940 30324 44996
rect 30716 44828 30772 44884
rect 30716 44268 30772 44324
rect 30604 43708 30660 43764
rect 29820 43260 29876 43316
rect 30044 41804 30100 41860
rect 29596 41186 29652 41188
rect 29596 41134 29598 41186
rect 29598 41134 29650 41186
rect 29650 41134 29652 41186
rect 29596 41132 29652 41134
rect 27468 39394 27524 39396
rect 27468 39342 27470 39394
rect 27470 39342 27522 39394
rect 27522 39342 27524 39394
rect 27468 39340 27524 39342
rect 27804 38668 27860 38724
rect 27468 38332 27524 38388
rect 27020 37266 27076 37268
rect 27020 37214 27022 37266
rect 27022 37214 27074 37266
rect 27074 37214 27076 37266
rect 27020 37212 27076 37214
rect 27692 38050 27748 38052
rect 27692 37998 27694 38050
rect 27694 37998 27746 38050
rect 27746 37998 27748 38050
rect 27692 37996 27748 37998
rect 27468 37212 27524 37268
rect 27580 37436 27636 37492
rect 27356 36988 27412 37044
rect 26908 36540 26964 36596
rect 27020 36876 27076 36932
rect 26124 35196 26180 35252
rect 26684 35586 26740 35588
rect 26684 35534 26686 35586
rect 26686 35534 26738 35586
rect 26738 35534 26740 35586
rect 26684 35532 26740 35534
rect 26684 35196 26740 35252
rect 26908 34860 26964 34916
rect 26236 34018 26292 34020
rect 26236 33966 26238 34018
rect 26238 33966 26290 34018
rect 26290 33966 26292 34018
rect 26236 33964 26292 33966
rect 26236 32562 26292 32564
rect 26236 32510 26238 32562
rect 26238 32510 26290 32562
rect 26290 32510 26292 32562
rect 26236 32508 26292 32510
rect 26460 31106 26516 31108
rect 26460 31054 26462 31106
rect 26462 31054 26514 31106
rect 26514 31054 26516 31106
rect 26460 31052 26516 31054
rect 26684 34188 26740 34244
rect 27580 36988 27636 37044
rect 27468 35586 27524 35588
rect 27468 35534 27470 35586
rect 27470 35534 27522 35586
rect 27522 35534 27524 35586
rect 27468 35532 27524 35534
rect 27468 35196 27524 35252
rect 27468 34914 27524 34916
rect 27468 34862 27470 34914
rect 27470 34862 27522 34914
rect 27522 34862 27524 34914
rect 27468 34860 27524 34862
rect 26908 34300 26964 34356
rect 27132 33404 27188 33460
rect 26236 29986 26292 29988
rect 26236 29934 26238 29986
rect 26238 29934 26290 29986
rect 26290 29934 26292 29986
rect 26236 29932 26292 29934
rect 26012 29426 26068 29428
rect 26012 29374 26014 29426
rect 26014 29374 26066 29426
rect 26066 29374 26068 29426
rect 26012 29372 26068 29374
rect 26012 28812 26068 28868
rect 26124 27746 26180 27748
rect 26124 27694 26126 27746
rect 26126 27694 26178 27746
rect 26178 27694 26180 27746
rect 26124 27692 26180 27694
rect 25004 24668 25060 24724
rect 23324 23548 23380 23604
rect 21756 20524 21812 20580
rect 21532 20300 21588 20356
rect 22428 20300 22484 20356
rect 20972 19906 21028 19908
rect 20972 19854 20974 19906
rect 20974 19854 21026 19906
rect 21026 19854 21028 19906
rect 20972 19852 21028 19854
rect 22652 19964 22708 20020
rect 22764 20524 22820 20580
rect 21980 19852 22036 19908
rect 20860 18060 20916 18116
rect 19292 17612 19348 17668
rect 20076 17388 20132 17444
rect 19628 17276 19684 17332
rect 19068 17106 19124 17108
rect 19068 17054 19070 17106
rect 19070 17054 19122 17106
rect 19122 17054 19124 17106
rect 19068 17052 19124 17054
rect 18508 16604 18564 16660
rect 18620 16380 18676 16436
rect 19068 16828 19124 16884
rect 17164 14924 17220 14980
rect 17276 14588 17332 14644
rect 17164 14530 17220 14532
rect 17164 14478 17166 14530
rect 17166 14478 17218 14530
rect 17218 14478 17220 14530
rect 17164 14476 17220 14478
rect 17724 14530 17780 14532
rect 17724 14478 17726 14530
rect 17726 14478 17778 14530
rect 17778 14478 17780 14530
rect 17724 14476 17780 14478
rect 17052 14418 17108 14420
rect 17052 14366 17054 14418
rect 17054 14366 17106 14418
rect 17106 14366 17108 14418
rect 17052 14364 17108 14366
rect 17388 14364 17444 14420
rect 16268 13804 16324 13860
rect 16044 13244 16100 13300
rect 16156 13746 16212 13748
rect 16156 13694 16158 13746
rect 16158 13694 16210 13746
rect 16210 13694 16212 13746
rect 16156 13692 16212 13694
rect 16380 13074 16436 13076
rect 16380 13022 16382 13074
rect 16382 13022 16434 13074
rect 16434 13022 16436 13074
rect 16380 13020 16436 13022
rect 15820 12908 15876 12964
rect 15932 12850 15988 12852
rect 15932 12798 15934 12850
rect 15934 12798 15986 12850
rect 15986 12798 15988 12850
rect 15932 12796 15988 12798
rect 15932 12460 15988 12516
rect 17612 13746 17668 13748
rect 17612 13694 17614 13746
rect 17614 13694 17666 13746
rect 17666 13694 17668 13746
rect 17612 13692 17668 13694
rect 17500 13634 17556 13636
rect 17500 13582 17502 13634
rect 17502 13582 17554 13634
rect 17554 13582 17556 13634
rect 17500 13580 17556 13582
rect 17836 13468 17892 13524
rect 16940 12962 16996 12964
rect 16940 12910 16942 12962
rect 16942 12910 16994 12962
rect 16994 12910 16996 12962
rect 16940 12908 16996 12910
rect 17388 12962 17444 12964
rect 17388 12910 17390 12962
rect 17390 12910 17442 12962
rect 17442 12910 17444 12962
rect 17388 12908 17444 12910
rect 16492 12850 16548 12852
rect 16492 12798 16494 12850
rect 16494 12798 16546 12850
rect 16546 12798 16548 12850
rect 16492 12796 16548 12798
rect 16156 12738 16212 12740
rect 16156 12686 16158 12738
rect 16158 12686 16210 12738
rect 16210 12686 16212 12738
rect 16156 12684 16212 12686
rect 16268 12290 16324 12292
rect 16268 12238 16270 12290
rect 16270 12238 16322 12290
rect 16322 12238 16324 12290
rect 16268 12236 16324 12238
rect 15596 12066 15652 12068
rect 15596 12014 15598 12066
rect 15598 12014 15650 12066
rect 15650 12014 15652 12066
rect 15596 12012 15652 12014
rect 15372 11618 15428 11620
rect 15372 11566 15374 11618
rect 15374 11566 15426 11618
rect 15426 11566 15428 11618
rect 15372 11564 15428 11566
rect 16044 11676 16100 11732
rect 15260 11004 15316 11060
rect 15260 10834 15316 10836
rect 15260 10782 15262 10834
rect 15262 10782 15314 10834
rect 15314 10782 15316 10834
rect 15260 10780 15316 10782
rect 16156 10780 16212 10836
rect 15820 10332 15876 10388
rect 16268 9996 16324 10052
rect 15260 9602 15316 9604
rect 15260 9550 15262 9602
rect 15262 9550 15314 9602
rect 15314 9550 15316 9602
rect 15260 9548 15316 9550
rect 14924 9436 14980 9492
rect 14588 8204 14644 8260
rect 14028 7756 14084 7812
rect 13916 7474 13972 7476
rect 13916 7422 13918 7474
rect 13918 7422 13970 7474
rect 13970 7422 13972 7474
rect 13916 7420 13972 7422
rect 16044 9436 16100 9492
rect 16268 9212 16324 9268
rect 16492 12460 16548 12516
rect 17836 12796 17892 12852
rect 17724 12402 17780 12404
rect 17724 12350 17726 12402
rect 17726 12350 17778 12402
rect 17778 12350 17780 12402
rect 17724 12348 17780 12350
rect 17948 12012 18004 12068
rect 16604 9548 16660 9604
rect 15372 8930 15428 8932
rect 15372 8878 15374 8930
rect 15374 8878 15426 8930
rect 15426 8878 15428 8930
rect 15372 8876 15428 8878
rect 15484 8316 15540 8372
rect 15260 8146 15316 8148
rect 15260 8094 15262 8146
rect 15262 8094 15314 8146
rect 15314 8094 15316 8146
rect 15260 8092 15316 8094
rect 14924 7084 14980 7140
rect 14588 6748 14644 6804
rect 14140 6636 14196 6692
rect 14476 6578 14532 6580
rect 14476 6526 14478 6578
rect 14478 6526 14530 6578
rect 14530 6526 14532 6578
rect 14476 6524 14532 6526
rect 16492 8482 16548 8484
rect 16492 8430 16494 8482
rect 16494 8430 16546 8482
rect 16546 8430 16548 8482
rect 16492 8428 16548 8430
rect 16044 8316 16100 8372
rect 16380 8316 16436 8372
rect 16492 7980 16548 8036
rect 16380 7698 16436 7700
rect 16380 7646 16382 7698
rect 16382 7646 16434 7698
rect 16434 7646 16436 7698
rect 16380 7644 16436 7646
rect 16044 7308 16100 7364
rect 15820 7196 15876 7252
rect 15372 7084 15428 7140
rect 15484 6914 15540 6916
rect 15484 6862 15486 6914
rect 15486 6862 15538 6914
rect 15538 6862 15540 6914
rect 15484 6860 15540 6862
rect 15036 6524 15092 6580
rect 15148 6300 15204 6356
rect 15036 6018 15092 6020
rect 15036 5966 15038 6018
rect 15038 5966 15090 6018
rect 15090 5966 15092 6018
rect 15036 5964 15092 5966
rect 14364 5794 14420 5796
rect 14364 5742 14366 5794
rect 14366 5742 14418 5794
rect 14418 5742 14420 5794
rect 14364 5740 14420 5742
rect 14812 5180 14868 5236
rect 14364 5068 14420 5124
rect 14140 3724 14196 3780
rect 13244 3612 13300 3668
rect 12460 3442 12516 3444
rect 12460 3390 12462 3442
rect 12462 3390 12514 3442
rect 12514 3390 12516 3442
rect 12460 3388 12516 3390
rect 7756 2940 7812 2996
rect 14476 3948 14532 4004
rect 15484 5740 15540 5796
rect 15596 5516 15652 5572
rect 16268 5404 16324 5460
rect 16380 5068 16436 5124
rect 16828 8930 16884 8932
rect 16828 8878 16830 8930
rect 16830 8878 16882 8930
rect 16882 8878 16884 8930
rect 16828 8876 16884 8878
rect 16716 7698 16772 7700
rect 16716 7646 16718 7698
rect 16718 7646 16770 7698
rect 16770 7646 16772 7698
rect 16716 7644 16772 7646
rect 16716 7084 16772 7140
rect 17500 9714 17556 9716
rect 17500 9662 17502 9714
rect 17502 9662 17554 9714
rect 17554 9662 17556 9714
rect 17500 9660 17556 9662
rect 18060 11452 18116 11508
rect 17836 11394 17892 11396
rect 17836 11342 17838 11394
rect 17838 11342 17890 11394
rect 17890 11342 17892 11394
rect 17836 11340 17892 11342
rect 18956 15986 19012 15988
rect 18956 15934 18958 15986
rect 18958 15934 19010 15986
rect 19010 15934 19012 15986
rect 18956 15932 19012 15934
rect 19292 16716 19348 16772
rect 19516 16380 19572 16436
rect 18620 12572 18676 12628
rect 18620 12012 18676 12068
rect 18172 9996 18228 10052
rect 17836 9660 17892 9716
rect 17164 9212 17220 9268
rect 17276 9042 17332 9044
rect 17276 8990 17278 9042
rect 17278 8990 17330 9042
rect 17330 8990 17332 9042
rect 17276 8988 17332 8990
rect 18172 9436 18228 9492
rect 18284 9324 18340 9380
rect 17612 9266 17668 9268
rect 17612 9214 17614 9266
rect 17614 9214 17666 9266
rect 17666 9214 17668 9266
rect 17612 9212 17668 9214
rect 17276 8428 17332 8484
rect 17052 7868 17108 7924
rect 17948 8764 18004 8820
rect 17724 7532 17780 7588
rect 18732 11340 18788 11396
rect 19180 13916 19236 13972
rect 19068 13468 19124 13524
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19852 17106 19908 17108
rect 19852 17054 19854 17106
rect 19854 17054 19906 17106
rect 19906 17054 19908 17106
rect 19852 17052 19908 17054
rect 20076 16770 20132 16772
rect 20076 16718 20078 16770
rect 20078 16718 20130 16770
rect 20130 16718 20132 16770
rect 20076 16716 20132 16718
rect 19628 15932 19684 15988
rect 20860 16716 20916 16772
rect 20412 16044 20468 16100
rect 20636 16604 20692 16660
rect 20188 15820 20244 15876
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19516 15484 19572 15540
rect 21308 16994 21364 16996
rect 21308 16942 21310 16994
rect 21310 16942 21362 16994
rect 21362 16942 21364 16994
rect 21308 16940 21364 16942
rect 24668 23660 24724 23716
rect 24220 22540 24276 22596
rect 23436 22482 23492 22484
rect 23436 22430 23438 22482
rect 23438 22430 23490 22482
rect 23490 22430 23492 22482
rect 23436 22428 23492 22430
rect 24332 23548 24388 23604
rect 23436 21980 23492 22036
rect 23772 21698 23828 21700
rect 23772 21646 23774 21698
rect 23774 21646 23826 21698
rect 23826 21646 23828 21698
rect 23772 21644 23828 21646
rect 25228 22764 25284 22820
rect 24668 21644 24724 21700
rect 25452 21698 25508 21700
rect 25452 21646 25454 21698
rect 25454 21646 25506 21698
rect 25506 21646 25508 21698
rect 25452 21644 25508 21646
rect 22988 20524 23044 20580
rect 23436 20412 23492 20468
rect 23660 20524 23716 20580
rect 23436 20018 23492 20020
rect 23436 19966 23438 20018
rect 23438 19966 23490 20018
rect 23490 19966 23492 20018
rect 23436 19964 23492 19966
rect 21868 19068 21924 19124
rect 21756 18396 21812 18452
rect 21532 17666 21588 17668
rect 21532 17614 21534 17666
rect 21534 17614 21586 17666
rect 21586 17614 21588 17666
rect 21532 17612 21588 17614
rect 21868 17554 21924 17556
rect 21868 17502 21870 17554
rect 21870 17502 21922 17554
rect 21922 17502 21924 17554
rect 21868 17500 21924 17502
rect 22092 17948 22148 18004
rect 22092 17554 22148 17556
rect 22092 17502 22094 17554
rect 22094 17502 22146 17554
rect 22146 17502 22148 17554
rect 22092 17500 22148 17502
rect 21756 16828 21812 16884
rect 21980 16940 22036 16996
rect 21644 16770 21700 16772
rect 21644 16718 21646 16770
rect 21646 16718 21698 16770
rect 21698 16718 21700 16770
rect 21644 16716 21700 16718
rect 21420 16380 21476 16436
rect 19740 15202 19796 15204
rect 19740 15150 19742 15202
rect 19742 15150 19794 15202
rect 19794 15150 19796 15202
rect 19740 15148 19796 15150
rect 21756 16044 21812 16100
rect 20972 15148 21028 15204
rect 19852 14700 19908 14756
rect 20076 14812 20132 14868
rect 20300 14530 20356 14532
rect 20300 14478 20302 14530
rect 20302 14478 20354 14530
rect 20354 14478 20356 14530
rect 20300 14476 20356 14478
rect 20636 14754 20692 14756
rect 20636 14702 20638 14754
rect 20638 14702 20690 14754
rect 20690 14702 20692 14754
rect 20636 14700 20692 14702
rect 20188 14252 20244 14308
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20860 14588 20916 14644
rect 18620 9212 18676 9268
rect 18956 11506 19012 11508
rect 18956 11454 18958 11506
rect 18958 11454 19010 11506
rect 19010 11454 19012 11506
rect 18956 11452 19012 11454
rect 18956 11116 19012 11172
rect 18396 8988 18452 9044
rect 19068 11340 19124 11396
rect 18956 10834 19012 10836
rect 18956 10782 18958 10834
rect 18958 10782 19010 10834
rect 19010 10782 19012 10834
rect 18956 10780 19012 10782
rect 19068 10556 19124 10612
rect 18844 9884 18900 9940
rect 18844 9324 18900 9380
rect 19180 9996 19236 10052
rect 19516 10556 19572 10612
rect 20188 13468 20244 13524
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20748 13692 20804 13748
rect 20300 11900 20356 11956
rect 20748 11900 20804 11956
rect 20188 10892 20244 10948
rect 19740 10610 19796 10612
rect 19740 10558 19742 10610
rect 19742 10558 19794 10610
rect 19794 10558 19796 10610
rect 19740 10556 19796 10558
rect 21196 15484 21252 15540
rect 21420 15426 21476 15428
rect 21420 15374 21422 15426
rect 21422 15374 21474 15426
rect 21474 15374 21476 15426
rect 21420 15372 21476 15374
rect 21532 15148 21588 15204
rect 21308 14476 21364 14532
rect 21084 14252 21140 14308
rect 21980 15874 22036 15876
rect 21980 15822 21982 15874
rect 21982 15822 22034 15874
rect 22034 15822 22036 15874
rect 21980 15820 22036 15822
rect 21980 15314 22036 15316
rect 21980 15262 21982 15314
rect 21982 15262 22034 15314
rect 22034 15262 22036 15314
rect 21980 15260 22036 15262
rect 22204 16716 22260 16772
rect 22540 17164 22596 17220
rect 22428 16882 22484 16884
rect 22428 16830 22430 16882
rect 22430 16830 22482 16882
rect 22482 16830 22484 16882
rect 22428 16828 22484 16830
rect 22428 16380 22484 16436
rect 22204 15484 22260 15540
rect 21756 14588 21812 14644
rect 22204 15148 22260 15204
rect 22316 15260 22372 15316
rect 21308 13970 21364 13972
rect 21308 13918 21310 13970
rect 21310 13918 21362 13970
rect 21362 13918 21364 13970
rect 21308 13916 21364 13918
rect 21420 13746 21476 13748
rect 21420 13694 21422 13746
rect 21422 13694 21474 13746
rect 21474 13694 21476 13746
rect 21420 13692 21476 13694
rect 22540 14588 22596 14644
rect 22988 17836 23044 17892
rect 23884 20130 23940 20132
rect 23884 20078 23886 20130
rect 23886 20078 23938 20130
rect 23938 20078 23940 20130
rect 23884 20076 23940 20078
rect 23772 17948 23828 18004
rect 23772 16940 23828 16996
rect 22876 16716 22932 16772
rect 22988 16658 23044 16660
rect 22988 16606 22990 16658
rect 22990 16606 23042 16658
rect 23042 16606 23044 16658
rect 22988 16604 23044 16606
rect 22988 16156 23044 16212
rect 24780 20802 24836 20804
rect 24780 20750 24782 20802
rect 24782 20750 24834 20802
rect 24834 20750 24836 20802
rect 24780 20748 24836 20750
rect 24556 19794 24612 19796
rect 24556 19742 24558 19794
rect 24558 19742 24610 19794
rect 24610 19742 24612 19794
rect 24556 19740 24612 19742
rect 24444 18620 24500 18676
rect 25564 20636 25620 20692
rect 25116 20076 25172 20132
rect 25340 20130 25396 20132
rect 25340 20078 25342 20130
rect 25342 20078 25394 20130
rect 25394 20078 25396 20130
rect 25340 20076 25396 20078
rect 25004 18508 25060 18564
rect 24444 18172 24500 18228
rect 24108 17612 24164 17668
rect 25228 18396 25284 18452
rect 24780 18284 24836 18340
rect 24780 18060 24836 18116
rect 24556 17948 24612 18004
rect 24668 17612 24724 17668
rect 23996 16604 24052 16660
rect 23884 16380 23940 16436
rect 23548 15932 23604 15988
rect 23548 15314 23604 15316
rect 23548 15262 23550 15314
rect 23550 15262 23602 15314
rect 23602 15262 23604 15314
rect 23548 15260 23604 15262
rect 23212 14588 23268 14644
rect 22092 14306 22148 14308
rect 22092 14254 22094 14306
rect 22094 14254 22146 14306
rect 22146 14254 22148 14306
rect 22092 14252 22148 14254
rect 23548 14530 23604 14532
rect 23548 14478 23550 14530
rect 23550 14478 23602 14530
rect 23602 14478 23604 14530
rect 23548 14476 23604 14478
rect 25228 16994 25284 16996
rect 25228 16942 25230 16994
rect 25230 16942 25282 16994
rect 25282 16942 25284 16994
rect 25228 16940 25284 16942
rect 25564 19068 25620 19124
rect 25564 18674 25620 18676
rect 25564 18622 25566 18674
rect 25566 18622 25618 18674
rect 25618 18622 25620 18674
rect 25564 18620 25620 18622
rect 26012 27580 26068 27636
rect 26124 25228 26180 25284
rect 26236 25340 26292 25396
rect 26012 22876 26068 22932
rect 26572 27298 26628 27300
rect 26572 27246 26574 27298
rect 26574 27246 26626 27298
rect 26626 27246 26628 27298
rect 26572 27244 26628 27246
rect 27020 29820 27076 29876
rect 27692 37324 27748 37380
rect 27916 37826 27972 37828
rect 27916 37774 27918 37826
rect 27918 37774 27970 37826
rect 27970 37774 27972 37826
rect 27916 37772 27972 37774
rect 27916 37324 27972 37380
rect 27916 36370 27972 36372
rect 27916 36318 27918 36370
rect 27918 36318 27970 36370
rect 27970 36318 27972 36370
rect 27916 36316 27972 36318
rect 27692 35868 27748 35924
rect 27804 35308 27860 35364
rect 28700 38668 28756 38724
rect 29036 38946 29092 38948
rect 29036 38894 29038 38946
rect 29038 38894 29090 38946
rect 29090 38894 29092 38946
rect 29036 38892 29092 38894
rect 28252 36988 28308 37044
rect 28364 36876 28420 36932
rect 28140 35420 28196 35476
rect 27804 34188 27860 34244
rect 27804 34018 27860 34020
rect 27804 33966 27806 34018
rect 27806 33966 27858 34018
rect 27858 33966 27860 34018
rect 27804 33964 27860 33966
rect 28252 35084 28308 35140
rect 28028 34300 28084 34356
rect 28028 34130 28084 34132
rect 28028 34078 28030 34130
rect 28030 34078 28082 34130
rect 28082 34078 28084 34130
rect 28028 34076 28084 34078
rect 29596 40348 29652 40404
rect 28700 37212 28756 37268
rect 29484 38332 29540 38388
rect 28588 36258 28644 36260
rect 28588 36206 28590 36258
rect 28590 36206 28642 36258
rect 28642 36206 28644 36258
rect 28588 36204 28644 36206
rect 28588 35420 28644 35476
rect 29036 36764 29092 36820
rect 28924 36204 28980 36260
rect 29484 37212 29540 37268
rect 29148 35980 29204 36036
rect 30156 41580 30212 41636
rect 30492 40348 30548 40404
rect 30268 40124 30324 40180
rect 31612 44492 31668 44548
rect 33404 45052 33460 45108
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35532 47068 35588 47124
rect 33740 46956 33796 47012
rect 31948 44268 32004 44324
rect 32956 43708 33012 43764
rect 32508 43596 32564 43652
rect 32060 43538 32116 43540
rect 32060 43486 32062 43538
rect 32062 43486 32114 43538
rect 32114 43486 32116 43538
rect 32060 43484 32116 43486
rect 31500 43314 31556 43316
rect 31500 43262 31502 43314
rect 31502 43262 31554 43314
rect 31554 43262 31556 43314
rect 31500 43260 31556 43262
rect 30716 41858 30772 41860
rect 30716 41806 30718 41858
rect 30718 41806 30770 41858
rect 30770 41806 30772 41858
rect 30716 41804 30772 41806
rect 31052 41580 31108 41636
rect 34300 44156 34356 44212
rect 33404 43708 33460 43764
rect 33628 43596 33684 43652
rect 31724 40908 31780 40964
rect 31052 40178 31108 40180
rect 31052 40126 31054 40178
rect 31054 40126 31106 40178
rect 31106 40126 31108 40178
rect 31052 40124 31108 40126
rect 30268 38892 30324 38948
rect 29708 36764 29764 36820
rect 29820 36428 29876 36484
rect 29932 36988 29988 37044
rect 29372 36370 29428 36372
rect 29372 36318 29374 36370
rect 29374 36318 29426 36370
rect 29426 36318 29428 36370
rect 29372 36316 29428 36318
rect 29932 36370 29988 36372
rect 29932 36318 29934 36370
rect 29934 36318 29986 36370
rect 29986 36318 29988 36370
rect 29932 36316 29988 36318
rect 32508 40962 32564 40964
rect 32508 40910 32510 40962
rect 32510 40910 32562 40962
rect 32562 40910 32564 40962
rect 32508 40908 32564 40910
rect 31836 40348 31892 40404
rect 32508 40402 32564 40404
rect 32508 40350 32510 40402
rect 32510 40350 32562 40402
rect 32562 40350 32564 40402
rect 32508 40348 32564 40350
rect 31724 40236 31780 40292
rect 31948 40236 32004 40292
rect 31612 38834 31668 38836
rect 31612 38782 31614 38834
rect 31614 38782 31666 38834
rect 31666 38782 31668 38834
rect 31612 38780 31668 38782
rect 32284 38444 32340 38500
rect 30940 37772 30996 37828
rect 30828 36988 30884 37044
rect 31500 37100 31556 37156
rect 30492 36876 30548 36932
rect 30156 36428 30212 36484
rect 29036 35810 29092 35812
rect 29036 35758 29038 35810
rect 29038 35758 29090 35810
rect 29090 35758 29092 35810
rect 29036 35756 29092 35758
rect 29596 35420 29652 35476
rect 28700 35196 28756 35252
rect 29260 35084 29316 35140
rect 28700 34748 28756 34804
rect 28588 34412 28644 34468
rect 28140 33516 28196 33572
rect 28140 33122 28196 33124
rect 28140 33070 28142 33122
rect 28142 33070 28194 33122
rect 28194 33070 28196 33122
rect 28140 33068 28196 33070
rect 28812 34412 28868 34468
rect 28812 34188 28868 34244
rect 28476 33234 28532 33236
rect 28476 33182 28478 33234
rect 28478 33182 28530 33234
rect 28530 33182 28532 33234
rect 28476 33180 28532 33182
rect 27916 32620 27972 32676
rect 27916 31724 27972 31780
rect 27804 29820 27860 29876
rect 27468 29148 27524 29204
rect 27356 28140 27412 28196
rect 27020 28028 27076 28084
rect 27692 27916 27748 27972
rect 27468 27858 27524 27860
rect 27468 27806 27470 27858
rect 27470 27806 27522 27858
rect 27522 27806 27524 27858
rect 27468 27804 27524 27806
rect 27580 27692 27636 27748
rect 26572 25788 26628 25844
rect 26572 25506 26628 25508
rect 26572 25454 26574 25506
rect 26574 25454 26626 25506
rect 26626 25454 26628 25506
rect 26572 25452 26628 25454
rect 26348 25116 26404 25172
rect 25900 21026 25956 21028
rect 25900 20974 25902 21026
rect 25902 20974 25954 21026
rect 25954 20974 25956 21026
rect 25900 20972 25956 20974
rect 26348 24834 26404 24836
rect 26348 24782 26350 24834
rect 26350 24782 26402 24834
rect 26402 24782 26404 24834
rect 26348 24780 26404 24782
rect 26236 24444 26292 24500
rect 26460 22876 26516 22932
rect 26908 25618 26964 25620
rect 26908 25566 26910 25618
rect 26910 25566 26962 25618
rect 26962 25566 26964 25618
rect 26908 25564 26964 25566
rect 27132 25676 27188 25732
rect 26796 25116 26852 25172
rect 27020 25116 27076 25172
rect 26796 24892 26852 24948
rect 26796 24108 26852 24164
rect 27468 25116 27524 25172
rect 27580 25452 27636 25508
rect 27692 25282 27748 25284
rect 27692 25230 27694 25282
rect 27694 25230 27746 25282
rect 27746 25230 27748 25282
rect 27692 25228 27748 25230
rect 27580 24556 27636 24612
rect 27804 24444 27860 24500
rect 27468 24220 27524 24276
rect 27020 23884 27076 23940
rect 27356 24108 27412 24164
rect 26572 22428 26628 22484
rect 26796 21698 26852 21700
rect 26796 21646 26798 21698
rect 26798 21646 26850 21698
rect 26850 21646 26852 21698
rect 26796 21644 26852 21646
rect 26908 21644 26964 21700
rect 26460 21532 26516 21588
rect 26236 20972 26292 21028
rect 26124 20300 26180 20356
rect 25900 19852 25956 19908
rect 26236 20076 26292 20132
rect 25676 18396 25732 18452
rect 24668 16828 24724 16884
rect 22988 14364 23044 14420
rect 21196 13020 21252 13076
rect 21644 13074 21700 13076
rect 21644 13022 21646 13074
rect 21646 13022 21698 13074
rect 21698 13022 21700 13074
rect 21644 13020 21700 13022
rect 21084 11676 21140 11732
rect 21980 12290 22036 12292
rect 21980 12238 21982 12290
rect 21982 12238 22034 12290
rect 22034 12238 22036 12290
rect 21980 12236 22036 12238
rect 21756 11676 21812 11732
rect 22316 12290 22372 12292
rect 22316 12238 22318 12290
rect 22318 12238 22370 12290
rect 22370 12238 22372 12290
rect 22316 12236 22372 12238
rect 22092 12012 22148 12068
rect 22652 11900 22708 11956
rect 21868 11564 21924 11620
rect 20972 11004 21028 11060
rect 21196 11116 21252 11172
rect 20748 10892 20804 10948
rect 22316 11004 22372 11060
rect 19292 9714 19348 9716
rect 19292 9662 19294 9714
rect 19294 9662 19346 9714
rect 19346 9662 19348 9714
rect 19292 9660 19348 9662
rect 19404 9266 19460 9268
rect 19404 9214 19406 9266
rect 19406 9214 19458 9266
rect 19458 9214 19460 9266
rect 19404 9212 19460 9214
rect 18956 9100 19012 9156
rect 18284 8764 18340 8820
rect 18844 8876 18900 8932
rect 18508 8764 18564 8820
rect 18732 8370 18788 8372
rect 18732 8318 18734 8370
rect 18734 8318 18786 8370
rect 18786 8318 18788 8370
rect 18732 8316 18788 8318
rect 19180 9042 19236 9044
rect 19180 8990 19182 9042
rect 19182 8990 19234 9042
rect 19234 8990 19236 9042
rect 19180 8988 19236 8990
rect 19292 8764 19348 8820
rect 19516 8204 19572 8260
rect 18060 7868 18116 7924
rect 18284 7532 18340 7588
rect 17276 7308 17332 7364
rect 17164 6578 17220 6580
rect 17164 6526 17166 6578
rect 17166 6526 17218 6578
rect 17218 6526 17220 6578
rect 17164 6524 17220 6526
rect 16940 6076 16996 6132
rect 15372 3836 15428 3892
rect 16828 3778 16884 3780
rect 16828 3726 16830 3778
rect 16830 3726 16882 3778
rect 16882 3726 16884 3778
rect 16828 3724 16884 3726
rect 18844 7474 18900 7476
rect 18844 7422 18846 7474
rect 18846 7422 18898 7474
rect 18898 7422 18900 7474
rect 18844 7420 18900 7422
rect 18060 7196 18116 7252
rect 18396 7084 18452 7140
rect 18732 6860 18788 6916
rect 18956 6802 19012 6804
rect 18956 6750 18958 6802
rect 18958 6750 19010 6802
rect 19010 6750 19012 6802
rect 18956 6748 19012 6750
rect 18620 6690 18676 6692
rect 18620 6638 18622 6690
rect 18622 6638 18674 6690
rect 18674 6638 18676 6690
rect 18620 6636 18676 6638
rect 18396 6524 18452 6580
rect 17724 6130 17780 6132
rect 17724 6078 17726 6130
rect 17726 6078 17778 6130
rect 17778 6078 17780 6130
rect 17724 6076 17780 6078
rect 17388 5628 17444 5684
rect 17500 4450 17556 4452
rect 17500 4398 17502 4450
rect 17502 4398 17554 4450
rect 17554 4398 17556 4450
rect 17500 4396 17556 4398
rect 19180 6300 19236 6356
rect 18732 6188 18788 6244
rect 18732 5852 18788 5908
rect 19068 5964 19124 6020
rect 18732 5234 18788 5236
rect 18732 5182 18734 5234
rect 18734 5182 18786 5234
rect 18786 5182 18788 5234
rect 18732 5180 18788 5182
rect 18508 4956 18564 5012
rect 19292 5682 19348 5684
rect 19292 5630 19294 5682
rect 19294 5630 19346 5682
rect 19346 5630 19348 5682
rect 19292 5628 19348 5630
rect 19852 9602 19908 9604
rect 19852 9550 19854 9602
rect 19854 9550 19906 9602
rect 19906 9550 19908 9602
rect 19852 9548 19908 9550
rect 21084 10610 21140 10612
rect 21084 10558 21086 10610
rect 21086 10558 21138 10610
rect 21138 10558 21140 10610
rect 21084 10556 21140 10558
rect 20636 10108 20692 10164
rect 21532 10108 21588 10164
rect 20748 9772 20804 9828
rect 21308 9996 21364 10052
rect 21644 9996 21700 10052
rect 21980 10444 22036 10500
rect 21644 9772 21700 9828
rect 22652 9938 22708 9940
rect 22652 9886 22654 9938
rect 22654 9886 22706 9938
rect 22706 9886 22708 9938
rect 22652 9884 22708 9886
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20188 9212 20244 9268
rect 19852 9154 19908 9156
rect 19852 9102 19854 9154
rect 19854 9102 19906 9154
rect 19906 9102 19908 9154
rect 19852 9100 19908 9102
rect 21308 9548 21364 9604
rect 20524 8204 20580 8260
rect 20748 9324 20804 9380
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19628 7532 19684 7588
rect 20412 7980 20468 8036
rect 20412 7362 20468 7364
rect 20412 7310 20414 7362
rect 20414 7310 20466 7362
rect 20466 7310 20468 7362
rect 20412 7308 20468 7310
rect 20188 6636 20244 6692
rect 20300 6578 20356 6580
rect 20300 6526 20302 6578
rect 20302 6526 20354 6578
rect 20354 6526 20356 6578
rect 20300 6524 20356 6526
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20188 6300 20244 6356
rect 20044 6244 20100 6246
rect 21196 9100 21252 9156
rect 20972 8092 21028 8148
rect 20748 7420 20804 7476
rect 21644 9324 21700 9380
rect 21532 9212 21588 9268
rect 21644 9154 21700 9156
rect 21644 9102 21646 9154
rect 21646 9102 21698 9154
rect 21698 9102 21700 9154
rect 21644 9100 21700 9102
rect 21308 8876 21364 8932
rect 22204 8930 22260 8932
rect 22204 8878 22206 8930
rect 22206 8878 22258 8930
rect 22258 8878 22260 8930
rect 22204 8876 22260 8878
rect 21644 8428 21700 8484
rect 21084 7196 21140 7252
rect 20748 6636 20804 6692
rect 19740 5740 19796 5796
rect 20636 5852 20692 5908
rect 19292 5068 19348 5124
rect 17388 3724 17444 3780
rect 13580 3442 13636 3444
rect 13580 3390 13582 3442
rect 13582 3390 13634 3442
rect 13634 3390 13636 3442
rect 13580 3388 13636 3390
rect 15708 3612 15764 3668
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20748 5740 20804 5796
rect 21308 7698 21364 7700
rect 21308 7646 21310 7698
rect 21310 7646 21362 7698
rect 21362 7646 21364 7698
rect 21308 7644 21364 7646
rect 21420 7084 21476 7140
rect 21196 5740 21252 5796
rect 21420 5122 21476 5124
rect 21420 5070 21422 5122
rect 21422 5070 21474 5122
rect 21474 5070 21476 5122
rect 21420 5068 21476 5070
rect 20188 4396 20244 4452
rect 20972 4396 21028 4452
rect 19964 4060 20020 4116
rect 20748 3778 20804 3780
rect 20748 3726 20750 3778
rect 20750 3726 20802 3778
rect 20802 3726 20804 3778
rect 20748 3724 20804 3726
rect 20188 3442 20244 3444
rect 20188 3390 20190 3442
rect 20190 3390 20242 3442
rect 20242 3390 20244 3442
rect 20188 3388 20244 3390
rect 21756 5740 21812 5796
rect 21532 4284 21588 4340
rect 21084 3778 21140 3780
rect 21084 3726 21086 3778
rect 21086 3726 21138 3778
rect 21138 3726 21140 3778
rect 21084 3724 21140 3726
rect 22652 7980 22708 8036
rect 23996 14418 24052 14420
rect 23996 14366 23998 14418
rect 23998 14366 24050 14418
rect 24050 14366 24052 14418
rect 23996 14364 24052 14366
rect 22988 13692 23044 13748
rect 23772 13132 23828 13188
rect 22876 11618 22932 11620
rect 22876 11566 22878 11618
rect 22878 11566 22930 11618
rect 22930 11566 22932 11618
rect 22876 11564 22932 11566
rect 23548 12066 23604 12068
rect 23548 12014 23550 12066
rect 23550 12014 23602 12066
rect 23602 12014 23604 12066
rect 23548 12012 23604 12014
rect 22876 10498 22932 10500
rect 22876 10446 22878 10498
rect 22878 10446 22930 10498
rect 22930 10446 22932 10498
rect 22876 10444 22932 10446
rect 22988 9042 23044 9044
rect 22988 8990 22990 9042
rect 22990 8990 23042 9042
rect 23042 8990 23044 9042
rect 22988 8988 23044 8990
rect 23324 11676 23380 11732
rect 23212 11282 23268 11284
rect 23212 11230 23214 11282
rect 23214 11230 23266 11282
rect 23266 11230 23268 11282
rect 23212 11228 23268 11230
rect 24332 13580 24388 13636
rect 24108 13020 24164 13076
rect 23884 12738 23940 12740
rect 23884 12686 23886 12738
rect 23886 12686 23938 12738
rect 23938 12686 23940 12738
rect 23884 12684 23940 12686
rect 24220 12236 24276 12292
rect 23884 12124 23940 12180
rect 24332 11282 24388 11284
rect 24332 11230 24334 11282
rect 24334 11230 24386 11282
rect 24386 11230 24388 11282
rect 24332 11228 24388 11230
rect 23772 11004 23828 11060
rect 24220 9772 24276 9828
rect 22764 7868 22820 7924
rect 22092 7308 22148 7364
rect 22092 6412 22148 6468
rect 22428 5068 22484 5124
rect 22540 6076 22596 6132
rect 23212 7196 23268 7252
rect 23324 6748 23380 6804
rect 23772 8876 23828 8932
rect 23884 9100 23940 9156
rect 23436 7644 23492 7700
rect 23212 6300 23268 6356
rect 23660 8764 23716 8820
rect 23660 8092 23716 8148
rect 23548 6524 23604 6580
rect 23772 6466 23828 6468
rect 23772 6414 23774 6466
rect 23774 6414 23826 6466
rect 23826 6414 23828 6466
rect 23772 6412 23828 6414
rect 24556 15260 24612 15316
rect 24668 15202 24724 15204
rect 24668 15150 24670 15202
rect 24670 15150 24722 15202
rect 24722 15150 24724 15202
rect 24668 15148 24724 15150
rect 24668 14252 24724 14308
rect 25676 16716 25732 16772
rect 25900 15426 25956 15428
rect 25900 15374 25902 15426
rect 25902 15374 25954 15426
rect 25954 15374 25956 15426
rect 25900 15372 25956 15374
rect 25452 15148 25508 15204
rect 25228 14812 25284 14868
rect 25340 14924 25396 14980
rect 25004 14364 25060 14420
rect 25004 12684 25060 12740
rect 24892 9938 24948 9940
rect 24892 9886 24894 9938
rect 24894 9886 24946 9938
rect 24946 9886 24948 9938
rect 24892 9884 24948 9886
rect 24668 9154 24724 9156
rect 24668 9102 24670 9154
rect 24670 9102 24722 9154
rect 24722 9102 24724 9154
rect 24668 9100 24724 9102
rect 24556 8876 24612 8932
rect 23884 6300 23940 6356
rect 24108 6300 24164 6356
rect 24220 7532 24276 7588
rect 23996 6076 24052 6132
rect 25564 14252 25620 14308
rect 25676 14140 25732 14196
rect 26124 14812 26180 14868
rect 26572 21084 26628 21140
rect 26460 20802 26516 20804
rect 26460 20750 26462 20802
rect 26462 20750 26514 20802
rect 26514 20750 26516 20802
rect 26460 20748 26516 20750
rect 26348 19180 26404 19236
rect 26572 20524 26628 20580
rect 26460 18450 26516 18452
rect 26460 18398 26462 18450
rect 26462 18398 26514 18450
rect 26514 18398 26516 18450
rect 26460 18396 26516 18398
rect 26908 20524 26964 20580
rect 26684 20188 26740 20244
rect 26908 20018 26964 20020
rect 26908 19966 26910 20018
rect 26910 19966 26962 20018
rect 26962 19966 26964 20018
rect 26908 19964 26964 19966
rect 27468 22988 27524 23044
rect 29036 34130 29092 34132
rect 29036 34078 29038 34130
rect 29038 34078 29090 34130
rect 29090 34078 29092 34130
rect 29036 34076 29092 34078
rect 29260 34130 29316 34132
rect 29260 34078 29262 34130
rect 29262 34078 29314 34130
rect 29314 34078 29316 34130
rect 29260 34076 29316 34078
rect 28924 33964 28980 34020
rect 28924 33628 28980 33684
rect 28924 33068 28980 33124
rect 28476 30716 28532 30772
rect 28028 27916 28084 27972
rect 28252 25676 28308 25732
rect 28028 25618 28084 25620
rect 28028 25566 28030 25618
rect 28030 25566 28082 25618
rect 28082 25566 28084 25618
rect 28028 25564 28084 25566
rect 28140 25506 28196 25508
rect 28140 25454 28142 25506
rect 28142 25454 28194 25506
rect 28194 25454 28196 25506
rect 28140 25452 28196 25454
rect 27916 22652 27972 22708
rect 28028 25228 28084 25284
rect 28252 24610 28308 24612
rect 28252 24558 28254 24610
rect 28254 24558 28306 24610
rect 28306 24558 28308 24610
rect 28252 24556 28308 24558
rect 28476 26684 28532 26740
rect 28588 25452 28644 25508
rect 28364 24220 28420 24276
rect 28812 30156 28868 30212
rect 28140 22876 28196 22932
rect 27244 21980 27300 22036
rect 27804 21980 27860 22036
rect 27132 21756 27188 21812
rect 27580 21756 27636 21812
rect 28028 21586 28084 21588
rect 28028 21534 28030 21586
rect 28030 21534 28082 21586
rect 28082 21534 28084 21586
rect 28028 21532 28084 21534
rect 28364 21474 28420 21476
rect 28364 21422 28366 21474
rect 28366 21422 28418 21474
rect 28418 21422 28420 21474
rect 28364 21420 28420 21422
rect 28252 21308 28308 21364
rect 28252 21084 28308 21140
rect 27244 20802 27300 20804
rect 27244 20750 27246 20802
rect 27246 20750 27298 20802
rect 27298 20750 27300 20802
rect 27244 20748 27300 20750
rect 27804 20300 27860 20356
rect 28028 20636 28084 20692
rect 27132 19852 27188 19908
rect 26796 19628 26852 19684
rect 26684 18844 26740 18900
rect 25788 13356 25844 13412
rect 27020 18844 27076 18900
rect 25452 12850 25508 12852
rect 25452 12798 25454 12850
rect 25454 12798 25506 12850
rect 25506 12798 25508 12850
rect 25452 12796 25508 12798
rect 26460 17388 26516 17444
rect 26796 18060 26852 18116
rect 28028 20076 28084 20132
rect 27468 19964 27524 20020
rect 27692 19964 27748 20020
rect 27580 19852 27636 19908
rect 27692 19628 27748 19684
rect 28252 20018 28308 20020
rect 28252 19966 28254 20018
rect 28254 19966 28306 20018
rect 28306 19966 28308 20018
rect 28252 19964 28308 19966
rect 27356 19122 27412 19124
rect 27356 19070 27358 19122
rect 27358 19070 27410 19122
rect 27410 19070 27412 19122
rect 27356 19068 27412 19070
rect 27692 19122 27748 19124
rect 27692 19070 27694 19122
rect 27694 19070 27746 19122
rect 27746 19070 27748 19122
rect 27692 19068 27748 19070
rect 27132 18620 27188 18676
rect 27692 18674 27748 18676
rect 27692 18622 27694 18674
rect 27694 18622 27746 18674
rect 27746 18622 27748 18674
rect 27692 18620 27748 18622
rect 27020 17836 27076 17892
rect 27468 17724 27524 17780
rect 26684 17276 26740 17332
rect 26796 17500 26852 17556
rect 28252 18844 28308 18900
rect 28364 18732 28420 18788
rect 28812 24946 28868 24948
rect 28812 24894 28814 24946
rect 28814 24894 28866 24946
rect 28866 24894 28868 24946
rect 28812 24892 28868 24894
rect 28700 22092 28756 22148
rect 28812 23212 28868 23268
rect 28700 21644 28756 21700
rect 28700 21308 28756 21364
rect 28812 19964 28868 20020
rect 29148 33180 29204 33236
rect 29372 32956 29428 33012
rect 29820 35420 29876 35476
rect 31052 35980 31108 36036
rect 30940 35922 30996 35924
rect 30940 35870 30942 35922
rect 30942 35870 30994 35922
rect 30994 35870 30996 35922
rect 30940 35868 30996 35870
rect 30380 35644 30436 35700
rect 30492 35420 30548 35476
rect 29932 35308 29988 35364
rect 29820 34802 29876 34804
rect 29820 34750 29822 34802
rect 29822 34750 29874 34802
rect 29874 34750 29876 34802
rect 29820 34748 29876 34750
rect 29708 34524 29764 34580
rect 29708 34300 29764 34356
rect 29708 33628 29764 33684
rect 29932 33346 29988 33348
rect 29932 33294 29934 33346
rect 29934 33294 29986 33346
rect 29986 33294 29988 33346
rect 29932 33292 29988 33294
rect 29932 32956 29988 33012
rect 29596 32450 29652 32452
rect 29596 32398 29598 32450
rect 29598 32398 29650 32450
rect 29650 32398 29652 32450
rect 29596 32396 29652 32398
rect 30268 34412 30324 34468
rect 31388 35756 31444 35812
rect 30828 34524 30884 34580
rect 30604 33628 30660 33684
rect 30716 33964 30772 34020
rect 30380 33404 30436 33460
rect 31052 33964 31108 34020
rect 30940 33346 30996 33348
rect 30940 33294 30942 33346
rect 30942 33294 30994 33346
rect 30994 33294 30996 33346
rect 30940 33292 30996 33294
rect 30716 33234 30772 33236
rect 30716 33182 30718 33234
rect 30718 33182 30770 33234
rect 30770 33182 30772 33234
rect 30716 33180 30772 33182
rect 30604 32844 30660 32900
rect 30604 31554 30660 31556
rect 30604 31502 30606 31554
rect 30606 31502 30658 31554
rect 30658 31502 30660 31554
rect 30604 31500 30660 31502
rect 31164 31612 31220 31668
rect 30940 31500 30996 31556
rect 32396 38556 32452 38612
rect 32508 37154 32564 37156
rect 32508 37102 32510 37154
rect 32510 37102 32562 37154
rect 32562 37102 32564 37154
rect 32508 37100 32564 37102
rect 31948 35810 32004 35812
rect 31948 35758 31950 35810
rect 31950 35758 32002 35810
rect 32002 35758 32004 35810
rect 31948 35756 32004 35758
rect 31724 35644 31780 35700
rect 31612 34412 31668 34468
rect 31500 34188 31556 34244
rect 32396 35756 32452 35812
rect 32284 35698 32340 35700
rect 32284 35646 32286 35698
rect 32286 35646 32338 35698
rect 32338 35646 32340 35698
rect 32284 35644 32340 35646
rect 32060 34018 32116 34020
rect 32060 33966 32062 34018
rect 32062 33966 32114 34018
rect 32114 33966 32116 34018
rect 32060 33964 32116 33966
rect 31724 33180 31780 33236
rect 31500 33122 31556 33124
rect 31500 33070 31502 33122
rect 31502 33070 31554 33122
rect 31554 33070 31556 33122
rect 31500 33068 31556 33070
rect 33068 38668 33124 38724
rect 32956 37772 33012 37828
rect 33068 37100 33124 37156
rect 33068 36652 33124 36708
rect 33292 38444 33348 38500
rect 33852 38444 33908 38500
rect 35980 47234 36036 47236
rect 35980 47182 35982 47234
rect 35982 47182 36034 47234
rect 36034 47182 36036 47234
rect 35980 47180 36036 47182
rect 38892 48354 38948 48356
rect 38892 48302 38894 48354
rect 38894 48302 38946 48354
rect 38946 48302 38948 48354
rect 38892 48300 38948 48302
rect 38220 47346 38276 47348
rect 38220 47294 38222 47346
rect 38222 47294 38274 47346
rect 38274 47294 38276 47346
rect 38220 47292 38276 47294
rect 37996 47180 38052 47236
rect 38332 47180 38388 47236
rect 37100 46956 37156 47012
rect 34972 46562 35028 46564
rect 34972 46510 34974 46562
rect 34974 46510 35026 46562
rect 35026 46510 35028 46562
rect 34972 46508 35028 46510
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 38892 47292 38948 47348
rect 38668 46786 38724 46788
rect 38668 46734 38670 46786
rect 38670 46734 38722 46786
rect 38722 46734 38724 46786
rect 38668 46732 38724 46734
rect 40012 48300 40068 48356
rect 39228 46956 39284 47012
rect 40236 46956 40292 47012
rect 34636 43932 34692 43988
rect 34412 43596 34468 43652
rect 34076 43538 34132 43540
rect 34076 43486 34078 43538
rect 34078 43486 34130 43538
rect 34130 43486 34132 43538
rect 34076 43484 34132 43486
rect 34188 41356 34244 41412
rect 34076 41020 34132 41076
rect 34076 40236 34132 40292
rect 34524 39394 34580 39396
rect 34524 39342 34526 39394
rect 34526 39342 34578 39394
rect 34578 39342 34580 39394
rect 34524 39340 34580 39342
rect 34972 45276 35028 45332
rect 37436 45330 37492 45332
rect 37436 45278 37438 45330
rect 37438 45278 37490 45330
rect 37490 45278 37492 45330
rect 37436 45276 37492 45278
rect 34972 44210 35028 44212
rect 34972 44158 34974 44210
rect 34974 44158 35026 44210
rect 35026 44158 35028 44210
rect 34972 44156 35028 44158
rect 38108 45276 38164 45332
rect 40012 46732 40068 46788
rect 40012 46060 40068 46116
rect 41692 47180 41748 47236
rect 39788 45164 39844 45220
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35084 44044 35140 44100
rect 34860 43596 34916 43652
rect 35644 44098 35700 44100
rect 35644 44046 35646 44098
rect 35646 44046 35698 44098
rect 35698 44046 35700 44098
rect 35644 44044 35700 44046
rect 36316 43708 36372 43764
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 41132 46114 41188 46116
rect 41132 46062 41134 46114
rect 41134 46062 41186 46114
rect 41186 46062 41188 46114
rect 41132 46060 41188 46062
rect 37772 41916 37828 41972
rect 35644 41804 35700 41860
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35308 41410 35364 41412
rect 35308 41358 35310 41410
rect 35310 41358 35362 41410
rect 35362 41358 35364 41410
rect 35308 41356 35364 41358
rect 36092 41356 36148 41412
rect 34972 41020 35028 41076
rect 35532 41074 35588 41076
rect 35532 41022 35534 41074
rect 35534 41022 35586 41074
rect 35586 41022 35588 41074
rect 35532 41020 35588 41022
rect 38780 41804 38836 41860
rect 39340 41970 39396 41972
rect 39340 41918 39342 41970
rect 39342 41918 39394 41970
rect 39394 41918 39396 41970
rect 39340 41916 39396 41918
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35532 39340 35588 39396
rect 35084 38946 35140 38948
rect 35084 38894 35086 38946
rect 35086 38894 35138 38946
rect 35138 38894 35140 38946
rect 35084 38892 35140 38894
rect 34188 38610 34244 38612
rect 34188 38558 34190 38610
rect 34190 38558 34242 38610
rect 34242 38558 34244 38610
rect 34188 38556 34244 38558
rect 33964 38332 34020 38388
rect 33964 38108 34020 38164
rect 33628 37100 33684 37156
rect 32732 36316 32788 36372
rect 32396 33964 32452 34020
rect 32508 33628 32564 33684
rect 32172 32844 32228 32900
rect 32396 33122 32452 33124
rect 32396 33070 32398 33122
rect 32398 33070 32450 33122
rect 32450 33070 32452 33122
rect 32396 33068 32452 33070
rect 32060 32732 32116 32788
rect 31948 32674 32004 32676
rect 31948 32622 31950 32674
rect 31950 32622 32002 32674
rect 32002 32622 32004 32674
rect 31948 32620 32004 32622
rect 30828 31218 30884 31220
rect 30828 31166 30830 31218
rect 30830 31166 30882 31218
rect 30882 31166 30884 31218
rect 30828 31164 30884 31166
rect 29372 29538 29428 29540
rect 29372 29486 29374 29538
rect 29374 29486 29426 29538
rect 29426 29486 29428 29538
rect 29372 29484 29428 29486
rect 29484 29260 29540 29316
rect 29820 28700 29876 28756
rect 29484 28642 29540 28644
rect 29484 28590 29486 28642
rect 29486 28590 29538 28642
rect 29538 28590 29540 28642
rect 29484 28588 29540 28590
rect 29932 28140 29988 28196
rect 31388 32172 31444 32228
rect 30156 29484 30212 29540
rect 30492 29260 30548 29316
rect 30156 28642 30212 28644
rect 30156 28590 30158 28642
rect 30158 28590 30210 28642
rect 30210 28590 30212 28642
rect 30156 28588 30212 28590
rect 30380 28364 30436 28420
rect 30044 27468 30100 27524
rect 29372 25788 29428 25844
rect 29148 24892 29204 24948
rect 29148 24722 29204 24724
rect 29148 24670 29150 24722
rect 29150 24670 29202 24722
rect 29202 24670 29204 24722
rect 29148 24668 29204 24670
rect 29148 23938 29204 23940
rect 29148 23886 29150 23938
rect 29150 23886 29202 23938
rect 29202 23886 29204 23938
rect 29148 23884 29204 23886
rect 29036 20018 29092 20020
rect 29036 19966 29038 20018
rect 29038 19966 29090 20018
rect 29090 19966 29092 20018
rect 29036 19964 29092 19966
rect 30044 26460 30100 26516
rect 30044 25788 30100 25844
rect 29820 25452 29876 25508
rect 30268 25506 30324 25508
rect 30268 25454 30270 25506
rect 30270 25454 30322 25506
rect 30322 25454 30324 25506
rect 30268 25452 30324 25454
rect 32060 31890 32116 31892
rect 32060 31838 32062 31890
rect 32062 31838 32114 31890
rect 32114 31838 32116 31890
rect 32060 31836 32116 31838
rect 33292 34242 33348 34244
rect 33292 34190 33294 34242
rect 33294 34190 33346 34242
rect 33346 34190 33348 34242
rect 33292 34188 33348 34190
rect 33740 35420 33796 35476
rect 33852 35810 33908 35812
rect 33852 35758 33854 35810
rect 33854 35758 33906 35810
rect 33906 35758 33908 35810
rect 33852 35756 33908 35758
rect 33852 35308 33908 35364
rect 34300 37826 34356 37828
rect 34300 37774 34302 37826
rect 34302 37774 34354 37826
rect 34354 37774 34356 37826
rect 34300 37772 34356 37774
rect 34076 36370 34132 36372
rect 34076 36318 34078 36370
rect 34078 36318 34130 36370
rect 34130 36318 34132 36370
rect 34076 36316 34132 36318
rect 34188 34636 34244 34692
rect 33516 34018 33572 34020
rect 33516 33966 33518 34018
rect 33518 33966 33570 34018
rect 33570 33966 33572 34018
rect 33516 33964 33572 33966
rect 33180 33628 33236 33684
rect 32844 33234 32900 33236
rect 32844 33182 32846 33234
rect 32846 33182 32898 33234
rect 32898 33182 32900 33234
rect 32844 33180 32900 33182
rect 32732 33068 32788 33124
rect 32284 32060 32340 32116
rect 32396 32396 32452 32452
rect 31500 31554 31556 31556
rect 31500 31502 31502 31554
rect 31502 31502 31554 31554
rect 31554 31502 31556 31554
rect 31500 31500 31556 31502
rect 31164 29260 31220 29316
rect 31724 31218 31780 31220
rect 31724 31166 31726 31218
rect 31726 31166 31778 31218
rect 31778 31166 31780 31218
rect 31724 31164 31780 31166
rect 30604 28812 30660 28868
rect 30716 29036 30772 29092
rect 31948 30156 32004 30212
rect 31836 29708 31892 29764
rect 31164 28364 31220 28420
rect 31500 28700 31556 28756
rect 30604 27970 30660 27972
rect 30604 27918 30606 27970
rect 30606 27918 30658 27970
rect 30658 27918 30660 27970
rect 30604 27916 30660 27918
rect 30940 27580 30996 27636
rect 30940 27244 30996 27300
rect 29708 24668 29764 24724
rect 29596 24220 29652 24276
rect 29372 22988 29428 23044
rect 29372 22428 29428 22484
rect 30044 24220 30100 24276
rect 29708 22428 29764 22484
rect 30044 23324 30100 23380
rect 29596 22258 29652 22260
rect 29596 22206 29598 22258
rect 29598 22206 29650 22258
rect 29650 22206 29652 22258
rect 29596 22204 29652 22206
rect 29708 21698 29764 21700
rect 29708 21646 29710 21698
rect 29710 21646 29762 21698
rect 29762 21646 29764 21698
rect 29708 21644 29764 21646
rect 29596 21586 29652 21588
rect 29596 21534 29598 21586
rect 29598 21534 29650 21586
rect 29650 21534 29652 21586
rect 29596 21532 29652 21534
rect 29820 21420 29876 21476
rect 29260 20860 29316 20916
rect 29372 20076 29428 20132
rect 29260 19852 29316 19908
rect 28924 19404 28980 19460
rect 28588 19346 28644 19348
rect 28588 19294 28590 19346
rect 28590 19294 28642 19346
rect 28642 19294 28644 19346
rect 28588 19292 28644 19294
rect 29372 19292 29428 19348
rect 29484 19964 29540 20020
rect 28700 18732 28756 18788
rect 29036 18562 29092 18564
rect 29036 18510 29038 18562
rect 29038 18510 29090 18562
rect 29090 18510 29092 18562
rect 29036 18508 29092 18510
rect 28252 18284 28308 18340
rect 27692 17554 27748 17556
rect 27692 17502 27694 17554
rect 27694 17502 27746 17554
rect 27746 17502 27748 17554
rect 27692 17500 27748 17502
rect 27020 17388 27076 17444
rect 27468 17442 27524 17444
rect 27468 17390 27470 17442
rect 27470 17390 27522 17442
rect 27522 17390 27524 17442
rect 27468 17388 27524 17390
rect 27356 16828 27412 16884
rect 27244 16716 27300 16772
rect 29708 21362 29764 21364
rect 29708 21310 29710 21362
rect 29710 21310 29762 21362
rect 29762 21310 29764 21362
rect 29708 21308 29764 21310
rect 30380 24332 30436 24388
rect 30492 24220 30548 24276
rect 30044 22428 30100 22484
rect 30828 26796 30884 26852
rect 31276 27074 31332 27076
rect 31276 27022 31278 27074
rect 31278 27022 31330 27074
rect 31330 27022 31332 27074
rect 31276 27020 31332 27022
rect 31836 29036 31892 29092
rect 31164 26796 31220 26852
rect 30828 25788 30884 25844
rect 31500 25452 31556 25508
rect 31948 28082 32004 28084
rect 31948 28030 31950 28082
rect 31950 28030 32002 28082
rect 32002 28030 32004 28082
rect 31948 28028 32004 28030
rect 32508 31724 32564 31780
rect 32956 32396 33012 32452
rect 33292 33516 33348 33572
rect 34524 35308 34580 35364
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 36092 38892 36148 38948
rect 37212 38892 37268 38948
rect 39228 40908 39284 40964
rect 39004 38834 39060 38836
rect 39004 38782 39006 38834
rect 39006 38782 39058 38834
rect 39058 38782 39060 38834
rect 39004 38780 39060 38782
rect 35868 38108 35924 38164
rect 37996 38108 38052 38164
rect 35868 37938 35924 37940
rect 35868 37886 35870 37938
rect 35870 37886 35922 37938
rect 35922 37886 35924 37938
rect 35868 37884 35924 37886
rect 37660 37938 37716 37940
rect 37660 37886 37662 37938
rect 37662 37886 37714 37938
rect 37714 37886 37716 37938
rect 37660 37884 37716 37886
rect 39116 38050 39172 38052
rect 39116 37998 39118 38050
rect 39118 37998 39170 38050
rect 39170 37998 39172 38050
rect 39116 37996 39172 37998
rect 36988 37548 37044 37604
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 36092 35532 36148 35588
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35532 34914 35588 34916
rect 35532 34862 35534 34914
rect 35534 34862 35586 34914
rect 35586 34862 35588 34914
rect 35532 34860 35588 34862
rect 36092 34802 36148 34804
rect 36092 34750 36094 34802
rect 36094 34750 36146 34802
rect 36146 34750 36148 34802
rect 36092 34748 36148 34750
rect 34524 34242 34580 34244
rect 34524 34190 34526 34242
rect 34526 34190 34578 34242
rect 34578 34190 34580 34242
rect 34524 34188 34580 34190
rect 34524 33964 34580 34020
rect 34748 34076 34804 34132
rect 36204 34242 36260 34244
rect 36204 34190 36206 34242
rect 36206 34190 36258 34242
rect 36258 34190 36260 34242
rect 36204 34188 36260 34190
rect 35868 34076 35924 34132
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35084 33346 35140 33348
rect 35084 33294 35086 33346
rect 35086 33294 35138 33346
rect 35138 33294 35140 33346
rect 35084 33292 35140 33294
rect 33628 32450 33684 32452
rect 33628 32398 33630 32450
rect 33630 32398 33682 32450
rect 33682 32398 33684 32450
rect 33628 32396 33684 32398
rect 33964 32562 34020 32564
rect 33964 32510 33966 32562
rect 33966 32510 34018 32562
rect 34018 32510 34020 32562
rect 33964 32508 34020 32510
rect 33740 32172 33796 32228
rect 32844 31554 32900 31556
rect 32844 31502 32846 31554
rect 32846 31502 32898 31554
rect 32898 31502 32900 31554
rect 32844 31500 32900 31502
rect 32284 30210 32340 30212
rect 32284 30158 32286 30210
rect 32286 30158 32338 30210
rect 32338 30158 32340 30210
rect 32284 30156 32340 30158
rect 33292 29372 33348 29428
rect 33404 29314 33460 29316
rect 33404 29262 33406 29314
rect 33406 29262 33458 29314
rect 33458 29262 33460 29314
rect 33404 29260 33460 29262
rect 33628 31500 33684 31556
rect 32620 28642 32676 28644
rect 32620 28590 32622 28642
rect 32622 28590 32674 28642
rect 32674 28590 32676 28642
rect 32620 28588 32676 28590
rect 33628 30828 33684 30884
rect 33628 29036 33684 29092
rect 32284 28028 32340 28084
rect 32172 27580 32228 27636
rect 31836 27132 31892 27188
rect 31836 26962 31892 26964
rect 31836 26910 31838 26962
rect 31838 26910 31890 26962
rect 31890 26910 31892 26962
rect 31836 26908 31892 26910
rect 31836 25506 31892 25508
rect 31836 25454 31838 25506
rect 31838 25454 31890 25506
rect 31890 25454 31892 25506
rect 31836 25452 31892 25454
rect 31612 25340 31668 25396
rect 31164 25228 31220 25284
rect 31164 24444 31220 24500
rect 31276 24332 31332 24388
rect 30492 23212 30548 23268
rect 30380 22316 30436 22372
rect 30156 20972 30212 21028
rect 29932 20130 29988 20132
rect 29932 20078 29934 20130
rect 29934 20078 29986 20130
rect 29986 20078 29988 20130
rect 29932 20076 29988 20078
rect 30716 22258 30772 22260
rect 30716 22206 30718 22258
rect 30718 22206 30770 22258
rect 30770 22206 30772 22258
rect 30716 22204 30772 22206
rect 30604 21756 30660 21812
rect 30268 20018 30324 20020
rect 30268 19966 30270 20018
rect 30270 19966 30322 20018
rect 30322 19966 30324 20018
rect 30268 19964 30324 19966
rect 29596 19404 29652 19460
rect 29596 18732 29652 18788
rect 29372 18172 29428 18228
rect 29484 18396 29540 18452
rect 28812 17836 28868 17892
rect 29484 17666 29540 17668
rect 29484 17614 29486 17666
rect 29486 17614 29538 17666
rect 29538 17614 29540 17666
rect 29484 17612 29540 17614
rect 28028 16882 28084 16884
rect 28028 16830 28030 16882
rect 28030 16830 28082 16882
rect 28082 16830 28084 16882
rect 28028 16828 28084 16830
rect 27916 16156 27972 16212
rect 27020 15820 27076 15876
rect 27132 15596 27188 15652
rect 26460 13468 26516 13524
rect 25900 12348 25956 12404
rect 27244 15260 27300 15316
rect 27132 14700 27188 14756
rect 27580 15148 27636 15204
rect 27468 14642 27524 14644
rect 27468 14590 27470 14642
rect 27470 14590 27522 14642
rect 27522 14590 27524 14642
rect 27468 14588 27524 14590
rect 27692 14700 27748 14756
rect 27916 14924 27972 14980
rect 27132 13468 27188 13524
rect 26908 13020 26964 13076
rect 26124 12684 26180 12740
rect 26460 12236 26516 12292
rect 26236 10108 26292 10164
rect 26796 12572 26852 12628
rect 27020 12460 27076 12516
rect 26796 12236 26852 12292
rect 26684 9996 26740 10052
rect 25788 9772 25844 9828
rect 27356 12962 27412 12964
rect 27356 12910 27358 12962
rect 27358 12910 27410 12962
rect 27410 12910 27412 12962
rect 27356 12908 27412 12910
rect 27356 12348 27412 12404
rect 27356 12124 27412 12180
rect 27916 13132 27972 13188
rect 28700 16828 28756 16884
rect 28364 16210 28420 16212
rect 28364 16158 28366 16210
rect 28366 16158 28418 16210
rect 28418 16158 28420 16210
rect 28364 16156 28420 16158
rect 28924 16156 28980 16212
rect 28252 16098 28308 16100
rect 28252 16046 28254 16098
rect 28254 16046 28306 16098
rect 28306 16046 28308 16098
rect 28252 16044 28308 16046
rect 28252 15148 28308 15204
rect 28588 15484 28644 15540
rect 28364 14028 28420 14084
rect 29484 16098 29540 16100
rect 29484 16046 29486 16098
rect 29486 16046 29538 16098
rect 29538 16046 29540 16098
rect 29484 16044 29540 16046
rect 28588 14252 28644 14308
rect 28476 13804 28532 13860
rect 28364 13580 28420 13636
rect 28588 13746 28644 13748
rect 28588 13694 28590 13746
rect 28590 13694 28642 13746
rect 28642 13694 28644 13746
rect 28588 13692 28644 13694
rect 30604 20578 30660 20580
rect 30604 20526 30606 20578
rect 30606 20526 30658 20578
rect 30658 20526 30660 20578
rect 30604 20524 30660 20526
rect 29708 14140 29764 14196
rect 29820 17836 29876 17892
rect 29932 17276 29988 17332
rect 30044 17388 30100 17444
rect 29932 17106 29988 17108
rect 29932 17054 29934 17106
rect 29934 17054 29986 17106
rect 29986 17054 29988 17106
rect 29932 17052 29988 17054
rect 29932 16658 29988 16660
rect 29932 16606 29934 16658
rect 29934 16606 29986 16658
rect 29986 16606 29988 16658
rect 29932 16604 29988 16606
rect 28364 13244 28420 13300
rect 28252 13186 28308 13188
rect 28252 13134 28254 13186
rect 28254 13134 28306 13186
rect 28306 13134 28308 13186
rect 28252 13132 28308 13134
rect 29148 13244 29204 13300
rect 27692 12684 27748 12740
rect 28140 12290 28196 12292
rect 28140 12238 28142 12290
rect 28142 12238 28194 12290
rect 28194 12238 28196 12290
rect 28140 12236 28196 12238
rect 27916 11676 27972 11732
rect 27804 11340 27860 11396
rect 27804 10444 27860 10500
rect 26908 9660 26964 9716
rect 25228 9154 25284 9156
rect 25228 9102 25230 9154
rect 25230 9102 25282 9154
rect 25282 9102 25284 9154
rect 25228 9100 25284 9102
rect 25228 8652 25284 8708
rect 25228 8092 25284 8148
rect 25004 7420 25060 7476
rect 25004 6578 25060 6580
rect 25004 6526 25006 6578
rect 25006 6526 25058 6578
rect 25058 6526 25060 6578
rect 25004 6524 25060 6526
rect 25228 6412 25284 6468
rect 24668 6188 24724 6244
rect 24444 6130 24500 6132
rect 24444 6078 24446 6130
rect 24446 6078 24498 6130
rect 24498 6078 24500 6130
rect 24444 6076 24500 6078
rect 25340 6300 25396 6356
rect 27580 9042 27636 9044
rect 27580 8990 27582 9042
rect 27582 8990 27634 9042
rect 27634 8990 27636 9042
rect 27580 8988 27636 8990
rect 25676 8370 25732 8372
rect 25676 8318 25678 8370
rect 25678 8318 25730 8370
rect 25730 8318 25732 8370
rect 25676 8316 25732 8318
rect 25676 7532 25732 7588
rect 25564 7250 25620 7252
rect 25564 7198 25566 7250
rect 25566 7198 25618 7250
rect 25618 7198 25620 7250
rect 25564 7196 25620 7198
rect 25900 8316 25956 8372
rect 27132 8316 27188 8372
rect 27804 8316 27860 8372
rect 28364 12460 28420 12516
rect 28140 10444 28196 10500
rect 28364 12236 28420 12292
rect 28140 9996 28196 10052
rect 28140 9436 28196 9492
rect 28140 9100 28196 9156
rect 28140 8428 28196 8484
rect 29820 13916 29876 13972
rect 29484 13692 29540 13748
rect 29372 13132 29428 13188
rect 29372 12796 29428 12852
rect 29148 12178 29204 12180
rect 29148 12126 29150 12178
rect 29150 12126 29202 12178
rect 29202 12126 29204 12178
rect 29148 12124 29204 12126
rect 29260 12684 29316 12740
rect 29260 12460 29316 12516
rect 28476 10332 28532 10388
rect 29596 12908 29652 12964
rect 29932 15596 29988 15652
rect 29596 12124 29652 12180
rect 29484 10610 29540 10612
rect 29484 10558 29486 10610
rect 29486 10558 29538 10610
rect 29538 10558 29540 10610
rect 29484 10556 29540 10558
rect 28364 9436 28420 9492
rect 28476 8764 28532 8820
rect 28476 8428 28532 8484
rect 28812 7980 28868 8036
rect 26460 7474 26516 7476
rect 26460 7422 26462 7474
rect 26462 7422 26514 7474
rect 26514 7422 26516 7474
rect 26460 7420 26516 7422
rect 25788 6972 25844 7028
rect 25452 6076 25508 6132
rect 26124 6636 26180 6692
rect 26908 7474 26964 7476
rect 26908 7422 26910 7474
rect 26910 7422 26962 7474
rect 26962 7422 26964 7474
rect 26908 7420 26964 7422
rect 27468 7474 27524 7476
rect 27468 7422 27470 7474
rect 27470 7422 27522 7474
rect 27522 7422 27524 7474
rect 27468 7420 27524 7422
rect 26908 6972 26964 7028
rect 26460 6636 26516 6692
rect 26796 6636 26852 6692
rect 26348 6524 26404 6580
rect 25788 5906 25844 5908
rect 25788 5854 25790 5906
rect 25790 5854 25842 5906
rect 25842 5854 25844 5906
rect 25788 5852 25844 5854
rect 24556 5794 24612 5796
rect 24556 5742 24558 5794
rect 24558 5742 24610 5794
rect 24610 5742 24612 5794
rect 24556 5740 24612 5742
rect 26012 5794 26068 5796
rect 26012 5742 26014 5794
rect 26014 5742 26066 5794
rect 26066 5742 26068 5794
rect 26012 5740 26068 5742
rect 27804 6578 27860 6580
rect 27804 6526 27806 6578
rect 27806 6526 27858 6578
rect 27858 6526 27860 6578
rect 27804 6524 27860 6526
rect 30156 13692 30212 13748
rect 30828 21308 30884 21364
rect 31052 22652 31108 22708
rect 30940 20972 30996 21028
rect 32172 25282 32228 25284
rect 32172 25230 32174 25282
rect 32174 25230 32226 25282
rect 32226 25230 32228 25282
rect 32172 25228 32228 25230
rect 31388 23324 31444 23380
rect 31500 21532 31556 21588
rect 30940 20636 30996 20692
rect 30828 19234 30884 19236
rect 30828 19182 30830 19234
rect 30830 19182 30882 19234
rect 30882 19182 30884 19234
rect 30828 19180 30884 19182
rect 31164 20188 31220 20244
rect 31276 20636 31332 20692
rect 31164 19740 31220 19796
rect 30940 18508 30996 18564
rect 31052 18172 31108 18228
rect 30940 17442 30996 17444
rect 30940 17390 30942 17442
rect 30942 17390 30994 17442
rect 30994 17390 30996 17442
rect 30940 17388 30996 17390
rect 31164 17388 31220 17444
rect 30940 16716 30996 16772
rect 30492 16604 30548 16660
rect 30940 15708 30996 15764
rect 31276 16716 31332 16772
rect 31500 20690 31556 20692
rect 31500 20638 31502 20690
rect 31502 20638 31554 20690
rect 31554 20638 31556 20690
rect 31500 20636 31556 20638
rect 32508 27020 32564 27076
rect 32956 27132 33012 27188
rect 33180 27020 33236 27076
rect 33180 26348 33236 26404
rect 32284 24722 32340 24724
rect 32284 24670 32286 24722
rect 32286 24670 32338 24722
rect 32338 24670 32340 24722
rect 32284 24668 32340 24670
rect 31836 24556 31892 24612
rect 31948 24108 32004 24164
rect 32732 25394 32788 25396
rect 32732 25342 32734 25394
rect 32734 25342 32786 25394
rect 32786 25342 32788 25394
rect 32732 25340 32788 25342
rect 32620 25282 32676 25284
rect 32620 25230 32622 25282
rect 32622 25230 32674 25282
rect 32674 25230 32676 25282
rect 32620 25228 32676 25230
rect 32508 24444 32564 24500
rect 32172 23714 32228 23716
rect 32172 23662 32174 23714
rect 32174 23662 32226 23714
rect 32226 23662 32228 23714
rect 32172 23660 32228 23662
rect 31724 22988 31780 23044
rect 31836 22876 31892 22932
rect 31836 22652 31892 22708
rect 31724 21980 31780 22036
rect 32396 23660 32452 23716
rect 32620 24050 32676 24052
rect 32620 23998 32622 24050
rect 32622 23998 32674 24050
rect 32674 23998 32676 24050
rect 32620 23996 32676 23998
rect 33180 23938 33236 23940
rect 33180 23886 33182 23938
rect 33182 23886 33234 23938
rect 33234 23886 33236 23938
rect 33180 23884 33236 23886
rect 33628 28476 33684 28532
rect 33516 27356 33572 27412
rect 34076 31778 34132 31780
rect 34076 31726 34078 31778
rect 34078 31726 34130 31778
rect 34130 31726 34132 31778
rect 34076 31724 34132 31726
rect 33852 31388 33908 31444
rect 34524 31388 34580 31444
rect 36316 33292 36372 33348
rect 37324 37154 37380 37156
rect 37324 37102 37326 37154
rect 37326 37102 37378 37154
rect 37378 37102 37380 37154
rect 37324 37100 37380 37102
rect 37436 36652 37492 36708
rect 39228 35586 39284 35588
rect 39228 35534 39230 35586
rect 39230 35534 39282 35586
rect 39282 35534 39284 35586
rect 39228 35532 39284 35534
rect 38220 35084 38276 35140
rect 37100 34802 37156 34804
rect 37100 34750 37102 34802
rect 37102 34750 37154 34802
rect 37154 34750 37156 34802
rect 37100 34748 37156 34750
rect 37884 34690 37940 34692
rect 37884 34638 37886 34690
rect 37886 34638 37938 34690
rect 37938 34638 37940 34690
rect 37884 34636 37940 34638
rect 38220 34914 38276 34916
rect 38220 34862 38222 34914
rect 38222 34862 38274 34914
rect 38274 34862 38276 34914
rect 38220 34860 38276 34862
rect 38892 35084 38948 35140
rect 38556 34188 38612 34244
rect 38332 34130 38388 34132
rect 38332 34078 38334 34130
rect 38334 34078 38386 34130
rect 38386 34078 38388 34130
rect 38332 34076 38388 34078
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34076 29484 34132 29540
rect 33964 29314 34020 29316
rect 33964 29262 33966 29314
rect 33966 29262 34018 29314
rect 34018 29262 34020 29314
rect 33964 29260 34020 29262
rect 33964 28476 34020 28532
rect 33852 27356 33908 27412
rect 33852 27132 33908 27188
rect 33516 26684 33572 26740
rect 34524 29538 34580 29540
rect 34524 29486 34526 29538
rect 34526 29486 34578 29538
rect 34578 29486 34580 29538
rect 34524 29484 34580 29486
rect 35532 30210 35588 30212
rect 35532 30158 35534 30210
rect 35534 30158 35586 30210
rect 35586 30158 35588 30210
rect 35532 30156 35588 30158
rect 36316 30044 36372 30100
rect 36428 32620 36484 32676
rect 35980 29596 36036 29652
rect 34188 28924 34244 28980
rect 34524 28530 34580 28532
rect 34524 28478 34526 28530
rect 34526 28478 34578 28530
rect 34578 28478 34580 28530
rect 34524 28476 34580 28478
rect 34860 28028 34916 28084
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 39004 34412 39060 34468
rect 37436 30940 37492 30996
rect 36428 29036 36484 29092
rect 36764 29650 36820 29652
rect 36764 29598 36766 29650
rect 36766 29598 36818 29650
rect 36818 29598 36820 29650
rect 36764 29596 36820 29598
rect 36204 28812 36260 28868
rect 36092 28754 36148 28756
rect 36092 28702 36094 28754
rect 36094 28702 36146 28754
rect 36146 28702 36148 28754
rect 36092 28700 36148 28702
rect 35196 28476 35252 28532
rect 34188 27356 34244 27412
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 33516 26348 33572 26404
rect 32620 23324 32676 23380
rect 35308 26348 35364 26404
rect 34188 24444 34244 24500
rect 34412 26178 34468 26180
rect 34412 26126 34414 26178
rect 34414 26126 34466 26178
rect 34466 26126 34468 26178
rect 34412 26124 34468 26126
rect 33852 24050 33908 24052
rect 33852 23998 33854 24050
rect 33854 23998 33906 24050
rect 33906 23998 33908 24050
rect 33852 23996 33908 23998
rect 32508 22876 32564 22932
rect 32732 22204 32788 22260
rect 32172 21756 32228 21812
rect 32284 21698 32340 21700
rect 32284 21646 32286 21698
rect 32286 21646 32338 21698
rect 32338 21646 32340 21698
rect 32284 21644 32340 21646
rect 31724 21362 31780 21364
rect 31724 21310 31726 21362
rect 31726 21310 31778 21362
rect 31778 21310 31780 21362
rect 31724 21308 31780 21310
rect 32172 21308 32228 21364
rect 32284 20972 32340 21028
rect 31948 20914 32004 20916
rect 31948 20862 31950 20914
rect 31950 20862 32002 20914
rect 32002 20862 32004 20914
rect 31948 20860 32004 20862
rect 32396 20748 32452 20804
rect 31836 20636 31892 20692
rect 32284 20690 32340 20692
rect 32284 20638 32286 20690
rect 32286 20638 32338 20690
rect 32338 20638 32340 20690
rect 32284 20636 32340 20638
rect 31724 20300 31780 20356
rect 32172 20130 32228 20132
rect 32172 20078 32174 20130
rect 32174 20078 32226 20130
rect 32226 20078 32228 20130
rect 32172 20076 32228 20078
rect 31948 19122 32004 19124
rect 31948 19070 31950 19122
rect 31950 19070 32002 19122
rect 32002 19070 32004 19122
rect 31948 19068 32004 19070
rect 31948 18450 32004 18452
rect 31948 18398 31950 18450
rect 31950 18398 32002 18450
rect 32002 18398 32004 18450
rect 31948 18396 32004 18398
rect 31612 17836 31668 17892
rect 31724 17442 31780 17444
rect 31724 17390 31726 17442
rect 31726 17390 31778 17442
rect 31778 17390 31780 17442
rect 31724 17388 31780 17390
rect 32172 17052 32228 17108
rect 31164 15932 31220 15988
rect 30492 14924 30548 14980
rect 31276 15596 31332 15652
rect 30380 14028 30436 14084
rect 30940 14588 30996 14644
rect 31052 14418 31108 14420
rect 31052 14366 31054 14418
rect 31054 14366 31106 14418
rect 31106 14366 31108 14418
rect 31052 14364 31108 14366
rect 30492 13692 30548 13748
rect 30380 12684 30436 12740
rect 29820 12012 29876 12068
rect 29932 11676 29988 11732
rect 29372 9324 29428 9380
rect 29484 9548 29540 9604
rect 29148 9042 29204 9044
rect 29148 8990 29150 9042
rect 29150 8990 29202 9042
rect 29202 8990 29204 9042
rect 29148 8988 29204 8990
rect 29260 8764 29316 8820
rect 30268 11452 30324 11508
rect 30604 13356 30660 13412
rect 30940 14028 30996 14084
rect 30716 13132 30772 13188
rect 30716 12962 30772 12964
rect 30716 12910 30718 12962
rect 30718 12910 30770 12962
rect 30770 12910 30772 12962
rect 30716 12908 30772 12910
rect 30604 11394 30660 11396
rect 30604 11342 30606 11394
rect 30606 11342 30658 11394
rect 30658 11342 30660 11394
rect 30604 11340 30660 11342
rect 30828 11340 30884 11396
rect 30044 9212 30100 9268
rect 31164 13580 31220 13636
rect 31052 12236 31108 12292
rect 31388 14530 31444 14532
rect 31388 14478 31390 14530
rect 31390 14478 31442 14530
rect 31442 14478 31444 14530
rect 31388 14476 31444 14478
rect 31948 15260 32004 15316
rect 31500 14418 31556 14420
rect 31500 14366 31502 14418
rect 31502 14366 31554 14418
rect 31554 14366 31556 14418
rect 31500 14364 31556 14366
rect 31612 13580 31668 13636
rect 31948 14476 32004 14532
rect 31500 12290 31556 12292
rect 31500 12238 31502 12290
rect 31502 12238 31554 12290
rect 31554 12238 31556 12290
rect 31500 12236 31556 12238
rect 31612 12012 31668 12068
rect 31724 11676 31780 11732
rect 31948 12012 32004 12068
rect 31948 11676 32004 11732
rect 31052 10610 31108 10612
rect 31052 10558 31054 10610
rect 31054 10558 31106 10610
rect 31106 10558 31108 10610
rect 31052 10556 31108 10558
rect 30716 9548 30772 9604
rect 30828 10220 30884 10276
rect 29708 8316 29764 8372
rect 30380 9212 30436 9268
rect 30716 8988 30772 9044
rect 29932 8034 29988 8036
rect 29932 7982 29934 8034
rect 29934 7982 29986 8034
rect 29986 7982 29988 8034
rect 29932 7980 29988 7982
rect 29708 7586 29764 7588
rect 29708 7534 29710 7586
rect 29710 7534 29762 7586
rect 29762 7534 29764 7586
rect 29708 7532 29764 7534
rect 31052 9884 31108 9940
rect 31388 9826 31444 9828
rect 31388 9774 31390 9826
rect 31390 9774 31442 9826
rect 31442 9774 31444 9826
rect 31388 9772 31444 9774
rect 31836 9884 31892 9940
rect 31052 8540 31108 8596
rect 30940 7644 30996 7700
rect 28364 6690 28420 6692
rect 28364 6638 28366 6690
rect 28366 6638 28418 6690
rect 28418 6638 28420 6690
rect 28364 6636 28420 6638
rect 29148 6690 29204 6692
rect 29148 6638 29150 6690
rect 29150 6638 29202 6690
rect 29202 6638 29204 6690
rect 29148 6636 29204 6638
rect 29260 6524 29316 6580
rect 28028 6466 28084 6468
rect 28028 6414 28030 6466
rect 28030 6414 28082 6466
rect 28082 6414 28084 6466
rect 28028 6412 28084 6414
rect 28252 6018 28308 6020
rect 28252 5966 28254 6018
rect 28254 5966 28306 6018
rect 28306 5966 28308 6018
rect 28252 5964 28308 5966
rect 26684 5794 26740 5796
rect 26684 5742 26686 5794
rect 26686 5742 26738 5794
rect 26738 5742 26740 5794
rect 26684 5740 26740 5742
rect 25228 5628 25284 5684
rect 23212 4956 23268 5012
rect 22092 3724 22148 3780
rect 21420 3554 21476 3556
rect 21420 3502 21422 3554
rect 21422 3502 21474 3554
rect 21474 3502 21476 3554
rect 21420 3500 21476 3502
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 24780 4956 24836 5012
rect 24668 4226 24724 4228
rect 24668 4174 24670 4226
rect 24670 4174 24722 4226
rect 24722 4174 24724 4226
rect 24668 4172 24724 4174
rect 24556 3778 24612 3780
rect 24556 3726 24558 3778
rect 24558 3726 24610 3778
rect 24610 3726 24612 3778
rect 24556 3724 24612 3726
rect 27580 5122 27636 5124
rect 27580 5070 27582 5122
rect 27582 5070 27634 5122
rect 27634 5070 27636 5122
rect 27580 5068 27636 5070
rect 28812 5682 28868 5684
rect 28812 5630 28814 5682
rect 28814 5630 28866 5682
rect 28866 5630 28868 5682
rect 28812 5628 28868 5630
rect 28364 5180 28420 5236
rect 25228 4732 25284 4788
rect 24892 4396 24948 4452
rect 26236 4450 26292 4452
rect 26236 4398 26238 4450
rect 26238 4398 26290 4450
rect 26290 4398 26292 4450
rect 26236 4396 26292 4398
rect 25900 4284 25956 4340
rect 26908 4338 26964 4340
rect 26908 4286 26910 4338
rect 26910 4286 26962 4338
rect 26962 4286 26964 4338
rect 26908 4284 26964 4286
rect 25676 4226 25732 4228
rect 25676 4174 25678 4226
rect 25678 4174 25730 4226
rect 25730 4174 25732 4226
rect 25676 4172 25732 4174
rect 25340 4114 25396 4116
rect 25340 4062 25342 4114
rect 25342 4062 25394 4114
rect 25394 4062 25396 4114
rect 25340 4060 25396 4062
rect 26684 4060 26740 4116
rect 25228 3388 25284 3444
rect 27916 4114 27972 4116
rect 27916 4062 27918 4114
rect 27918 4062 27970 4114
rect 27970 4062 27972 4114
rect 27916 4060 27972 4062
rect 27804 3612 27860 3668
rect 28588 5122 28644 5124
rect 28588 5070 28590 5122
rect 28590 5070 28642 5122
rect 28642 5070 28644 5122
rect 28588 5068 28644 5070
rect 28364 4172 28420 4228
rect 28924 4060 28980 4116
rect 29260 5122 29316 5124
rect 29260 5070 29262 5122
rect 29262 5070 29314 5122
rect 29314 5070 29316 5122
rect 29260 5068 29316 5070
rect 32172 16658 32228 16660
rect 32172 16606 32174 16658
rect 32174 16606 32226 16658
rect 32226 16606 32228 16658
rect 32172 16604 32228 16606
rect 32508 21644 32564 21700
rect 32620 20690 32676 20692
rect 32620 20638 32622 20690
rect 32622 20638 32674 20690
rect 32674 20638 32676 20690
rect 32620 20636 32676 20638
rect 32396 20130 32452 20132
rect 32396 20078 32398 20130
rect 32398 20078 32450 20130
rect 32450 20078 32452 20130
rect 32396 20076 32452 20078
rect 32508 18674 32564 18676
rect 32508 18622 32510 18674
rect 32510 18622 32562 18674
rect 32562 18622 32564 18674
rect 32508 18620 32564 18622
rect 33068 21980 33124 22036
rect 33292 23324 33348 23380
rect 32844 20972 32900 21028
rect 32844 20524 32900 20580
rect 32844 20076 32900 20132
rect 32284 15596 32340 15652
rect 32844 19628 32900 19684
rect 32284 15314 32340 15316
rect 32284 15262 32286 15314
rect 32286 15262 32338 15314
rect 32338 15262 32340 15314
rect 32284 15260 32340 15262
rect 32732 17836 32788 17892
rect 32620 15596 32676 15652
rect 33740 22258 33796 22260
rect 33740 22206 33742 22258
rect 33742 22206 33794 22258
rect 33794 22206 33796 22258
rect 33740 22204 33796 22206
rect 33292 20972 33348 21028
rect 33068 19852 33124 19908
rect 33068 19068 33124 19124
rect 33068 18620 33124 18676
rect 33516 20860 33572 20916
rect 33404 20802 33460 20804
rect 33404 20750 33406 20802
rect 33406 20750 33458 20802
rect 33458 20750 33460 20802
rect 33404 20748 33460 20750
rect 33516 20076 33572 20132
rect 33740 20802 33796 20804
rect 33740 20750 33742 20802
rect 33742 20750 33794 20802
rect 33794 20750 33796 20802
rect 33740 20748 33796 20750
rect 34076 23378 34132 23380
rect 34076 23326 34078 23378
rect 34078 23326 34130 23378
rect 34130 23326 34132 23378
rect 34076 23324 34132 23326
rect 33964 22370 34020 22372
rect 33964 22318 33966 22370
rect 33966 22318 34018 22370
rect 34018 22318 34020 22370
rect 33964 22316 34020 22318
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34524 24668 34580 24724
rect 34748 24444 34804 24500
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34412 22764 34468 22820
rect 34076 21756 34132 21812
rect 34860 22204 34916 22260
rect 34412 21756 34468 21812
rect 34524 21586 34580 21588
rect 34524 21534 34526 21586
rect 34526 21534 34578 21586
rect 34578 21534 34580 21586
rect 34524 21532 34580 21534
rect 34188 21026 34244 21028
rect 34188 20974 34190 21026
rect 34190 20974 34242 21026
rect 34242 20974 34244 21026
rect 34188 20972 34244 20974
rect 34636 20748 34692 20804
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35756 25452 35812 25508
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34972 20748 35028 20804
rect 33852 20188 33908 20244
rect 34524 20524 34580 20580
rect 33852 19964 33908 20020
rect 34076 19964 34132 20020
rect 34188 19852 34244 19908
rect 33964 18396 34020 18452
rect 33068 17276 33124 17332
rect 33516 17276 33572 17332
rect 33516 16940 33572 16996
rect 33740 16994 33796 16996
rect 33740 16942 33742 16994
rect 33742 16942 33794 16994
rect 33794 16942 33796 16994
rect 33740 16940 33796 16942
rect 34860 20076 34916 20132
rect 34412 20018 34468 20020
rect 34412 19966 34414 20018
rect 34414 19966 34466 20018
rect 34466 19966 34468 20018
rect 34412 19964 34468 19966
rect 34524 17724 34580 17780
rect 34748 17778 34804 17780
rect 34748 17726 34750 17778
rect 34750 17726 34802 17778
rect 34802 17726 34804 17778
rect 34748 17724 34804 17726
rect 34076 17052 34132 17108
rect 34300 16994 34356 16996
rect 34300 16942 34302 16994
rect 34302 16942 34354 16994
rect 34354 16942 34356 16994
rect 34300 16940 34356 16942
rect 34636 17164 34692 17220
rect 36988 29260 37044 29316
rect 36988 27132 37044 27188
rect 37100 28700 37156 28756
rect 36540 24722 36596 24724
rect 36540 24670 36542 24722
rect 36542 24670 36594 24722
rect 36594 24670 36596 24722
rect 36540 24668 36596 24670
rect 36428 24050 36484 24052
rect 36428 23998 36430 24050
rect 36430 23998 36482 24050
rect 36482 23998 36484 24050
rect 36428 23996 36484 23998
rect 36988 26348 37044 26404
rect 38108 30210 38164 30212
rect 38108 30158 38110 30210
rect 38110 30158 38162 30210
rect 38162 30158 38164 30210
rect 38108 30156 38164 30158
rect 37436 28812 37492 28868
rect 38556 32562 38612 32564
rect 38556 32510 38558 32562
rect 38558 32510 38610 32562
rect 38610 32510 38612 32562
rect 38556 32508 38612 32510
rect 38668 30994 38724 30996
rect 38668 30942 38670 30994
rect 38670 30942 38722 30994
rect 38722 30942 38724 30994
rect 38668 30940 38724 30942
rect 38668 30098 38724 30100
rect 38668 30046 38670 30098
rect 38670 30046 38722 30098
rect 38722 30046 38724 30098
rect 38668 30044 38724 30046
rect 40012 40908 40068 40964
rect 40124 41020 40180 41076
rect 40012 40514 40068 40516
rect 40012 40462 40014 40514
rect 40014 40462 40066 40514
rect 40066 40462 40068 40514
rect 40012 40460 40068 40462
rect 39340 34300 39396 34356
rect 40684 40908 40740 40964
rect 40684 40460 40740 40516
rect 40012 38780 40068 38836
rect 39788 37772 39844 37828
rect 39788 37212 39844 37268
rect 39900 37938 39956 37940
rect 39900 37886 39902 37938
rect 39902 37886 39954 37938
rect 39954 37886 39956 37938
rect 39900 37884 39956 37886
rect 39900 37100 39956 37156
rect 40460 37266 40516 37268
rect 40460 37214 40462 37266
rect 40462 37214 40514 37266
rect 40514 37214 40516 37266
rect 40460 37212 40516 37214
rect 39788 36652 39844 36708
rect 40572 35532 40628 35588
rect 40572 34914 40628 34916
rect 40572 34862 40574 34914
rect 40574 34862 40626 34914
rect 40626 34862 40628 34914
rect 40572 34860 40628 34862
rect 40012 33404 40068 33460
rect 39452 32508 39508 32564
rect 39452 31948 39508 32004
rect 40124 32508 40180 32564
rect 39564 31612 39620 31668
rect 39004 29820 39060 29876
rect 39228 30156 39284 30212
rect 38332 29148 38388 29204
rect 38220 28812 38276 28868
rect 38780 28812 38836 28868
rect 38668 28588 38724 28644
rect 38556 28140 38612 28196
rect 37996 27916 38052 27972
rect 37660 27468 37716 27524
rect 37212 26962 37268 26964
rect 37212 26910 37214 26962
rect 37214 26910 37266 26962
rect 37266 26910 37268 26962
rect 37212 26908 37268 26910
rect 36652 23996 36708 24052
rect 36988 24108 37044 24164
rect 36428 23492 36484 23548
rect 36764 22876 36820 22932
rect 36204 22316 36260 22372
rect 35756 21586 35812 21588
rect 35756 21534 35758 21586
rect 35758 21534 35810 21586
rect 35810 21534 35812 21586
rect 35756 21532 35812 21534
rect 35644 21308 35700 21364
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35308 19010 35364 19012
rect 35308 18958 35310 19010
rect 35310 18958 35362 19010
rect 35362 18958 35364 19010
rect 35308 18956 35364 18958
rect 34972 18844 35028 18900
rect 35420 18844 35476 18900
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35084 17836 35140 17892
rect 35420 17836 35476 17892
rect 35756 18956 35812 19012
rect 36092 21868 36148 21924
rect 36316 21756 36372 21812
rect 36204 19740 36260 19796
rect 35868 18844 35924 18900
rect 36540 19628 36596 19684
rect 36428 19234 36484 19236
rect 36428 19182 36430 19234
rect 36430 19182 36482 19234
rect 36482 19182 36484 19234
rect 36428 19180 36484 19182
rect 35980 18508 36036 18564
rect 36652 18396 36708 18452
rect 36428 18284 36484 18340
rect 36428 17948 36484 18004
rect 35756 17500 35812 17556
rect 34748 16940 34804 16996
rect 33516 16604 33572 16660
rect 33180 15874 33236 15876
rect 33180 15822 33182 15874
rect 33182 15822 33234 15874
rect 33234 15822 33236 15874
rect 33180 15820 33236 15822
rect 33180 15596 33236 15652
rect 33404 15314 33460 15316
rect 33404 15262 33406 15314
rect 33406 15262 33458 15314
rect 33458 15262 33460 15314
rect 33404 15260 33460 15262
rect 32284 14476 32340 14532
rect 32732 13692 32788 13748
rect 34076 15148 34132 15204
rect 33964 14924 34020 14980
rect 33404 14530 33460 14532
rect 33404 14478 33406 14530
rect 33406 14478 33458 14530
rect 33458 14478 33460 14530
rect 33404 14476 33460 14478
rect 33740 14812 33796 14868
rect 33180 13634 33236 13636
rect 33180 13582 33182 13634
rect 33182 13582 33234 13634
rect 33234 13582 33236 13634
rect 33180 13580 33236 13582
rect 33628 13580 33684 13636
rect 33292 13468 33348 13524
rect 33180 13074 33236 13076
rect 33180 13022 33182 13074
rect 33182 13022 33234 13074
rect 33234 13022 33236 13074
rect 33180 13020 33236 13022
rect 32620 12738 32676 12740
rect 32620 12686 32622 12738
rect 32622 12686 32674 12738
rect 32674 12686 32676 12738
rect 32620 12684 32676 12686
rect 33292 12348 33348 12404
rect 33516 12908 33572 12964
rect 32060 9660 32116 9716
rect 32396 12236 32452 12292
rect 33068 12236 33124 12292
rect 32508 12178 32564 12180
rect 32508 12126 32510 12178
rect 32510 12126 32562 12178
rect 32562 12126 32564 12178
rect 32508 12124 32564 12126
rect 33964 14418 34020 14420
rect 33964 14366 33966 14418
rect 33966 14366 34018 14418
rect 34018 14366 34020 14418
rect 33964 14364 34020 14366
rect 34860 16770 34916 16772
rect 34860 16718 34862 16770
rect 34862 16718 34914 16770
rect 34914 16718 34916 16770
rect 34860 16716 34916 16718
rect 34300 15986 34356 15988
rect 34300 15934 34302 15986
rect 34302 15934 34354 15986
rect 34354 15934 34356 15986
rect 34300 15932 34356 15934
rect 34636 15314 34692 15316
rect 34636 15262 34638 15314
rect 34638 15262 34690 15314
rect 34690 15262 34692 15314
rect 34636 15260 34692 15262
rect 35756 16770 35812 16772
rect 35756 16718 35758 16770
rect 35758 16718 35810 16770
rect 35810 16718 35812 16770
rect 35756 16716 35812 16718
rect 34972 14812 35028 14868
rect 35532 16604 35588 16660
rect 34860 14700 34916 14756
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35420 15596 35476 15652
rect 35980 17164 36036 17220
rect 35980 16940 36036 16996
rect 38444 27186 38500 27188
rect 38444 27134 38446 27186
rect 38446 27134 38498 27186
rect 38498 27134 38500 27186
rect 38444 27132 38500 27134
rect 37324 26402 37380 26404
rect 37324 26350 37326 26402
rect 37326 26350 37378 26402
rect 37378 26350 37380 26402
rect 37324 26348 37380 26350
rect 37436 24668 37492 24724
rect 37884 24780 37940 24836
rect 37548 23772 37604 23828
rect 37324 22876 37380 22932
rect 40236 31612 40292 31668
rect 40908 45218 40964 45220
rect 40908 45166 40910 45218
rect 40910 45166 40962 45218
rect 40962 45166 40964 45218
rect 40908 45164 40964 45166
rect 41132 44044 41188 44100
rect 41020 41970 41076 41972
rect 41020 41918 41022 41970
rect 41022 41918 41074 41970
rect 41074 41918 41076 41970
rect 41020 41916 41076 41918
rect 42364 47234 42420 47236
rect 42364 47182 42366 47234
rect 42366 47182 42418 47234
rect 42418 47182 42420 47234
rect 42364 47180 42420 47182
rect 41804 46956 41860 47012
rect 41468 44994 41524 44996
rect 41468 44942 41470 44994
rect 41470 44942 41522 44994
rect 41522 44942 41524 44994
rect 41468 44940 41524 44942
rect 43036 44940 43092 44996
rect 41468 44156 41524 44212
rect 41804 44044 41860 44100
rect 43372 44210 43428 44212
rect 43372 44158 43374 44210
rect 43374 44158 43426 44210
rect 43426 44158 43428 44210
rect 43372 44156 43428 44158
rect 45164 44156 45220 44212
rect 42028 43314 42084 43316
rect 42028 43262 42030 43314
rect 42030 43262 42082 43314
rect 42082 43262 42084 43314
rect 42028 43260 42084 43262
rect 41692 41916 41748 41972
rect 42924 43260 42980 43316
rect 42924 42140 42980 42196
rect 42364 41970 42420 41972
rect 42364 41918 42366 41970
rect 42366 41918 42418 41970
rect 42418 41918 42420 41970
rect 42364 41916 42420 41918
rect 41804 40962 41860 40964
rect 41804 40910 41806 40962
rect 41806 40910 41858 40962
rect 41858 40910 41860 40962
rect 41804 40908 41860 40910
rect 41356 40348 41412 40404
rect 42364 40348 42420 40404
rect 41468 37884 41524 37940
rect 42252 37436 42308 37492
rect 41916 37100 41972 37156
rect 42812 41074 42868 41076
rect 42812 41022 42814 41074
rect 42814 41022 42866 41074
rect 42866 41022 42868 41074
rect 42812 41020 42868 41022
rect 42588 40908 42644 40964
rect 42812 40348 42868 40404
rect 41020 34354 41076 34356
rect 41020 34302 41022 34354
rect 41022 34302 41074 34354
rect 41074 34302 41076 34354
rect 41020 34300 41076 34302
rect 41244 33516 41300 33572
rect 41580 33906 41636 33908
rect 41580 33854 41582 33906
rect 41582 33854 41634 33906
rect 41634 33854 41636 33906
rect 41580 33852 41636 33854
rect 41356 32620 41412 32676
rect 41580 32732 41636 32788
rect 40908 32562 40964 32564
rect 40908 32510 40910 32562
rect 40910 32510 40962 32562
rect 40962 32510 40964 32562
rect 40908 32508 40964 32510
rect 40572 31778 40628 31780
rect 40572 31726 40574 31778
rect 40574 31726 40626 31778
rect 40626 31726 40628 31778
rect 40572 31724 40628 31726
rect 40348 31164 40404 31220
rect 40348 30882 40404 30884
rect 40348 30830 40350 30882
rect 40350 30830 40402 30882
rect 40402 30830 40404 30882
rect 40348 30828 40404 30830
rect 39788 29426 39844 29428
rect 39788 29374 39790 29426
rect 39790 29374 39842 29426
rect 39842 29374 39844 29426
rect 39788 29372 39844 29374
rect 39116 28700 39172 28756
rect 38892 28642 38948 28644
rect 38892 28590 38894 28642
rect 38894 28590 38946 28642
rect 38946 28590 38948 28642
rect 38892 28588 38948 28590
rect 39340 28476 39396 28532
rect 40236 28476 40292 28532
rect 39228 28028 39284 28084
rect 38892 27580 38948 27636
rect 39564 27580 39620 27636
rect 38892 27244 38948 27300
rect 39452 27074 39508 27076
rect 39452 27022 39454 27074
rect 39454 27022 39506 27074
rect 39506 27022 39508 27074
rect 39452 27020 39508 27022
rect 38556 24834 38612 24836
rect 38556 24782 38558 24834
rect 38558 24782 38610 24834
rect 38610 24782 38612 24834
rect 38556 24780 38612 24782
rect 38332 24220 38388 24276
rect 37996 23826 38052 23828
rect 37996 23774 37998 23826
rect 37998 23774 38050 23826
rect 38050 23774 38052 23826
rect 37996 23772 38052 23774
rect 37884 22988 37940 23044
rect 38444 24332 38500 24388
rect 38780 24722 38836 24724
rect 38780 24670 38782 24722
rect 38782 24670 38834 24722
rect 38834 24670 38836 24722
rect 38780 24668 38836 24670
rect 39788 27356 39844 27412
rect 40012 27356 40068 27412
rect 40124 27020 40180 27076
rect 39788 26908 39844 26964
rect 39676 26850 39732 26852
rect 39676 26798 39678 26850
rect 39678 26798 39730 26850
rect 39730 26798 39732 26850
rect 39676 26796 39732 26798
rect 40460 30268 40516 30324
rect 40572 31500 40628 31556
rect 40348 27746 40404 27748
rect 40348 27694 40350 27746
rect 40350 27694 40402 27746
rect 40402 27694 40404 27746
rect 40348 27692 40404 27694
rect 40908 31666 40964 31668
rect 40908 31614 40910 31666
rect 40910 31614 40962 31666
rect 40962 31614 40964 31666
rect 40908 31612 40964 31614
rect 40796 31164 40852 31220
rect 41132 31724 41188 31780
rect 41132 31218 41188 31220
rect 41132 31166 41134 31218
rect 41134 31166 41186 31218
rect 41186 31166 41188 31218
rect 41132 31164 41188 31166
rect 40796 30322 40852 30324
rect 40796 30270 40798 30322
rect 40798 30270 40850 30322
rect 40850 30270 40852 30322
rect 40796 30268 40852 30270
rect 40796 30044 40852 30100
rect 41356 31500 41412 31556
rect 41468 30828 41524 30884
rect 41020 30156 41076 30212
rect 40908 29708 40964 29764
rect 41244 30098 41300 30100
rect 41244 30046 41246 30098
rect 41246 30046 41298 30098
rect 41298 30046 41300 30098
rect 41244 30044 41300 30046
rect 41244 29538 41300 29540
rect 41244 29486 41246 29538
rect 41246 29486 41298 29538
rect 41298 29486 41300 29538
rect 41244 29484 41300 29486
rect 41132 28476 41188 28532
rect 40908 27916 40964 27972
rect 41020 27804 41076 27860
rect 40684 27244 40740 27300
rect 40348 26684 40404 26740
rect 40236 26236 40292 26292
rect 38556 23826 38612 23828
rect 38556 23774 38558 23826
rect 38558 23774 38610 23826
rect 38610 23774 38612 23826
rect 38556 23772 38612 23774
rect 38444 23660 38500 23716
rect 39340 24556 39396 24612
rect 38780 23378 38836 23380
rect 38780 23326 38782 23378
rect 38782 23326 38834 23378
rect 38834 23326 38836 23378
rect 38780 23324 38836 23326
rect 37996 22652 38052 22708
rect 36876 21644 36932 21700
rect 37212 21868 37268 21924
rect 36876 21420 36932 21476
rect 37212 21362 37268 21364
rect 37212 21310 37214 21362
rect 37214 21310 37266 21362
rect 37266 21310 37268 21362
rect 37212 21308 37268 21310
rect 37436 21586 37492 21588
rect 37436 21534 37438 21586
rect 37438 21534 37490 21586
rect 37490 21534 37492 21586
rect 37436 21532 37492 21534
rect 36988 18396 37044 18452
rect 36652 17164 36708 17220
rect 36764 17388 36820 17444
rect 37100 18060 37156 18116
rect 37212 18508 37268 18564
rect 37772 21698 37828 21700
rect 37772 21646 37774 21698
rect 37774 21646 37826 21698
rect 37826 21646 37828 21698
rect 37772 21644 37828 21646
rect 39004 22146 39060 22148
rect 39004 22094 39006 22146
rect 39006 22094 39058 22146
rect 39058 22094 39060 22146
rect 39004 22092 39060 22094
rect 38444 21644 38500 21700
rect 38668 21586 38724 21588
rect 38668 21534 38670 21586
rect 38670 21534 38722 21586
rect 38722 21534 38724 21586
rect 38668 21532 38724 21534
rect 38780 21196 38836 21252
rect 37996 20578 38052 20580
rect 37996 20526 37998 20578
rect 37998 20526 38050 20578
rect 38050 20526 38052 20578
rect 37996 20524 38052 20526
rect 38108 20018 38164 20020
rect 38108 19966 38110 20018
rect 38110 19966 38162 20018
rect 38162 19966 38164 20018
rect 38108 19964 38164 19966
rect 37996 19628 38052 19684
rect 37548 19234 37604 19236
rect 37548 19182 37550 19234
rect 37550 19182 37602 19234
rect 37602 19182 37604 19234
rect 37548 19180 37604 19182
rect 37660 18732 37716 18788
rect 37212 17778 37268 17780
rect 37212 17726 37214 17778
rect 37214 17726 37266 17778
rect 37266 17726 37268 17778
rect 37212 17724 37268 17726
rect 36988 17500 37044 17556
rect 36876 16940 36932 16996
rect 37100 16940 37156 16996
rect 36764 16882 36820 16884
rect 36764 16830 36766 16882
rect 36766 16830 36818 16882
rect 36818 16830 36820 16882
rect 36764 16828 36820 16830
rect 36876 16770 36932 16772
rect 36876 16718 36878 16770
rect 36878 16718 36930 16770
rect 36930 16718 36932 16770
rect 36876 16716 36932 16718
rect 36652 16604 36708 16660
rect 37436 17948 37492 18004
rect 37436 17612 37492 17668
rect 37436 17164 37492 17220
rect 37772 18396 37828 18452
rect 37996 18284 38052 18340
rect 37660 17106 37716 17108
rect 37660 17054 37662 17106
rect 37662 17054 37714 17106
rect 37714 17054 37716 17106
rect 37660 17052 37716 17054
rect 38444 20690 38500 20692
rect 38444 20638 38446 20690
rect 38446 20638 38498 20690
rect 38498 20638 38500 20690
rect 38444 20636 38500 20638
rect 38668 20076 38724 20132
rect 38332 19180 38388 19236
rect 38556 19180 38612 19236
rect 38444 19068 38500 19124
rect 38444 18620 38500 18676
rect 38332 18172 38388 18228
rect 37100 16380 37156 16436
rect 36316 16044 36372 16100
rect 36092 15986 36148 15988
rect 36092 15934 36094 15986
rect 36094 15934 36146 15986
rect 36146 15934 36148 15986
rect 36092 15932 36148 15934
rect 36988 15932 37044 15988
rect 36540 15820 36596 15876
rect 37100 15708 37156 15764
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 14364 35252 14420
rect 34524 13970 34580 13972
rect 34524 13918 34526 13970
rect 34526 13918 34578 13970
rect 34578 13918 34580 13970
rect 34524 13916 34580 13918
rect 34972 13916 35028 13972
rect 34860 13858 34916 13860
rect 34860 13806 34862 13858
rect 34862 13806 34914 13858
rect 34914 13806 34916 13858
rect 34860 13804 34916 13806
rect 34188 13692 34244 13748
rect 33852 13020 33908 13076
rect 33628 12460 33684 12516
rect 32508 11676 32564 11732
rect 34972 12908 35028 12964
rect 34188 12850 34244 12852
rect 34188 12798 34190 12850
rect 34190 12798 34242 12850
rect 34242 12798 34244 12850
rect 34188 12796 34244 12798
rect 34412 12850 34468 12852
rect 34412 12798 34414 12850
rect 34414 12798 34466 12850
rect 34466 12798 34468 12850
rect 34412 12796 34468 12798
rect 34860 12796 34916 12852
rect 35644 14642 35700 14644
rect 35644 14590 35646 14642
rect 35646 14590 35698 14642
rect 35698 14590 35700 14642
rect 35644 14588 35700 14590
rect 35308 13468 35364 13524
rect 36652 15314 36708 15316
rect 36652 15262 36654 15314
rect 36654 15262 36706 15314
rect 36706 15262 36708 15314
rect 36652 15260 36708 15262
rect 37324 16604 37380 16660
rect 37548 15484 37604 15540
rect 37212 15372 37268 15428
rect 37436 15372 37492 15428
rect 37548 15314 37604 15316
rect 37548 15262 37550 15314
rect 37550 15262 37602 15314
rect 37602 15262 37604 15314
rect 37548 15260 37604 15262
rect 36092 14924 36148 14980
rect 36204 14812 36260 14868
rect 36988 14700 37044 14756
rect 35532 13804 35588 13860
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 13074 35252 13076
rect 35196 13022 35198 13074
rect 35198 13022 35250 13074
rect 35250 13022 35252 13074
rect 35196 13020 35252 13022
rect 35980 14476 36036 14532
rect 34524 12684 34580 12740
rect 34076 12460 34132 12516
rect 33068 9996 33124 10052
rect 32844 9714 32900 9716
rect 32844 9662 32846 9714
rect 32846 9662 32898 9714
rect 32898 9662 32900 9714
rect 32844 9660 32900 9662
rect 34412 12460 34468 12516
rect 34300 12178 34356 12180
rect 34300 12126 34302 12178
rect 34302 12126 34354 12178
rect 34354 12126 34356 12178
rect 34300 12124 34356 12126
rect 34524 12178 34580 12180
rect 34524 12126 34526 12178
rect 34526 12126 34578 12178
rect 34578 12126 34580 12178
rect 34524 12124 34580 12126
rect 34860 11900 34916 11956
rect 34636 11564 34692 11620
rect 33852 9772 33908 9828
rect 32620 9602 32676 9604
rect 32620 9550 32622 9602
rect 32622 9550 32674 9602
rect 32674 9550 32676 9602
rect 32620 9548 32676 9550
rect 32284 9436 32340 9492
rect 29820 6412 29876 6468
rect 30044 5180 30100 5236
rect 29596 4956 29652 5012
rect 31052 5964 31108 6020
rect 34076 9660 34132 9716
rect 33404 9042 33460 9044
rect 33404 8990 33406 9042
rect 33406 8990 33458 9042
rect 33458 8990 33460 9042
rect 33404 8988 33460 8990
rect 34300 9436 34356 9492
rect 34524 11004 34580 11060
rect 32284 8876 32340 8932
rect 33068 8930 33124 8932
rect 33068 8878 33070 8930
rect 33070 8878 33122 8930
rect 33122 8878 33124 8930
rect 33068 8876 33124 8878
rect 32172 8316 32228 8372
rect 33292 8428 33348 8484
rect 32508 7698 32564 7700
rect 32508 7646 32510 7698
rect 32510 7646 32562 7698
rect 32562 7646 32564 7698
rect 32508 7644 32564 7646
rect 32060 6300 32116 6356
rect 34076 8428 34132 8484
rect 34412 8428 34468 8484
rect 34636 10892 34692 10948
rect 35196 11900 35252 11956
rect 34972 11564 35028 11620
rect 34636 9602 34692 9604
rect 34636 9550 34638 9602
rect 34638 9550 34690 9602
rect 34690 9550 34692 9602
rect 34636 9548 34692 9550
rect 34860 9996 34916 10052
rect 34748 8258 34804 8260
rect 34748 8206 34750 8258
rect 34750 8206 34802 8258
rect 34802 8206 34804 8258
rect 34748 8204 34804 8206
rect 34076 7586 34132 7588
rect 34076 7534 34078 7586
rect 34078 7534 34130 7586
rect 34130 7534 34132 7586
rect 34076 7532 34132 7534
rect 32508 7420 32564 7476
rect 32620 6690 32676 6692
rect 32620 6638 32622 6690
rect 32622 6638 32674 6690
rect 32674 6638 32676 6690
rect 32620 6636 32676 6638
rect 32172 6076 32228 6132
rect 33516 6412 33572 6468
rect 31948 5852 32004 5908
rect 32508 5906 32564 5908
rect 32508 5854 32510 5906
rect 32510 5854 32562 5906
rect 32562 5854 32564 5906
rect 32508 5852 32564 5854
rect 31724 5628 31780 5684
rect 30828 5122 30884 5124
rect 30828 5070 30830 5122
rect 30830 5070 30882 5122
rect 30882 5070 30884 5122
rect 30828 5068 30884 5070
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35420 11506 35476 11508
rect 35420 11454 35422 11506
rect 35422 11454 35474 11506
rect 35474 11454 35476 11506
rect 35420 11452 35476 11454
rect 35756 13020 35812 13076
rect 35868 12850 35924 12852
rect 35868 12798 35870 12850
rect 35870 12798 35922 12850
rect 35922 12798 35924 12850
rect 35868 12796 35924 12798
rect 35084 10892 35140 10948
rect 35532 10780 35588 10836
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35532 9826 35588 9828
rect 35532 9774 35534 9826
rect 35534 9774 35586 9826
rect 35586 9774 35588 9826
rect 35532 9772 35588 9774
rect 35756 9884 35812 9940
rect 35868 9996 35924 10052
rect 35644 9660 35700 9716
rect 35532 9324 35588 9380
rect 35420 8764 35476 8820
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 8092 35252 8148
rect 34972 7698 35028 7700
rect 34972 7646 34974 7698
rect 34974 7646 35026 7698
rect 35026 7646 35028 7698
rect 34972 7644 35028 7646
rect 35756 8258 35812 8260
rect 35756 8206 35758 8258
rect 35758 8206 35810 8258
rect 35810 8206 35812 8258
rect 35756 8204 35812 8206
rect 35532 7698 35588 7700
rect 35532 7646 35534 7698
rect 35534 7646 35586 7698
rect 35586 7646 35588 7698
rect 35532 7644 35588 7646
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 36092 14364 36148 14420
rect 36316 13692 36372 13748
rect 37436 15148 37492 15204
rect 37212 14028 37268 14084
rect 36540 13634 36596 13636
rect 36540 13582 36542 13634
rect 36542 13582 36594 13634
rect 36594 13582 36596 13634
rect 36540 13580 36596 13582
rect 36316 12572 36372 12628
rect 36428 12796 36484 12852
rect 36092 12348 36148 12404
rect 36092 11954 36148 11956
rect 36092 11902 36094 11954
rect 36094 11902 36146 11954
rect 36146 11902 36148 11954
rect 36092 11900 36148 11902
rect 36092 9884 36148 9940
rect 37212 11394 37268 11396
rect 37212 11342 37214 11394
rect 37214 11342 37266 11394
rect 37266 11342 37268 11394
rect 37212 11340 37268 11342
rect 37324 13746 37380 13748
rect 37324 13694 37326 13746
rect 37326 13694 37378 13746
rect 37378 13694 37380 13746
rect 37324 13692 37380 13694
rect 38108 17612 38164 17668
rect 38668 17948 38724 18004
rect 38556 17612 38612 17668
rect 38220 17106 38276 17108
rect 38220 17054 38222 17106
rect 38222 17054 38274 17106
rect 38274 17054 38276 17106
rect 38220 17052 38276 17054
rect 38444 16716 38500 16772
rect 38220 16604 38276 16660
rect 37996 15484 38052 15540
rect 37884 15314 37940 15316
rect 37884 15262 37886 15314
rect 37886 15262 37938 15314
rect 37938 15262 37940 15314
rect 37884 15260 37940 15262
rect 39788 24108 39844 24164
rect 39452 23884 39508 23940
rect 39676 23548 39732 23604
rect 40908 26796 40964 26852
rect 41580 29484 41636 29540
rect 42476 34690 42532 34692
rect 42476 34638 42478 34690
rect 42478 34638 42530 34690
rect 42530 34638 42532 34690
rect 42476 34636 42532 34638
rect 42476 34300 42532 34356
rect 42140 33964 42196 34020
rect 41916 33516 41972 33572
rect 42028 33292 42084 33348
rect 42364 33292 42420 33348
rect 42028 32732 42084 32788
rect 41804 31948 41860 32004
rect 42140 31164 42196 31220
rect 42700 36316 42756 36372
rect 42700 34242 42756 34244
rect 42700 34190 42702 34242
rect 42702 34190 42754 34242
rect 42754 34190 42756 34242
rect 42700 34188 42756 34190
rect 42700 33740 42756 33796
rect 43820 42140 43876 42196
rect 45724 42194 45780 42196
rect 45724 42142 45726 42194
rect 45726 42142 45778 42194
rect 45778 42142 45780 42194
rect 45724 42140 45780 42142
rect 43484 41020 43540 41076
rect 43148 40348 43204 40404
rect 45052 40402 45108 40404
rect 45052 40350 45054 40402
rect 45054 40350 45106 40402
rect 45106 40350 45108 40402
rect 45052 40348 45108 40350
rect 43484 37436 43540 37492
rect 43148 37378 43204 37380
rect 43148 37326 43150 37378
rect 43150 37326 43202 37378
rect 43202 37326 43204 37378
rect 43148 37324 43204 37326
rect 43372 37266 43428 37268
rect 43372 37214 43374 37266
rect 43374 37214 43426 37266
rect 43426 37214 43428 37266
rect 43372 37212 43428 37214
rect 44044 37324 44100 37380
rect 44156 37212 44212 37268
rect 43708 37100 43764 37156
rect 43260 36316 43316 36372
rect 44156 36370 44212 36372
rect 44156 36318 44158 36370
rect 44158 36318 44210 36370
rect 44210 36318 44212 36370
rect 44156 36316 44212 36318
rect 44828 36316 44884 36372
rect 46508 36316 46564 36372
rect 43036 34802 43092 34804
rect 43036 34750 43038 34802
rect 43038 34750 43090 34802
rect 43090 34750 43092 34802
rect 43036 34748 43092 34750
rect 42924 34636 42980 34692
rect 43036 33740 43092 33796
rect 44156 34690 44212 34692
rect 44156 34638 44158 34690
rect 44158 34638 44210 34690
rect 44210 34638 44212 34690
rect 44156 34636 44212 34638
rect 43932 34188 43988 34244
rect 43260 33628 43316 33684
rect 43036 32786 43092 32788
rect 43036 32734 43038 32786
rect 43038 32734 43090 32786
rect 43090 32734 43092 32786
rect 43036 32732 43092 32734
rect 43372 33346 43428 33348
rect 43372 33294 43374 33346
rect 43374 33294 43426 33346
rect 43426 33294 43428 33346
rect 43372 33292 43428 33294
rect 43148 31836 43204 31892
rect 42700 31554 42756 31556
rect 42700 31502 42702 31554
rect 42702 31502 42754 31554
rect 42754 31502 42756 31554
rect 42700 31500 42756 31502
rect 41916 30268 41972 30324
rect 42364 30044 42420 30100
rect 42476 29820 42532 29876
rect 41916 29708 41972 29764
rect 41580 27916 41636 27972
rect 41468 27132 41524 27188
rect 41244 26908 41300 26964
rect 42700 27692 42756 27748
rect 42364 27468 42420 27524
rect 42700 27186 42756 27188
rect 42700 27134 42702 27186
rect 42702 27134 42754 27186
rect 42754 27134 42756 27186
rect 42700 27132 42756 27134
rect 42252 27074 42308 27076
rect 42252 27022 42254 27074
rect 42254 27022 42306 27074
rect 42306 27022 42308 27074
rect 42252 27020 42308 27022
rect 41916 26684 41972 26740
rect 43036 30380 43092 30436
rect 43596 30380 43652 30436
rect 43148 30268 43204 30324
rect 43036 28028 43092 28084
rect 43036 27356 43092 27412
rect 44156 30210 44212 30212
rect 44156 30158 44158 30210
rect 44158 30158 44210 30210
rect 44210 30158 44212 30210
rect 44156 30156 44212 30158
rect 43932 30098 43988 30100
rect 43932 30046 43934 30098
rect 43934 30046 43986 30098
rect 43986 30046 43988 30098
rect 43932 30044 43988 30046
rect 43372 29372 43428 29428
rect 44044 29932 44100 29988
rect 44044 28140 44100 28196
rect 43596 27916 43652 27972
rect 43484 27468 43540 27524
rect 43372 26908 43428 26964
rect 41468 26124 41524 26180
rect 40796 25900 40852 25956
rect 41132 24722 41188 24724
rect 41132 24670 41134 24722
rect 41134 24670 41186 24722
rect 41186 24670 41188 24722
rect 41132 24668 41188 24670
rect 39900 23884 39956 23940
rect 40124 23154 40180 23156
rect 40124 23102 40126 23154
rect 40126 23102 40178 23154
rect 40178 23102 40180 23154
rect 40124 23100 40180 23102
rect 39452 22146 39508 22148
rect 39452 22094 39454 22146
rect 39454 22094 39506 22146
rect 39506 22094 39508 22146
rect 39452 22092 39508 22094
rect 39788 22092 39844 22148
rect 42028 25228 42084 25284
rect 41356 23212 41412 23268
rect 41020 23154 41076 23156
rect 41020 23102 41022 23154
rect 41022 23102 41074 23154
rect 41074 23102 41076 23154
rect 41020 23100 41076 23102
rect 40460 22092 40516 22148
rect 41132 22092 41188 22148
rect 39452 21698 39508 21700
rect 39452 21646 39454 21698
rect 39454 21646 39506 21698
rect 39506 21646 39508 21698
rect 39452 21644 39508 21646
rect 39116 21532 39172 21588
rect 39340 21474 39396 21476
rect 39340 21422 39342 21474
rect 39342 21422 39394 21474
rect 39394 21422 39396 21474
rect 39340 21420 39396 21422
rect 39228 21362 39284 21364
rect 39228 21310 39230 21362
rect 39230 21310 39282 21362
rect 39282 21310 39284 21362
rect 39228 21308 39284 21310
rect 39004 20076 39060 20132
rect 38892 19964 38948 20020
rect 39452 19794 39508 19796
rect 39452 19742 39454 19794
rect 39454 19742 39506 19794
rect 39506 19742 39508 19794
rect 39452 19740 39508 19742
rect 38892 18620 38948 18676
rect 39228 18450 39284 18452
rect 39228 18398 39230 18450
rect 39230 18398 39282 18450
rect 39282 18398 39284 18450
rect 39228 18396 39284 18398
rect 39004 18060 39060 18116
rect 39004 17666 39060 17668
rect 39004 17614 39006 17666
rect 39006 17614 39058 17666
rect 39058 17614 39060 17666
rect 39004 17612 39060 17614
rect 39340 17612 39396 17668
rect 39228 17276 39284 17332
rect 39228 16940 39284 16996
rect 39452 16994 39508 16996
rect 39452 16942 39454 16994
rect 39454 16942 39506 16994
rect 39506 16942 39508 16994
rect 39452 16940 39508 16942
rect 39340 16828 39396 16884
rect 40124 21698 40180 21700
rect 40124 21646 40126 21698
rect 40126 21646 40178 21698
rect 40178 21646 40180 21698
rect 40124 21644 40180 21646
rect 42028 23884 42084 23940
rect 41692 23212 41748 23268
rect 41916 23436 41972 23492
rect 42140 24668 42196 24724
rect 42028 22428 42084 22484
rect 41468 21644 41524 21700
rect 41804 21644 41860 21700
rect 39676 21196 39732 21252
rect 39676 20524 39732 20580
rect 40348 19234 40404 19236
rect 40348 19182 40350 19234
rect 40350 19182 40402 19234
rect 40402 19182 40404 19234
rect 40348 19180 40404 19182
rect 41020 18956 41076 19012
rect 39676 18450 39732 18452
rect 39676 18398 39678 18450
rect 39678 18398 39730 18450
rect 39730 18398 39732 18450
rect 39676 18396 39732 18398
rect 41020 18562 41076 18564
rect 41020 18510 41022 18562
rect 41022 18510 41074 18562
rect 41074 18510 41076 18562
rect 41020 18508 41076 18510
rect 40908 18450 40964 18452
rect 40908 18398 40910 18450
rect 40910 18398 40962 18450
rect 40962 18398 40964 18450
rect 40908 18396 40964 18398
rect 40012 17948 40068 18004
rect 40796 18284 40852 18340
rect 41468 18284 41524 18340
rect 40012 17276 40068 17332
rect 41132 17666 41188 17668
rect 41132 17614 41134 17666
rect 41134 17614 41186 17666
rect 41186 17614 41188 17666
rect 41132 17612 41188 17614
rect 41020 17276 41076 17332
rect 41356 17164 41412 17220
rect 40908 17106 40964 17108
rect 40908 17054 40910 17106
rect 40910 17054 40962 17106
rect 40962 17054 40964 17106
rect 40908 17052 40964 17054
rect 40572 16940 40628 16996
rect 38780 16492 38836 16548
rect 39340 16492 39396 16548
rect 38556 15708 38612 15764
rect 38780 15484 38836 15540
rect 38332 15202 38388 15204
rect 38332 15150 38334 15202
rect 38334 15150 38386 15202
rect 38386 15150 38388 15202
rect 38332 15148 38388 15150
rect 38892 15202 38948 15204
rect 38892 15150 38894 15202
rect 38894 15150 38946 15202
rect 38946 15150 38948 15202
rect 38892 15148 38948 15150
rect 39788 16658 39844 16660
rect 39788 16606 39790 16658
rect 39790 16606 39842 16658
rect 39842 16606 39844 16658
rect 39788 16604 39844 16606
rect 39900 16492 39956 16548
rect 37884 14924 37940 14980
rect 37436 12796 37492 12852
rect 37548 13580 37604 13636
rect 37996 13074 38052 13076
rect 37996 13022 37998 13074
rect 37998 13022 38050 13074
rect 38050 13022 38052 13074
rect 37996 13020 38052 13022
rect 38556 14588 38612 14644
rect 38444 13916 38500 13972
rect 38220 13746 38276 13748
rect 38220 13694 38222 13746
rect 38222 13694 38274 13746
rect 38274 13694 38276 13746
rect 38220 13692 38276 13694
rect 37884 12796 37940 12852
rect 37548 12124 37604 12180
rect 37324 10722 37380 10724
rect 37324 10670 37326 10722
rect 37326 10670 37378 10722
rect 37378 10670 37380 10722
rect 37324 10668 37380 10670
rect 37772 10610 37828 10612
rect 37772 10558 37774 10610
rect 37774 10558 37826 10610
rect 37826 10558 37828 10610
rect 37772 10556 37828 10558
rect 36988 9996 37044 10052
rect 37212 9996 37268 10052
rect 37212 9548 37268 9604
rect 36428 8652 36484 8708
rect 38668 13634 38724 13636
rect 38668 13582 38670 13634
rect 38670 13582 38722 13634
rect 38722 13582 38724 13634
rect 38668 13580 38724 13582
rect 38668 12796 38724 12852
rect 39228 12402 39284 12404
rect 39228 12350 39230 12402
rect 39230 12350 39282 12402
rect 39282 12350 39284 12402
rect 39228 12348 39284 12350
rect 38780 12066 38836 12068
rect 38780 12014 38782 12066
rect 38782 12014 38834 12066
rect 38834 12014 38836 12066
rect 38780 12012 38836 12014
rect 38108 11394 38164 11396
rect 38108 11342 38110 11394
rect 38110 11342 38162 11394
rect 38162 11342 38164 11394
rect 38108 11340 38164 11342
rect 37996 11116 38052 11172
rect 38108 10834 38164 10836
rect 38108 10782 38110 10834
rect 38110 10782 38162 10834
rect 38162 10782 38164 10834
rect 38108 10780 38164 10782
rect 37996 9996 38052 10052
rect 37212 9100 37268 9156
rect 38780 10722 38836 10724
rect 38780 10670 38782 10722
rect 38782 10670 38834 10722
rect 38834 10670 38836 10722
rect 38780 10668 38836 10670
rect 38108 9602 38164 9604
rect 38108 9550 38110 9602
rect 38110 9550 38162 9602
rect 38162 9550 38164 9602
rect 38108 9548 38164 9550
rect 37324 8876 37380 8932
rect 38444 10444 38500 10500
rect 42812 21644 42868 21700
rect 42364 21586 42420 21588
rect 42364 21534 42366 21586
rect 42366 21534 42418 21586
rect 42418 21534 42420 21586
rect 42364 21532 42420 21534
rect 43036 26290 43092 26292
rect 43036 26238 43038 26290
rect 43038 26238 43090 26290
rect 43090 26238 43092 26290
rect 43036 26236 43092 26238
rect 43036 24668 43092 24724
rect 41804 19346 41860 19348
rect 41804 19294 41806 19346
rect 41806 19294 41858 19346
rect 41858 19294 41860 19346
rect 41804 19292 41860 19294
rect 41916 18284 41972 18340
rect 41916 18060 41972 18116
rect 41916 17612 41972 17668
rect 41580 16716 41636 16772
rect 41356 16156 41412 16212
rect 39564 14812 39620 14868
rect 40796 13916 40852 13972
rect 41132 13970 41188 13972
rect 41132 13918 41134 13970
rect 41134 13918 41186 13970
rect 41186 13918 41188 13970
rect 41132 13916 41188 13918
rect 40124 12012 40180 12068
rect 39340 10892 39396 10948
rect 39452 11116 39508 11172
rect 39116 9938 39172 9940
rect 39116 9886 39118 9938
rect 39118 9886 39170 9938
rect 39170 9886 39172 9938
rect 39116 9884 39172 9886
rect 39004 9660 39060 9716
rect 38108 8876 38164 8932
rect 38108 8652 38164 8708
rect 35196 6466 35252 6468
rect 35196 6414 35198 6466
rect 35198 6414 35250 6466
rect 35250 6414 35252 6466
rect 35196 6412 35252 6414
rect 36092 8092 36148 8148
rect 37660 8204 37716 8260
rect 36092 6690 36148 6692
rect 36092 6638 36094 6690
rect 36094 6638 36146 6690
rect 36146 6638 36148 6690
rect 36092 6636 36148 6638
rect 36316 6578 36372 6580
rect 36316 6526 36318 6578
rect 36318 6526 36370 6578
rect 36370 6526 36372 6578
rect 36316 6524 36372 6526
rect 35980 6412 36036 6468
rect 34076 5906 34132 5908
rect 34076 5854 34078 5906
rect 34078 5854 34130 5906
rect 34130 5854 34132 5906
rect 34076 5852 34132 5854
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34076 5180 34132 5236
rect 34636 5180 34692 5236
rect 33628 5068 33684 5124
rect 35532 5234 35588 5236
rect 35532 5182 35534 5234
rect 35534 5182 35586 5234
rect 35586 5182 35588 5234
rect 35532 5180 35588 5182
rect 35084 5122 35140 5124
rect 35084 5070 35086 5122
rect 35086 5070 35138 5122
rect 35138 5070 35140 5122
rect 35084 5068 35140 5070
rect 31388 4898 31444 4900
rect 31388 4846 31390 4898
rect 31390 4846 31442 4898
rect 31442 4846 31444 4898
rect 31388 4844 31444 4846
rect 33740 4844 33796 4900
rect 33292 4732 33348 4788
rect 32284 4396 32340 4452
rect 30044 4114 30100 4116
rect 30044 4062 30046 4114
rect 30046 4062 30098 4114
rect 30098 4062 30100 4114
rect 30044 4060 30100 4062
rect 31164 3836 31220 3892
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
rect 29148 3500 29204 3556
rect 30044 3388 30100 3444
rect 31276 3554 31332 3556
rect 31276 3502 31278 3554
rect 31278 3502 31330 3554
rect 31330 3502 31332 3554
rect 31276 3500 31332 3502
rect 33404 4060 33460 4116
rect 34860 4450 34916 4452
rect 34860 4398 34862 4450
rect 34862 4398 34914 4450
rect 34914 4398 34916 4450
rect 34860 4396 34916 4398
rect 35308 4114 35364 4116
rect 35308 4062 35310 4114
rect 35310 4062 35362 4114
rect 35362 4062 35364 4114
rect 35308 4060 35364 4062
rect 34412 3836 34468 3892
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34524 3612 34580 3668
rect 33740 3442 33796 3444
rect 33740 3390 33742 3442
rect 33742 3390 33794 3442
rect 33794 3390 33796 3442
rect 33740 3388 33796 3390
rect 37212 7980 37268 8036
rect 37548 8092 37604 8148
rect 37212 7756 37268 7812
rect 36652 7698 36708 7700
rect 36652 7646 36654 7698
rect 36654 7646 36706 7698
rect 36706 7646 36708 7698
rect 36652 7644 36708 7646
rect 37548 6690 37604 6692
rect 37548 6638 37550 6690
rect 37550 6638 37602 6690
rect 37602 6638 37604 6690
rect 37548 6636 37604 6638
rect 37884 8034 37940 8036
rect 37884 7982 37886 8034
rect 37886 7982 37938 8034
rect 37938 7982 37940 8034
rect 37884 7980 37940 7982
rect 37884 7644 37940 7700
rect 39788 10610 39844 10612
rect 39788 10558 39790 10610
rect 39790 10558 39842 10610
rect 39842 10558 39844 10610
rect 39788 10556 39844 10558
rect 41468 15596 41524 15652
rect 41692 16210 41748 16212
rect 41692 16158 41694 16210
rect 41694 16158 41746 16210
rect 41746 16158 41748 16210
rect 41692 16156 41748 16158
rect 41132 12684 41188 12740
rect 41020 11340 41076 11396
rect 41132 10780 41188 10836
rect 40796 10444 40852 10500
rect 39676 9436 39732 9492
rect 40796 9660 40852 9716
rect 39452 9266 39508 9268
rect 39452 9214 39454 9266
rect 39454 9214 39506 9266
rect 39506 9214 39508 9266
rect 39452 9212 39508 9214
rect 38780 8930 38836 8932
rect 38780 8878 38782 8930
rect 38782 8878 38834 8930
rect 38834 8878 38836 8930
rect 38780 8876 38836 8878
rect 41244 9212 41300 9268
rect 40796 8876 40852 8932
rect 42476 20300 42532 20356
rect 42364 19740 42420 19796
rect 42588 20188 42644 20244
rect 42364 17276 42420 17332
rect 41692 13916 41748 13972
rect 41916 11394 41972 11396
rect 41916 11342 41918 11394
rect 41918 11342 41970 11394
rect 41970 11342 41972 11394
rect 41916 11340 41972 11342
rect 42924 19180 42980 19236
rect 43820 26908 43876 26964
rect 44156 27132 44212 27188
rect 44716 27858 44772 27860
rect 44716 27806 44718 27858
rect 44718 27806 44770 27858
rect 44770 27806 44772 27858
rect 44716 27804 44772 27806
rect 44268 26236 44324 26292
rect 43596 23436 43652 23492
rect 43260 22482 43316 22484
rect 43260 22430 43262 22482
rect 43262 22430 43314 22482
rect 43314 22430 43316 22482
rect 43260 22428 43316 22430
rect 43484 21532 43540 21588
rect 43148 20860 43204 20916
rect 43596 20860 43652 20916
rect 43484 20188 43540 20244
rect 43148 19964 43204 20020
rect 43036 18620 43092 18676
rect 43596 19180 43652 19236
rect 44044 22258 44100 22260
rect 44044 22206 44046 22258
rect 44046 22206 44098 22258
rect 44098 22206 44100 22258
rect 44044 22204 44100 22206
rect 44268 22092 44324 22148
rect 44492 22428 44548 22484
rect 44044 20914 44100 20916
rect 44044 20862 44046 20914
rect 44046 20862 44098 20914
rect 44098 20862 44100 20914
rect 44044 20860 44100 20862
rect 42812 18060 42868 18116
rect 43820 17724 43876 17780
rect 43148 16658 43204 16660
rect 43148 16606 43150 16658
rect 43150 16606 43202 16658
rect 43202 16606 43204 16658
rect 43148 16604 43204 16606
rect 43596 16882 43652 16884
rect 43596 16830 43598 16882
rect 43598 16830 43650 16882
rect 43650 16830 43652 16882
rect 43596 16828 43652 16830
rect 42700 15932 42756 15988
rect 43820 15986 43876 15988
rect 43820 15934 43822 15986
rect 43822 15934 43874 15986
rect 43874 15934 43876 15986
rect 43820 15932 43876 15934
rect 44044 19068 44100 19124
rect 44156 18284 44212 18340
rect 44044 17836 44100 17892
rect 44716 23266 44772 23268
rect 44716 23214 44718 23266
rect 44718 23214 44770 23266
rect 44770 23214 44772 23266
rect 44716 23212 44772 23214
rect 44716 17836 44772 17892
rect 44268 17778 44324 17780
rect 44268 17726 44270 17778
rect 44270 17726 44322 17778
rect 44322 17726 44324 17778
rect 44268 17724 44324 17726
rect 42588 12348 42644 12404
rect 45276 33516 45332 33572
rect 46172 34242 46228 34244
rect 46172 34190 46174 34242
rect 46174 34190 46226 34242
rect 46226 34190 46228 34242
rect 46172 34188 46228 34190
rect 46956 34188 47012 34244
rect 46956 32396 47012 32452
rect 44940 29932 44996 29988
rect 47516 32396 47572 32452
rect 48300 32396 48356 32452
rect 47516 31388 47572 31444
rect 48300 31388 48356 31444
rect 45612 29986 45668 29988
rect 45612 29934 45614 29986
rect 45614 29934 45666 29986
rect 45666 29934 45668 29986
rect 45612 29932 45668 29934
rect 47180 30156 47236 30212
rect 46732 29986 46788 29988
rect 46732 29934 46734 29986
rect 46734 29934 46786 29986
rect 46786 29934 46788 29986
rect 46732 29932 46788 29934
rect 45500 28642 45556 28644
rect 45500 28590 45502 28642
rect 45502 28590 45554 28642
rect 45554 28590 45556 28642
rect 45500 28588 45556 28590
rect 46284 28642 46340 28644
rect 46284 28590 46286 28642
rect 46286 28590 46338 28642
rect 46338 28590 46340 28642
rect 46284 28588 46340 28590
rect 46732 28588 46788 28644
rect 46844 29372 46900 29428
rect 46956 28588 47012 28644
rect 46396 28140 46452 28196
rect 45500 28082 45556 28084
rect 45500 28030 45502 28082
rect 45502 28030 45554 28082
rect 45554 28030 45556 28082
rect 45500 28028 45556 28030
rect 46060 27970 46116 27972
rect 46060 27918 46062 27970
rect 46062 27918 46114 27970
rect 46114 27918 46116 27970
rect 46060 27916 46116 27918
rect 45836 27244 45892 27300
rect 45276 26908 45332 26964
rect 44940 25228 44996 25284
rect 45388 27132 45444 27188
rect 45612 27020 45668 27076
rect 45388 25618 45444 25620
rect 45388 25566 45390 25618
rect 45390 25566 45442 25618
rect 45442 25566 45444 25618
rect 45388 25564 45444 25566
rect 44940 22482 44996 22484
rect 44940 22430 44942 22482
rect 44942 22430 44994 22482
rect 44994 22430 44996 22482
rect 44940 22428 44996 22430
rect 45164 22204 45220 22260
rect 45500 22092 45556 22148
rect 46508 25564 46564 25620
rect 46172 23884 46228 23940
rect 45948 21644 46004 21700
rect 45052 19292 45108 19348
rect 44940 18396 44996 18452
rect 45052 17778 45108 17780
rect 45052 17726 45054 17778
rect 45054 17726 45106 17778
rect 45106 17726 45108 17778
rect 45052 17724 45108 17726
rect 44716 16770 44772 16772
rect 44716 16718 44718 16770
rect 44718 16718 44770 16770
rect 44770 16718 44772 16770
rect 44716 16716 44772 16718
rect 44604 16604 44660 16660
rect 44604 15820 44660 15876
rect 44828 15932 44884 15988
rect 44268 15036 44324 15092
rect 45052 15874 45108 15876
rect 45052 15822 45054 15874
rect 45054 15822 45106 15874
rect 45106 15822 45108 15874
rect 45052 15820 45108 15822
rect 45500 15932 45556 15988
rect 45164 13970 45220 13972
rect 45164 13918 45166 13970
rect 45166 13918 45218 13970
rect 45218 13918 45220 13970
rect 45164 13916 45220 13918
rect 44940 12738 44996 12740
rect 44940 12686 44942 12738
rect 44942 12686 44994 12738
rect 44994 12686 44996 12738
rect 44940 12684 44996 12686
rect 44828 12348 44884 12404
rect 43596 12066 43652 12068
rect 43596 12014 43598 12066
rect 43598 12014 43650 12066
rect 43650 12014 43652 12066
rect 43596 12012 43652 12014
rect 44380 11788 44436 11844
rect 42140 10444 42196 10500
rect 41916 9660 41972 9716
rect 40572 8146 40628 8148
rect 40572 8094 40574 8146
rect 40574 8094 40626 8146
rect 40626 8094 40628 8146
rect 40572 8092 40628 8094
rect 38780 7532 38836 7588
rect 37100 6524 37156 6580
rect 36988 6076 37044 6132
rect 37100 5292 37156 5348
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 36428 3554 36484 3556
rect 36428 3502 36430 3554
rect 36430 3502 36482 3554
rect 36482 3502 36484 3554
rect 36428 3500 36484 3502
rect 38668 6412 38724 6468
rect 39004 6188 39060 6244
rect 38556 5964 38612 6020
rect 37996 5346 38052 5348
rect 37996 5294 37998 5346
rect 37998 5294 38050 5346
rect 38050 5294 38052 5346
rect 37996 5292 38052 5294
rect 38444 5068 38500 5124
rect 37100 3500 37156 3556
rect 37884 3612 37940 3668
rect 36764 3276 36820 3332
rect 38780 5010 38836 5012
rect 38780 4958 38782 5010
rect 38782 4958 38834 5010
rect 38834 4958 38836 5010
rect 38780 4956 38836 4958
rect 40236 7196 40292 7252
rect 39788 6466 39844 6468
rect 39788 6414 39790 6466
rect 39790 6414 39842 6466
rect 39842 6414 39844 6466
rect 39788 6412 39844 6414
rect 39676 6018 39732 6020
rect 39676 5966 39678 6018
rect 39678 5966 39730 6018
rect 39730 5966 39732 6018
rect 39676 5964 39732 5966
rect 43484 10332 43540 10388
rect 41692 8204 41748 8260
rect 43820 8316 43876 8372
rect 42364 8092 42420 8148
rect 43148 8092 43204 8148
rect 39452 4956 39508 5012
rect 39116 4396 39172 4452
rect 39788 3554 39844 3556
rect 39788 3502 39790 3554
rect 39790 3502 39842 3554
rect 39842 3502 39844 3554
rect 39788 3500 39844 3502
rect 38892 3330 38948 3332
rect 38892 3278 38894 3330
rect 38894 3278 38946 3330
rect 38946 3278 38948 3330
rect 38892 3276 38948 3278
rect 38444 2940 38500 2996
rect 41580 7250 41636 7252
rect 41580 7198 41582 7250
rect 41582 7198 41634 7250
rect 41634 7198 41636 7250
rect 41580 7196 41636 7198
rect 40012 4450 40068 4452
rect 40012 4398 40014 4450
rect 40014 4398 40066 4450
rect 40066 4398 40068 4450
rect 40012 4396 40068 4398
rect 40348 4450 40404 4452
rect 40348 4398 40350 4450
rect 40350 4398 40402 4450
rect 40402 4398 40404 4450
rect 40348 4396 40404 4398
rect 41020 4284 41076 4340
rect 40796 3666 40852 3668
rect 40796 3614 40798 3666
rect 40798 3614 40850 3666
rect 40850 3614 40852 3666
rect 40796 3612 40852 3614
rect 40124 3276 40180 3332
rect 42476 7532 42532 7588
rect 44268 7586 44324 7588
rect 44268 7534 44270 7586
rect 44270 7534 44322 7586
rect 44322 7534 44324 7586
rect 44268 7532 44324 7534
rect 43148 7474 43204 7476
rect 43148 7422 43150 7474
rect 43150 7422 43202 7474
rect 43202 7422 43204 7474
rect 43148 7420 43204 7422
rect 43148 6748 43204 6804
rect 42364 6636 42420 6692
rect 42028 5964 42084 6020
rect 42924 5964 42980 6020
rect 43708 6690 43764 6692
rect 43708 6638 43710 6690
rect 43710 6638 43762 6690
rect 43762 6638 43764 6690
rect 43708 6636 43764 6638
rect 43260 6076 43316 6132
rect 46060 20018 46116 20020
rect 46060 19966 46062 20018
rect 46062 19966 46114 20018
rect 46114 19966 46116 20018
rect 46060 19964 46116 19966
rect 45836 19122 45892 19124
rect 45836 19070 45838 19122
rect 45838 19070 45890 19122
rect 45890 19070 45892 19122
rect 45836 19068 45892 19070
rect 46060 18620 46116 18676
rect 45836 18450 45892 18452
rect 45836 18398 45838 18450
rect 45838 18398 45890 18450
rect 45890 18398 45892 18450
rect 45836 18396 45892 18398
rect 45724 17890 45780 17892
rect 45724 17838 45726 17890
rect 45726 17838 45778 17890
rect 45778 17838 45780 17890
rect 45724 17836 45780 17838
rect 45724 16828 45780 16884
rect 46284 17724 46340 17780
rect 46060 16156 46116 16212
rect 46956 25394 47012 25396
rect 46956 25342 46958 25394
rect 46958 25342 47010 25394
rect 47010 25342 47012 25394
rect 46956 25340 47012 25342
rect 47180 23884 47236 23940
rect 47292 23660 47348 23716
rect 46620 18284 46676 18340
rect 46732 16882 46788 16884
rect 46732 16830 46734 16882
rect 46734 16830 46786 16882
rect 46786 16830 46788 16882
rect 46732 16828 46788 16830
rect 48300 29426 48356 29428
rect 48300 29374 48302 29426
rect 48302 29374 48354 29426
rect 48354 29374 48356 29426
rect 48300 29372 48356 29374
rect 47964 28642 48020 28644
rect 47964 28590 47966 28642
rect 47966 28590 48018 28642
rect 48018 28590 48020 28642
rect 47964 28588 48020 28590
rect 47292 16716 47348 16772
rect 46620 15538 46676 15540
rect 46620 15486 46622 15538
rect 46622 15486 46674 15538
rect 46674 15486 46676 15538
rect 46620 15484 46676 15486
rect 47292 15484 47348 15540
rect 47740 26012 47796 26068
rect 48300 25340 48356 25396
rect 47628 23212 47684 23268
rect 48412 23884 48468 23940
rect 47964 21698 48020 21700
rect 47964 21646 47966 21698
rect 47966 21646 48018 21698
rect 48018 21646 48020 21698
rect 47964 21644 48020 21646
rect 47740 18284 47796 18340
rect 48300 18338 48356 18340
rect 48300 18286 48302 18338
rect 48302 18286 48354 18338
rect 48354 18286 48356 18338
rect 48300 18284 48356 18286
rect 47740 16770 47796 16772
rect 47740 16718 47742 16770
rect 47742 16718 47794 16770
rect 47794 16718 47796 16770
rect 47740 16716 47796 16718
rect 48300 16210 48356 16212
rect 48300 16158 48302 16210
rect 48302 16158 48354 16210
rect 48354 16158 48356 16210
rect 48300 16156 48356 16158
rect 46508 13916 46564 13972
rect 45836 13746 45892 13748
rect 45836 13694 45838 13746
rect 45838 13694 45890 13746
rect 45890 13694 45892 13746
rect 45836 13692 45892 13694
rect 45276 12012 45332 12068
rect 46284 11788 46340 11844
rect 45276 10834 45332 10836
rect 45276 10782 45278 10834
rect 45278 10782 45330 10834
rect 45330 10782 45332 10834
rect 45276 10780 45332 10782
rect 44828 6636 44884 6692
rect 44940 10444 44996 10500
rect 45724 10780 45780 10836
rect 45948 10668 46004 10724
rect 45500 10444 45556 10500
rect 46956 11788 47012 11844
rect 47404 13692 47460 13748
rect 47740 13692 47796 13748
rect 48300 13692 48356 13748
rect 47292 10722 47348 10724
rect 47292 10670 47294 10722
rect 47294 10670 47346 10722
rect 47346 10670 47348 10722
rect 47292 10668 47348 10670
rect 46844 10386 46900 10388
rect 46844 10334 46846 10386
rect 46846 10334 46898 10386
rect 46898 10334 46900 10386
rect 46844 10332 46900 10334
rect 46508 9884 46564 9940
rect 48300 9938 48356 9940
rect 48300 9886 48302 9938
rect 48302 9886 48354 9938
rect 48354 9886 48356 9938
rect 48300 9884 48356 9886
rect 44156 6076 44212 6132
rect 42140 5122 42196 5124
rect 42140 5070 42142 5122
rect 42142 5070 42194 5122
rect 42194 5070 42196 5122
rect 42140 5068 42196 5070
rect 42364 3612 42420 3668
rect 43260 4396 43316 4452
rect 43820 4338 43876 4340
rect 43820 4286 43822 4338
rect 43822 4286 43874 4338
rect 43874 4286 43876 4338
rect 43820 4284 43876 4286
rect 45388 8204 45444 8260
rect 45052 7532 45108 7588
rect 45052 6690 45108 6692
rect 45052 6638 45054 6690
rect 45054 6638 45106 6690
rect 45106 6638 45108 6690
rect 45052 6636 45108 6638
rect 46956 7532 47012 7588
rect 45500 7420 45556 7476
rect 46844 6748 46900 6804
rect 47628 7586 47684 7588
rect 47628 7534 47630 7586
rect 47630 7534 47682 7586
rect 47682 7534 47684 7586
rect 47628 7532 47684 7534
rect 48300 7532 48356 7588
rect 45948 6524 46004 6580
rect 44940 6130 44996 6132
rect 44940 6078 44942 6130
rect 44942 6078 44994 6130
rect 44994 6078 44996 6130
rect 44940 6076 44996 6078
rect 44604 3666 44660 3668
rect 44604 3614 44606 3666
rect 44606 3614 44658 3666
rect 44658 3614 44660 3666
rect 44604 3612 44660 3614
rect 42476 3500 42532 3556
rect 43596 3554 43652 3556
rect 43596 3502 43598 3554
rect 43598 3502 43650 3554
rect 43650 3502 43652 3554
rect 43596 3500 43652 3502
rect 43484 3388 43540 3444
rect 42700 3330 42756 3332
rect 42700 3278 42702 3330
rect 42702 3278 42754 3330
rect 42754 3278 42756 3330
rect 42700 3276 42756 3278
rect 46508 3388 46564 3444
rect 45724 3276 45780 3332
rect 47180 6636 47236 6692
rect 48188 6636 48244 6692
rect 47516 6578 47572 6580
rect 47516 6526 47518 6578
rect 47518 6526 47570 6578
rect 47570 6526 47572 6578
rect 47516 6524 47572 6526
rect 48300 6524 48356 6580
rect 47404 3330 47460 3332
rect 47404 3278 47406 3330
rect 47406 3278 47458 3330
rect 47458 3278 47460 3330
rect 47404 3276 47460 3278
<< metal3 >>
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 14466 48972 14476 49028
rect 14532 48972 16828 49028
rect 16884 48972 17612 49028
rect 17668 48972 17678 49028
rect 29250 48972 29260 49028
rect 29316 48972 32396 49028
rect 32452 48972 32462 49028
rect 15026 48748 15036 48804
rect 15092 48748 16268 48804
rect 16324 48748 16334 48804
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 18386 48300 18396 48356
rect 18452 48300 20076 48356
rect 20132 48300 21532 48356
rect 21588 48300 21598 48356
rect 21970 48300 21980 48356
rect 22036 48300 22652 48356
rect 22708 48300 24332 48356
rect 24388 48300 24398 48356
rect 25666 48300 25676 48356
rect 25732 48300 28252 48356
rect 28308 48300 28318 48356
rect 30818 48300 30828 48356
rect 30884 48300 32172 48356
rect 32228 48300 32238 48356
rect 38882 48300 38892 48356
rect 38948 48300 40012 48356
rect 40068 48300 40078 48356
rect 16594 48188 16604 48244
rect 16660 48188 17276 48244
rect 17332 48188 17342 48244
rect 24332 48132 24388 48300
rect 30258 48188 30268 48244
rect 30324 48188 34076 48244
rect 34132 48188 35756 48244
rect 35812 48188 35822 48244
rect 24332 48076 26908 48132
rect 26964 48076 26974 48132
rect 30706 48076 30716 48132
rect 30772 48076 33740 48132
rect 33796 48076 33806 48132
rect 19842 47964 19852 48020
rect 19908 47964 20748 48020
rect 20804 47964 21308 48020
rect 21364 47964 21980 48020
rect 22036 47964 22046 48020
rect 27682 47964 27692 48020
rect 27748 47964 30828 48020
rect 30884 47964 30894 48020
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 32274 47404 32284 47460
rect 32340 47404 33068 47460
rect 33124 47404 33134 47460
rect 17378 47292 17388 47348
rect 17444 47292 18172 47348
rect 18228 47292 18620 47348
rect 18676 47292 19292 47348
rect 19348 47292 19358 47348
rect 38210 47292 38220 47348
rect 38276 47292 38892 47348
rect 38948 47292 38958 47348
rect 21410 47180 21420 47236
rect 21476 47180 22988 47236
rect 23044 47180 23054 47236
rect 32610 47180 32620 47236
rect 32676 47180 33516 47236
rect 33572 47180 35980 47236
rect 36036 47180 36046 47236
rect 37986 47180 37996 47236
rect 38052 47180 38332 47236
rect 38388 47180 41692 47236
rect 41748 47180 42364 47236
rect 42420 47180 42430 47236
rect 34972 47068 35532 47124
rect 35588 47068 35598 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 28466 46956 28476 47012
rect 28532 46956 30716 47012
rect 30772 46956 30782 47012
rect 31892 46956 33740 47012
rect 33796 46956 33806 47012
rect 9986 46844 9996 46900
rect 10052 46844 11004 46900
rect 11060 46844 11676 46900
rect 11732 46844 12908 46900
rect 12964 46844 12974 46900
rect 24434 46844 24444 46900
rect 24500 46844 25340 46900
rect 25396 46844 25406 46900
rect 31892 46788 31948 46956
rect 30146 46732 30156 46788
rect 30212 46732 31948 46788
rect 32004 46732 32014 46788
rect 32386 46732 32396 46788
rect 32452 46732 33404 46788
rect 33460 46732 33470 46788
rect 33404 46676 33460 46732
rect 34972 46676 35028 47068
rect 37090 46956 37100 47012
rect 37156 46956 39228 47012
rect 39284 46956 40236 47012
rect 40292 46956 41804 47012
rect 41860 46956 41870 47012
rect 38658 46732 38668 46788
rect 38724 46732 40012 46788
rect 40068 46732 40078 46788
rect 33404 46620 35028 46676
rect 34972 46564 35028 46620
rect 34962 46508 34972 46564
rect 35028 46508 35038 46564
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 16818 46060 16828 46116
rect 16884 46060 18732 46116
rect 18788 46060 19628 46116
rect 19684 46060 21196 46116
rect 21252 46060 21262 46116
rect 26898 46060 26908 46116
rect 26964 46060 27692 46116
rect 27748 46060 27758 46116
rect 40002 46060 40012 46116
rect 40068 46060 41132 46116
rect 41188 46060 41198 46116
rect 20738 45836 20748 45892
rect 20804 45836 21868 45892
rect 21924 45836 21934 45892
rect 11106 45724 11116 45780
rect 11172 45724 11676 45780
rect 11732 45724 12684 45780
rect 12740 45724 14364 45780
rect 14420 45724 14430 45780
rect 14802 45724 14812 45780
rect 14868 45724 15708 45780
rect 15764 45724 16156 45780
rect 16212 45724 16222 45780
rect 11218 45612 11228 45668
rect 11284 45612 12012 45668
rect 12068 45612 12078 45668
rect 22754 45612 22764 45668
rect 22820 45612 24332 45668
rect 24388 45612 24398 45668
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 17714 45388 17724 45444
rect 17780 45388 18508 45444
rect 18564 45388 19292 45444
rect 19348 45388 19358 45444
rect 28466 45276 28476 45332
rect 28532 45276 29036 45332
rect 29092 45276 29932 45332
rect 29988 45276 29998 45332
rect 34962 45276 34972 45332
rect 35028 45276 37436 45332
rect 37492 45276 38108 45332
rect 38164 45276 38174 45332
rect 30258 45164 30268 45220
rect 30324 45164 30604 45220
rect 30660 45164 39788 45220
rect 39844 45164 40908 45220
rect 40964 45164 40974 45220
rect 27010 45052 27020 45108
rect 27076 45052 30156 45108
rect 30212 45052 33404 45108
rect 33460 45052 33470 45108
rect 27906 44940 27916 44996
rect 27972 44940 30268 44996
rect 30324 44940 30334 44996
rect 41458 44940 41468 44996
rect 41524 44940 43036 44996
rect 43092 44940 43102 44996
rect 17826 44828 17836 44884
rect 17892 44828 19180 44884
rect 19236 44828 19246 44884
rect 25778 44828 25788 44884
rect 25844 44828 26348 44884
rect 26404 44828 26414 44884
rect 28354 44828 28364 44884
rect 28420 44828 29260 44884
rect 29316 44828 30716 44884
rect 30772 44828 30782 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 31602 44492 31612 44548
rect 31668 44492 41524 44548
rect 20962 44268 20972 44324
rect 21028 44268 23324 44324
rect 23380 44268 23390 44324
rect 30706 44268 30716 44324
rect 30772 44268 31948 44324
rect 32004 44268 32014 44324
rect 41468 44212 41524 44492
rect 34290 44156 34300 44212
rect 34356 44156 34972 44212
rect 35028 44156 35038 44212
rect 41458 44156 41468 44212
rect 41524 44156 43372 44212
rect 43428 44156 45164 44212
rect 45220 44156 45230 44212
rect 25666 44044 25676 44100
rect 25732 44044 26236 44100
rect 26292 44044 26302 44100
rect 35074 44044 35084 44100
rect 35140 44044 35644 44100
rect 35700 44044 35710 44100
rect 41122 44044 41132 44100
rect 41188 44044 41804 44100
rect 41860 44044 41870 44100
rect 31892 43932 34636 43988
rect 34692 43932 34702 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 31892 43764 31948 43932
rect 10882 43708 10892 43764
rect 10948 43708 12348 43764
rect 12404 43708 12414 43764
rect 30594 43708 30604 43764
rect 30660 43708 31948 43764
rect 32946 43708 32956 43764
rect 33012 43708 33404 43764
rect 33460 43708 36316 43764
rect 36372 43708 36382 43764
rect 12226 43596 12236 43652
rect 12292 43596 13132 43652
rect 13188 43596 13198 43652
rect 19394 43596 19404 43652
rect 19460 43596 20412 43652
rect 20468 43596 20478 43652
rect 32498 43596 32508 43652
rect 32564 43596 33628 43652
rect 33684 43596 34412 43652
rect 34468 43596 34860 43652
rect 34916 43596 34926 43652
rect 12002 43484 12012 43540
rect 12068 43484 13580 43540
rect 13636 43484 13646 43540
rect 28018 43484 28028 43540
rect 28084 43484 28700 43540
rect 28756 43484 28766 43540
rect 32050 43484 32060 43540
rect 32116 43484 34076 43540
rect 34132 43484 34142 43540
rect 7522 43372 7532 43428
rect 7588 43372 8316 43428
rect 8372 43372 8876 43428
rect 8932 43372 10892 43428
rect 10948 43372 11564 43428
rect 11620 43372 11630 43428
rect 12114 43372 12124 43428
rect 12180 43372 17948 43428
rect 18004 43372 18014 43428
rect 22082 43372 22092 43428
rect 22148 43372 22540 43428
rect 22596 43372 22606 43428
rect 29810 43260 29820 43316
rect 29876 43260 31500 43316
rect 31556 43260 31566 43316
rect 42018 43260 42028 43316
rect 42084 43260 42924 43316
rect 42980 43260 42990 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 20178 42924 20188 42980
rect 20244 42924 21420 42980
rect 21476 42924 21486 42980
rect 7634 42700 7644 42756
rect 7700 42700 8988 42756
rect 9044 42700 10220 42756
rect 10276 42700 10286 42756
rect 11106 42700 11116 42756
rect 11172 42700 12012 42756
rect 12068 42700 12078 42756
rect 13906 42700 13916 42756
rect 13972 42700 18396 42756
rect 18452 42700 18462 42756
rect 24546 42700 24556 42756
rect 24612 42700 25228 42756
rect 25284 42700 25294 42756
rect 9762 42588 9772 42644
rect 9828 42588 10668 42644
rect 10724 42588 10734 42644
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 9874 42252 9884 42308
rect 9940 42252 11452 42308
rect 11508 42252 11518 42308
rect 14018 42252 14028 42308
rect 14084 42252 14700 42308
rect 14756 42252 15148 42308
rect 9650 42140 9660 42196
rect 9716 42140 10444 42196
rect 10500 42140 10510 42196
rect 15092 42084 15148 42252
rect 42914 42140 42924 42196
rect 42980 42140 43820 42196
rect 43876 42140 45724 42196
rect 45780 42140 45790 42196
rect 8372 42028 9772 42084
rect 9828 42028 9838 42084
rect 15092 42028 15596 42084
rect 15652 42028 18284 42084
rect 18340 42028 18350 42084
rect 25554 42028 25564 42084
rect 25620 42028 26236 42084
rect 26292 42028 26908 42084
rect 26964 42028 26974 42084
rect 8372 41972 8428 42028
rect 7522 41916 7532 41972
rect 7588 41916 8428 41972
rect 15474 41916 15484 41972
rect 15540 41916 16268 41972
rect 16324 41916 18396 41972
rect 18452 41916 19180 41972
rect 19236 41916 19628 41972
rect 19684 41916 19694 41972
rect 37762 41916 37772 41972
rect 37828 41916 39340 41972
rect 39396 41916 41020 41972
rect 41076 41916 41692 41972
rect 41748 41916 42364 41972
rect 42420 41916 42430 41972
rect 21746 41804 21756 41860
rect 21812 41804 22316 41860
rect 22372 41804 22382 41860
rect 30034 41804 30044 41860
rect 30100 41804 30716 41860
rect 30772 41804 30782 41860
rect 35634 41804 35644 41860
rect 35700 41804 38780 41860
rect 38836 41804 38846 41860
rect 6850 41692 6860 41748
rect 6916 41692 7644 41748
rect 7700 41692 7710 41748
rect 30146 41580 30156 41636
rect 30212 41580 31052 41636
rect 31108 41580 31118 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 34178 41356 34188 41412
rect 34244 41356 35308 41412
rect 35364 41356 36092 41412
rect 36148 41356 36158 41412
rect 17826 41244 17836 41300
rect 17892 41244 19180 41300
rect 19236 41244 19246 41300
rect 27346 41132 27356 41188
rect 27412 41132 27804 41188
rect 27860 41132 29596 41188
rect 29652 41132 29662 41188
rect 24434 41020 24444 41076
rect 24500 41020 25340 41076
rect 25396 41020 25406 41076
rect 34066 41020 34076 41076
rect 34132 41020 34972 41076
rect 35028 41020 35532 41076
rect 35588 41020 35598 41076
rect 40114 41020 40124 41076
rect 40180 41020 42812 41076
rect 42868 41020 43484 41076
rect 43540 41020 43550 41076
rect 11554 40908 11564 40964
rect 11620 40908 12460 40964
rect 12516 40908 12526 40964
rect 15092 40908 15372 40964
rect 15428 40908 17052 40964
rect 17108 40908 17118 40964
rect 21746 40908 21756 40964
rect 21812 40908 23100 40964
rect 23156 40908 23166 40964
rect 31714 40908 31724 40964
rect 31780 40908 32508 40964
rect 32564 40908 32574 40964
rect 39218 40908 39228 40964
rect 39284 40908 40012 40964
rect 40068 40908 40078 40964
rect 40674 40908 40684 40964
rect 40740 40908 41804 40964
rect 41860 40908 42588 40964
rect 42644 40908 42654 40964
rect 15092 40740 15148 40908
rect 22418 40796 22428 40852
rect 22484 40796 24556 40852
rect 24612 40796 24622 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 14578 40684 14588 40740
rect 14644 40684 15148 40740
rect 12786 40572 12796 40628
rect 12852 40572 14476 40628
rect 14532 40572 14542 40628
rect 15026 40572 15036 40628
rect 15092 40572 15484 40628
rect 15540 40572 15550 40628
rect 8372 40460 8988 40516
rect 9044 40460 12236 40516
rect 12292 40460 12302 40516
rect 15698 40460 15708 40516
rect 15764 40460 17612 40516
rect 17668 40460 17678 40516
rect 40002 40460 40012 40516
rect 40068 40460 40684 40516
rect 40740 40460 40750 40516
rect 8372 40404 8428 40460
rect 4834 40348 4844 40404
rect 4900 40348 5740 40404
rect 5796 40348 5806 40404
rect 7634 40348 7644 40404
rect 7700 40348 8428 40404
rect 12114 40348 12124 40404
rect 12180 40348 12908 40404
rect 12964 40348 16268 40404
rect 16324 40348 16334 40404
rect 17490 40348 17500 40404
rect 17556 40348 19180 40404
rect 19236 40348 19246 40404
rect 20178 40348 20188 40404
rect 20244 40348 23548 40404
rect 23604 40348 23614 40404
rect 25666 40348 25676 40404
rect 25732 40348 25742 40404
rect 29586 40348 29596 40404
rect 29652 40348 30492 40404
rect 30548 40348 31836 40404
rect 31892 40348 32508 40404
rect 32564 40348 32574 40404
rect 41346 40348 41356 40404
rect 41412 40348 42364 40404
rect 42420 40348 42430 40404
rect 42802 40348 42812 40404
rect 42868 40348 43148 40404
rect 43204 40348 45052 40404
rect 45108 40348 45118 40404
rect 25676 40292 25732 40348
rect 25106 40236 25116 40292
rect 25172 40236 25732 40292
rect 31714 40236 31724 40292
rect 31780 40236 31948 40292
rect 32004 40236 34076 40292
rect 34132 40236 34142 40292
rect 9202 40124 9212 40180
rect 9268 40124 9996 40180
rect 10052 40124 10062 40180
rect 30258 40124 30268 40180
rect 30324 40124 31052 40180
rect 31108 40124 31118 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 7074 39788 7084 39844
rect 7140 39788 10556 39844
rect 10612 39788 11564 39844
rect 11620 39788 11630 39844
rect 5730 39676 5740 39732
rect 5796 39676 9324 39732
rect 9380 39676 9390 39732
rect 16930 39564 16940 39620
rect 16996 39564 20188 39620
rect 20244 39564 20254 39620
rect 22082 39564 22092 39620
rect 22148 39564 22764 39620
rect 22820 39564 24780 39620
rect 24836 39564 24846 39620
rect 12450 39452 12460 39508
rect 12516 39452 13244 39508
rect 13300 39452 14028 39508
rect 14084 39452 15148 39508
rect 20626 39452 20636 39508
rect 20692 39452 21756 39508
rect 21812 39452 21822 39508
rect 15092 39396 15148 39452
rect 10546 39340 10556 39396
rect 10612 39340 13132 39396
rect 13188 39340 14588 39396
rect 14644 39340 14654 39396
rect 15092 39340 21700 39396
rect 24322 39340 24332 39396
rect 24388 39340 26460 39396
rect 26516 39340 26526 39396
rect 27458 39340 27468 39396
rect 27524 39340 34524 39396
rect 34580 39340 35532 39396
rect 35588 39340 35598 39396
rect 21644 39284 21700 39340
rect 11778 39228 11788 39284
rect 11844 39228 12908 39284
rect 12964 39228 13692 39284
rect 13748 39228 13758 39284
rect 21634 39228 21644 39284
rect 21700 39228 21710 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 14690 39004 14700 39060
rect 14756 39004 15820 39060
rect 15876 39004 17948 39060
rect 18004 39004 18508 39060
rect 18564 39004 18574 39060
rect 21858 39004 21868 39060
rect 21924 39004 22652 39060
rect 22708 39004 22718 39060
rect 17602 38892 17612 38948
rect 17668 38892 19124 38948
rect 29026 38892 29036 38948
rect 29092 38892 30268 38948
rect 30324 38892 30334 38948
rect 35074 38892 35084 38948
rect 35140 38892 36092 38948
rect 36148 38892 37212 38948
rect 37268 38892 37278 38948
rect 19068 38836 19124 38892
rect 2146 38780 2156 38836
rect 2212 38780 5180 38836
rect 5236 38780 5740 38836
rect 5796 38780 5806 38836
rect 9650 38780 9660 38836
rect 9716 38780 10780 38836
rect 10836 38780 12124 38836
rect 12180 38780 12684 38836
rect 12740 38780 12750 38836
rect 14914 38780 14924 38836
rect 14980 38780 17388 38836
rect 17444 38780 17454 38836
rect 18050 38780 18060 38836
rect 18116 38780 18844 38836
rect 18900 38780 18910 38836
rect 19058 38780 19068 38836
rect 19124 38780 19516 38836
rect 19572 38780 19582 38836
rect 23100 38780 24332 38836
rect 24388 38780 24398 38836
rect 24658 38780 24668 38836
rect 24724 38780 24734 38836
rect 31602 38780 31612 38836
rect 31668 38780 31678 38836
rect 38994 38780 39004 38836
rect 39060 38780 40012 38836
rect 40068 38780 40078 38836
rect 23100 38724 23156 38780
rect 24668 38724 24724 38780
rect 31612 38724 31668 38780
rect 11666 38668 11676 38724
rect 11732 38668 12236 38724
rect 12292 38668 13580 38724
rect 13636 38668 13646 38724
rect 18610 38668 18620 38724
rect 18676 38668 23156 38724
rect 23314 38668 23324 38724
rect 23380 38668 24108 38724
rect 24164 38668 25452 38724
rect 25508 38668 25788 38724
rect 25844 38668 25854 38724
rect 27794 38668 27804 38724
rect 27860 38668 28700 38724
rect 28756 38668 28766 38724
rect 31612 38668 33068 38724
rect 33124 38668 33134 38724
rect 10098 38556 10108 38612
rect 10164 38556 19068 38612
rect 19124 38556 19134 38612
rect 19282 38556 19292 38612
rect 19348 38556 20076 38612
rect 20132 38556 20142 38612
rect 20962 38556 20972 38612
rect 21028 38556 24220 38612
rect 24276 38556 24286 38612
rect 32386 38556 32396 38612
rect 32452 38556 34188 38612
rect 34244 38556 34254 38612
rect 13234 38444 13244 38500
rect 13300 38444 14140 38500
rect 14196 38444 25228 38500
rect 25284 38444 25294 38500
rect 32274 38444 32284 38500
rect 32340 38444 33292 38500
rect 33348 38444 33852 38500
rect 33908 38444 33918 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 13570 38332 13580 38388
rect 13636 38332 24108 38388
rect 24164 38332 25340 38388
rect 25396 38332 27468 38388
rect 27524 38332 27534 38388
rect 29474 38332 29484 38388
rect 29540 38332 33964 38388
rect 34020 38332 34030 38388
rect 6626 38220 6636 38276
rect 6692 38220 7420 38276
rect 7476 38220 7486 38276
rect 17714 38220 17724 38276
rect 17780 38220 17836 38276
rect 17892 38220 17902 38276
rect 19058 38220 19068 38276
rect 19124 38220 26684 38276
rect 26740 38220 26750 38276
rect 4946 38108 4956 38164
rect 5012 38108 5516 38164
rect 5572 38108 6076 38164
rect 6132 38108 9660 38164
rect 9716 38108 9726 38164
rect 13346 38108 13356 38164
rect 13412 38108 14812 38164
rect 14868 38108 14878 38164
rect 15092 38108 21252 38164
rect 21634 38108 21644 38164
rect 21700 38108 22988 38164
rect 23044 38108 23324 38164
rect 23380 38108 23390 38164
rect 23762 38108 23772 38164
rect 23828 38108 25004 38164
rect 25060 38108 25070 38164
rect 33954 38108 33964 38164
rect 34020 38108 35868 38164
rect 35924 38108 37996 38164
rect 38052 38108 38668 38164
rect 15092 38052 15148 38108
rect 4834 37996 4844 38052
rect 4900 37996 5292 38052
rect 5348 37996 6300 38052
rect 6356 37996 6366 38052
rect 13682 37996 13692 38052
rect 13748 37996 15148 38052
rect 16044 37996 19180 38052
rect 19236 37996 20188 38052
rect 20244 37996 20254 38052
rect 16044 37940 16100 37996
rect 2594 37884 2604 37940
rect 2660 37884 5740 37940
rect 5796 37884 5806 37940
rect 9426 37884 9436 37940
rect 9492 37884 10332 37940
rect 10388 37884 11564 37940
rect 11620 37884 11630 37940
rect 12114 37884 12124 37940
rect 12180 37884 16100 37940
rect 16258 37884 16268 37940
rect 16324 37884 17220 37940
rect 17714 37884 17724 37940
rect 17780 37884 19628 37940
rect 19684 37884 19694 37940
rect 20402 37884 20412 37940
rect 20468 37884 20972 37940
rect 21028 37884 21038 37940
rect 14690 37772 14700 37828
rect 14756 37772 16156 37828
rect 16212 37772 16222 37828
rect 16380 37604 16436 37884
rect 17164 37828 17220 37884
rect 17164 37772 17612 37828
rect 17668 37772 19404 37828
rect 19460 37772 19470 37828
rect 19628 37772 19852 37828
rect 19908 37772 19918 37828
rect 20066 37772 20076 37828
rect 20132 37772 20356 37828
rect 19628 37716 19684 37772
rect 20300 37716 20356 37772
rect 19618 37660 19628 37716
rect 19684 37660 19694 37716
rect 20290 37660 20300 37716
rect 20356 37660 20366 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 12338 37548 12348 37604
rect 12404 37548 13020 37604
rect 13076 37548 16436 37604
rect 21196 37492 21252 38108
rect 23772 38052 23828 38108
rect 38612 38052 38668 38108
rect 22194 37996 22204 38052
rect 22260 37996 23828 38052
rect 24210 37996 24220 38052
rect 24276 37996 24286 38052
rect 24770 37996 24780 38052
rect 24836 37996 25676 38052
rect 25732 37996 25742 38052
rect 26338 37996 26348 38052
rect 26404 37996 27692 38052
rect 27748 37996 27758 38052
rect 38612 37996 39116 38052
rect 39172 37996 39182 38052
rect 24220 37940 24276 37996
rect 24220 37884 24668 37940
rect 24724 37884 24734 37940
rect 35858 37884 35868 37940
rect 35924 37884 37660 37940
rect 37716 37884 38668 37940
rect 39890 37884 39900 37940
rect 39956 37884 41468 37940
rect 41524 37884 41534 37940
rect 38612 37828 38668 37884
rect 21746 37772 21756 37828
rect 21812 37772 21980 37828
rect 22036 37772 22046 37828
rect 24434 37772 24444 37828
rect 24500 37772 25900 37828
rect 25956 37772 27916 37828
rect 27972 37772 27982 37828
rect 30930 37772 30940 37828
rect 30996 37772 32956 37828
rect 33012 37772 34300 37828
rect 34356 37772 34366 37828
rect 38612 37772 39788 37828
rect 39844 37772 39854 37828
rect 25778 37660 25788 37716
rect 25844 37660 26348 37716
rect 26404 37660 26414 37716
rect 25218 37548 25228 37604
rect 25284 37548 26124 37604
rect 26180 37548 26460 37604
rect 26516 37548 36988 37604
rect 37044 37548 37054 37604
rect 4274 37436 4284 37492
rect 4340 37436 4732 37492
rect 4788 37436 6860 37492
rect 6916 37436 11676 37492
rect 11732 37436 11742 37492
rect 15474 37436 15484 37492
rect 15540 37436 18172 37492
rect 18228 37436 18238 37492
rect 21196 37436 27580 37492
rect 27636 37436 27646 37492
rect 42242 37436 42252 37492
rect 42308 37436 43484 37492
rect 43540 37436 43550 37492
rect 9986 37324 9996 37380
rect 10052 37324 11004 37380
rect 11060 37324 11070 37380
rect 11218 37324 11228 37380
rect 11284 37324 12012 37380
rect 12068 37324 12078 37380
rect 12338 37324 12348 37380
rect 12404 37324 13692 37380
rect 13748 37324 13758 37380
rect 13906 37324 13916 37380
rect 13972 37324 15036 37380
rect 15092 37324 15102 37380
rect 26852 37324 27692 37380
rect 27748 37324 27758 37380
rect 27906 37324 27916 37380
rect 27972 37324 29540 37380
rect 43138 37324 43148 37380
rect 43204 37324 44044 37380
rect 44100 37324 44110 37380
rect 26852 37268 26908 37324
rect 29484 37268 29540 37324
rect 9090 37212 9100 37268
rect 9156 37212 10108 37268
rect 10164 37212 10174 37268
rect 10434 37212 10444 37268
rect 10500 37212 11788 37268
rect 11844 37212 11854 37268
rect 14130 37212 14140 37268
rect 14196 37212 15372 37268
rect 15428 37212 26908 37268
rect 27010 37212 27020 37268
rect 27076 37212 27468 37268
rect 27524 37212 28700 37268
rect 28756 37212 28766 37268
rect 29474 37212 29484 37268
rect 29540 37212 29820 37268
rect 29876 37212 29886 37268
rect 39778 37212 39788 37268
rect 39844 37212 40180 37268
rect 40450 37212 40460 37268
rect 40516 37212 43372 37268
rect 43428 37212 44156 37268
rect 44212 37212 44222 37268
rect 40124 37156 40180 37212
rect 4162 37100 4172 37156
rect 4228 37100 4732 37156
rect 4788 37100 6860 37156
rect 6916 37100 10668 37156
rect 10724 37100 10734 37156
rect 12898 37100 12908 37156
rect 12964 37100 13692 37156
rect 13748 37100 13758 37156
rect 18722 37100 18732 37156
rect 18788 37100 20076 37156
rect 20132 37100 21308 37156
rect 21364 37100 31500 37156
rect 31556 37100 32508 37156
rect 32564 37100 33068 37156
rect 33124 37100 33134 37156
rect 33618 37100 33628 37156
rect 33684 37100 37324 37156
rect 37380 37100 39900 37156
rect 39956 37100 39966 37156
rect 40124 37100 41916 37156
rect 41972 37100 43708 37156
rect 43764 37100 43774 37156
rect 10770 36988 10780 37044
rect 10836 36988 13468 37044
rect 13524 36988 13534 37044
rect 15698 36988 15708 37044
rect 15764 36988 16492 37044
rect 16548 36988 17500 37044
rect 17556 36988 17566 37044
rect 17826 36988 17836 37044
rect 17892 36988 20244 37044
rect 20962 36988 20972 37044
rect 21028 36988 22204 37044
rect 22260 36988 22270 37044
rect 23090 36988 23100 37044
rect 23156 36988 23884 37044
rect 23940 36988 23950 37044
rect 24994 36988 25004 37044
rect 25060 36988 27356 37044
rect 27412 36988 27422 37044
rect 27570 36988 27580 37044
rect 27636 36988 28252 37044
rect 28308 36988 28318 37044
rect 29922 36988 29932 37044
rect 29988 36988 30828 37044
rect 30884 36988 30894 37044
rect 20188 36932 20244 36988
rect 16930 36876 16940 36932
rect 16996 36876 19404 36932
rect 19460 36876 19470 36932
rect 20188 36876 24780 36932
rect 24836 36876 24846 36932
rect 26002 36876 26012 36932
rect 26068 36876 27020 36932
rect 27076 36876 27086 36932
rect 28354 36876 28364 36932
rect 28420 36876 30492 36932
rect 30548 36876 30558 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 26012 36820 26068 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 18834 36764 18844 36820
rect 18900 36764 19292 36820
rect 19348 36764 19358 36820
rect 23492 36764 26068 36820
rect 29026 36764 29036 36820
rect 29092 36764 29708 36820
rect 29764 36764 29774 36820
rect 23492 36708 23548 36764
rect 19030 36652 19068 36708
rect 19124 36652 19134 36708
rect 19292 36652 23548 36708
rect 24882 36652 24892 36708
rect 24948 36652 25340 36708
rect 25396 36652 25406 36708
rect 33058 36652 33068 36708
rect 33124 36652 37436 36708
rect 37492 36652 39788 36708
rect 39844 36652 39854 36708
rect 19292 36596 19348 36652
rect 14354 36540 14364 36596
rect 14420 36540 15148 36596
rect 15204 36540 15372 36596
rect 15428 36540 19348 36596
rect 19618 36540 19628 36596
rect 19684 36540 20636 36596
rect 20692 36540 20702 36596
rect 24770 36540 24780 36596
rect 24836 36540 26908 36596
rect 26964 36540 26974 36596
rect 12786 36428 12796 36484
rect 12852 36428 14028 36484
rect 14084 36428 14094 36484
rect 19506 36428 19516 36484
rect 19572 36428 19582 36484
rect 20738 36428 20748 36484
rect 20804 36428 22540 36484
rect 22596 36428 22606 36484
rect 23314 36428 23324 36484
rect 23380 36428 24332 36484
rect 24388 36428 24398 36484
rect 26450 36428 26460 36484
rect 26516 36428 29820 36484
rect 29876 36428 30156 36484
rect 30212 36428 30222 36484
rect 19516 36372 19572 36428
rect 2818 36316 2828 36372
rect 2884 36316 5740 36372
rect 5796 36316 5806 36372
rect 13346 36316 13356 36372
rect 13412 36316 14252 36372
rect 14308 36316 14318 36372
rect 18498 36316 18508 36372
rect 18564 36316 18956 36372
rect 19012 36316 19022 36372
rect 19516 36316 21420 36372
rect 21476 36316 21486 36372
rect 26562 36316 26572 36372
rect 26628 36316 27916 36372
rect 27972 36316 27982 36372
rect 29334 36316 29372 36372
rect 29428 36316 29438 36372
rect 29894 36316 29932 36372
rect 29988 36316 29998 36372
rect 32722 36316 32732 36372
rect 32788 36316 34076 36372
rect 34132 36316 34142 36372
rect 42690 36316 42700 36372
rect 42756 36316 43260 36372
rect 43316 36316 44156 36372
rect 44212 36316 44828 36372
rect 44884 36316 46508 36372
rect 46564 36316 46574 36372
rect 11890 36204 11900 36260
rect 11956 36204 13692 36260
rect 13748 36204 13758 36260
rect 14690 36204 14700 36260
rect 14756 36204 16156 36260
rect 16212 36204 16222 36260
rect 16370 36204 16380 36260
rect 16436 36204 18284 36260
rect 18340 36204 18844 36260
rect 18900 36204 18910 36260
rect 19180 36204 19964 36260
rect 20020 36204 20030 36260
rect 20850 36204 20860 36260
rect 20916 36204 23772 36260
rect 23828 36204 23838 36260
rect 26852 36204 28588 36260
rect 28644 36204 28924 36260
rect 28980 36204 28990 36260
rect 11900 36148 11956 36204
rect 10658 36092 10668 36148
rect 10724 36092 11956 36148
rect 13692 36148 13748 36204
rect 19180 36148 19236 36204
rect 13692 36092 18788 36148
rect 18946 36092 18956 36148
rect 19012 36092 19236 36148
rect 18732 36036 18788 36092
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 26852 36036 26908 36204
rect 18732 35980 19628 36036
rect 19684 35980 19694 36036
rect 20178 35980 20188 36036
rect 20244 35980 26908 36036
rect 29138 35980 29148 36036
rect 29204 35980 31052 36036
rect 31108 35980 31118 36036
rect 8530 35868 8540 35924
rect 8596 35868 8876 35924
rect 8932 35868 8942 35924
rect 13906 35868 13916 35924
rect 13972 35868 15820 35924
rect 15876 35868 18732 35924
rect 18788 35868 18798 35924
rect 21634 35868 21644 35924
rect 21700 35868 22764 35924
rect 22820 35868 22830 35924
rect 23650 35868 23660 35924
rect 23716 35868 26460 35924
rect 26516 35868 26526 35924
rect 27682 35868 27692 35924
rect 27748 35868 30940 35924
rect 30996 35868 31006 35924
rect 23660 35812 23716 35868
rect 15250 35756 15260 35812
rect 15316 35756 21700 35812
rect 22194 35756 22204 35812
rect 22260 35756 23716 35812
rect 24098 35756 24108 35812
rect 24164 35756 25452 35812
rect 25508 35756 25518 35812
rect 29026 35756 29036 35812
rect 29092 35756 31388 35812
rect 31444 35756 31948 35812
rect 32004 35756 32014 35812
rect 32386 35756 32396 35812
rect 32452 35756 33852 35812
rect 33908 35756 33918 35812
rect 21644 35700 21700 35756
rect 8418 35644 8428 35700
rect 8484 35644 10220 35700
rect 10276 35644 11900 35700
rect 11956 35644 11966 35700
rect 18610 35644 18620 35700
rect 18676 35644 19628 35700
rect 19684 35644 19694 35700
rect 21634 35644 21644 35700
rect 21700 35644 22764 35700
rect 22820 35644 22830 35700
rect 23090 35644 23100 35700
rect 23156 35644 24556 35700
rect 24612 35644 24622 35700
rect 30370 35644 30380 35700
rect 30436 35644 31724 35700
rect 31780 35644 32284 35700
rect 32340 35644 32350 35700
rect 8866 35532 8876 35588
rect 8932 35532 10444 35588
rect 10500 35532 10510 35588
rect 15586 35532 15596 35588
rect 15652 35532 18172 35588
rect 18228 35532 20188 35588
rect 20244 35532 21084 35588
rect 21140 35532 21150 35588
rect 23426 35532 23436 35588
rect 23492 35532 26684 35588
rect 26740 35532 27468 35588
rect 27524 35532 36092 35588
rect 36148 35532 36158 35588
rect 39218 35532 39228 35588
rect 39284 35532 40572 35588
rect 40628 35532 40638 35588
rect 9874 35420 9884 35476
rect 9940 35420 10668 35476
rect 10724 35420 11228 35476
rect 11284 35420 11294 35476
rect 18386 35420 18396 35476
rect 18452 35420 23324 35476
rect 23380 35420 23390 35476
rect 28130 35420 28140 35476
rect 28196 35420 28588 35476
rect 28644 35420 29596 35476
rect 29652 35420 29662 35476
rect 29810 35420 29820 35476
rect 29876 35420 29914 35476
rect 30482 35420 30492 35476
rect 30548 35420 33740 35476
rect 33796 35420 33806 35476
rect 11330 35308 11340 35364
rect 11396 35308 13468 35364
rect 13524 35308 13534 35364
rect 19618 35308 19628 35364
rect 19684 35308 24892 35364
rect 24948 35308 24958 35364
rect 27794 35308 27804 35364
rect 27860 35308 28476 35364
rect 28532 35308 28542 35364
rect 28700 35308 29932 35364
rect 29988 35308 29998 35364
rect 33842 35308 33852 35364
rect 33908 35308 34524 35364
rect 34580 35308 34590 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 28700 35252 28756 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 18834 35196 18844 35252
rect 18900 35196 23548 35252
rect 23604 35196 23614 35252
rect 25442 35196 25452 35252
rect 25508 35196 26012 35252
rect 26068 35196 26124 35252
rect 26180 35196 26684 35252
rect 26740 35196 26750 35252
rect 27458 35196 27468 35252
rect 27524 35196 28532 35252
rect 28690 35196 28700 35252
rect 28756 35196 28766 35252
rect 28476 35140 28532 35196
rect 10882 35084 10892 35140
rect 10948 35084 11676 35140
rect 11732 35084 12124 35140
rect 12180 35084 12190 35140
rect 13794 35084 13804 35140
rect 13860 35084 14588 35140
rect 14644 35084 14654 35140
rect 19506 35084 19516 35140
rect 19572 35084 20188 35140
rect 20244 35084 20254 35140
rect 22642 35084 22652 35140
rect 22708 35084 28252 35140
rect 28308 35084 28318 35140
rect 28476 35084 29260 35140
rect 29316 35084 29932 35140
rect 29988 35084 29998 35140
rect 38210 35084 38220 35140
rect 38276 35084 38892 35140
rect 38948 35084 38958 35140
rect 10322 34972 10332 35028
rect 10388 34972 12012 35028
rect 12068 34972 12078 35028
rect 12226 34972 12236 35028
rect 12292 34972 12330 35028
rect 13346 34972 13356 35028
rect 13412 34972 14140 35028
rect 14196 34972 14206 35028
rect 16930 34972 16940 35028
rect 16996 34972 17948 35028
rect 18004 34972 18014 35028
rect 21970 34972 21980 35028
rect 22036 34972 22764 35028
rect 22820 34972 22830 35028
rect 24994 34972 25004 35028
rect 25060 34972 25396 35028
rect 25890 34972 25900 35028
rect 25956 34972 43092 35028
rect 25340 34916 25396 34972
rect 3826 34860 3836 34916
rect 3892 34860 4732 34916
rect 4788 34860 5068 34916
rect 5124 34860 10780 34916
rect 10836 34860 10846 34916
rect 11106 34860 11116 34916
rect 11172 34860 11788 34916
rect 11844 34860 11854 34916
rect 18050 34860 18060 34916
rect 18116 34860 18620 34916
rect 18676 34860 18686 34916
rect 18946 34860 18956 34916
rect 19012 34860 19628 34916
rect 19684 34860 19694 34916
rect 23874 34860 23884 34916
rect 23940 34860 25116 34916
rect 25172 34860 25182 34916
rect 25340 34860 25676 34916
rect 25732 34860 26908 34916
rect 26964 34860 26974 34916
rect 27458 34860 27468 34916
rect 27524 34860 35532 34916
rect 35588 34860 38220 34916
rect 38276 34860 38286 34916
rect 40562 34860 40572 34916
rect 40628 34860 40638 34916
rect 6738 34748 6748 34804
rect 6804 34748 7980 34804
rect 8036 34748 8046 34804
rect 12114 34748 12124 34804
rect 12180 34748 22988 34804
rect 23044 34748 23054 34804
rect 25442 34748 25452 34804
rect 25508 34748 27804 34804
rect 27860 34748 27870 34804
rect 28690 34748 28700 34804
rect 28756 34748 29820 34804
rect 29876 34748 29886 34804
rect 36082 34748 36092 34804
rect 36148 34748 37100 34804
rect 37156 34748 37166 34804
rect 40572 34692 40628 34860
rect 43036 34804 43092 34972
rect 43026 34748 43036 34804
rect 43092 34748 43102 34804
rect 8306 34636 8316 34692
rect 8372 34636 9660 34692
rect 9716 34636 9726 34692
rect 15362 34636 15372 34692
rect 15428 34636 24556 34692
rect 24612 34636 25788 34692
rect 25844 34636 34188 34692
rect 34244 34636 34254 34692
rect 37874 34636 37884 34692
rect 37940 34636 40628 34692
rect 42466 34636 42476 34692
rect 42532 34636 42924 34692
rect 42980 34636 44156 34692
rect 44212 34636 44222 34692
rect 23492 34524 29708 34580
rect 29764 34524 30828 34580
rect 30884 34524 30894 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 23492 34468 23548 34524
rect 14466 34412 14476 34468
rect 14532 34412 15372 34468
rect 15428 34412 15438 34468
rect 20626 34412 20636 34468
rect 20692 34412 21532 34468
rect 21588 34412 23212 34468
rect 23268 34412 23548 34468
rect 28466 34412 28476 34468
rect 28532 34412 28588 34468
rect 28644 34412 28812 34468
rect 28868 34412 28878 34468
rect 30258 34412 30268 34468
rect 30324 34412 31612 34468
rect 31668 34412 39004 34468
rect 39060 34412 39070 34468
rect 15026 34300 15036 34356
rect 15092 34300 17388 34356
rect 17444 34300 17454 34356
rect 18610 34300 18620 34356
rect 18676 34300 25900 34356
rect 25956 34300 25966 34356
rect 26898 34300 26908 34356
rect 26964 34300 28028 34356
rect 28084 34300 29372 34356
rect 29428 34300 29708 34356
rect 29764 34300 29774 34356
rect 39330 34300 39340 34356
rect 39396 34300 41020 34356
rect 41076 34300 42476 34356
rect 42532 34300 42542 34356
rect 5282 34188 5292 34244
rect 5348 34188 5740 34244
rect 5796 34188 5806 34244
rect 15362 34188 15372 34244
rect 15428 34188 25452 34244
rect 25508 34188 25518 34244
rect 26674 34188 26684 34244
rect 26740 34188 27804 34244
rect 27860 34188 27870 34244
rect 28802 34188 28812 34244
rect 28868 34188 31500 34244
rect 31556 34188 31566 34244
rect 33282 34188 33292 34244
rect 33348 34188 34524 34244
rect 34580 34188 34590 34244
rect 36194 34188 36204 34244
rect 36260 34188 38556 34244
rect 38612 34188 38622 34244
rect 42690 34188 42700 34244
rect 42756 34188 43932 34244
rect 43988 34188 46172 34244
rect 46228 34188 46956 34244
rect 47012 34188 47022 34244
rect 2706 34076 2716 34132
rect 2772 34076 4172 34132
rect 4228 34076 4238 34132
rect 16818 34076 16828 34132
rect 16884 34076 18956 34132
rect 19012 34076 19022 34132
rect 28018 34076 28028 34132
rect 28084 34076 29036 34132
rect 29092 34076 29102 34132
rect 29250 34076 29260 34132
rect 29316 34076 34748 34132
rect 34804 34076 34814 34132
rect 35858 34076 35868 34132
rect 35924 34076 38332 34132
rect 38388 34076 38398 34132
rect 9650 33964 9660 34020
rect 9716 33964 17276 34020
rect 17332 33964 17342 34020
rect 17826 33964 17836 34020
rect 17892 33964 19964 34020
rect 20020 33964 20030 34020
rect 25890 33964 25900 34020
rect 25956 33964 26236 34020
rect 26292 33964 26302 34020
rect 27766 33964 27804 34020
rect 27860 33964 27870 34020
rect 28914 33964 28924 34020
rect 28980 33964 30716 34020
rect 30772 33964 30782 34020
rect 31042 33964 31052 34020
rect 31108 33964 32060 34020
rect 32116 33964 32126 34020
rect 32386 33964 32396 34020
rect 32452 33964 33516 34020
rect 33572 33964 33582 34020
rect 34514 33964 34524 34020
rect 34580 33964 42140 34020
rect 42196 33964 42206 34020
rect 38612 33852 41580 33908
rect 41636 33852 41646 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 28914 33628 28924 33684
rect 28980 33628 29708 33684
rect 29764 33628 29774 33684
rect 30594 33628 30604 33684
rect 30660 33628 32508 33684
rect 32564 33628 33180 33684
rect 33236 33628 33246 33684
rect 38612 33572 38668 33852
rect 42690 33740 42700 33796
rect 42756 33740 43036 33796
rect 43092 33740 43102 33796
rect 43250 33628 43260 33684
rect 43316 33628 43326 33684
rect 43260 33572 43316 33628
rect 6066 33516 6076 33572
rect 6132 33516 8652 33572
rect 8708 33516 8988 33572
rect 9044 33516 10332 33572
rect 10388 33516 10398 33572
rect 19506 33516 19516 33572
rect 19572 33516 24556 33572
rect 24612 33516 24622 33572
rect 28130 33516 28140 33572
rect 28196 33516 33124 33572
rect 33282 33516 33292 33572
rect 33348 33516 38668 33572
rect 41234 33516 41244 33572
rect 41300 33516 41916 33572
rect 41972 33516 45276 33572
rect 45332 33516 45342 33572
rect 33068 33460 33124 33516
rect 14466 33404 14476 33460
rect 14532 33404 15596 33460
rect 15652 33404 15662 33460
rect 20514 33404 20524 33460
rect 20580 33404 24332 33460
rect 24388 33404 24398 33460
rect 27122 33404 27132 33460
rect 27188 33404 30380 33460
rect 30436 33404 30446 33460
rect 33068 33404 40012 33460
rect 40068 33404 40078 33460
rect 15810 33292 15820 33348
rect 15876 33292 19516 33348
rect 19572 33292 19582 33348
rect 20262 33292 20300 33348
rect 20356 33292 20366 33348
rect 24098 33292 24108 33348
rect 24164 33292 25340 33348
rect 25396 33292 25406 33348
rect 29922 33292 29932 33348
rect 29988 33292 30940 33348
rect 30996 33292 31006 33348
rect 35074 33292 35084 33348
rect 35140 33292 36316 33348
rect 36372 33292 36382 33348
rect 42018 33292 42028 33348
rect 42084 33292 42364 33348
rect 42420 33292 43372 33348
rect 43428 33292 43438 33348
rect 4386 33180 4396 33236
rect 4452 33180 5068 33236
rect 5124 33180 5134 33236
rect 10210 33180 10220 33236
rect 10276 33180 10668 33236
rect 10724 33180 10734 33236
rect 14018 33180 14028 33236
rect 14084 33180 15260 33236
rect 15316 33180 15326 33236
rect 16034 33180 16044 33236
rect 16100 33180 16492 33236
rect 16548 33180 16558 33236
rect 28466 33180 28476 33236
rect 28532 33180 29148 33236
rect 29204 33180 29214 33236
rect 30706 33180 30716 33236
rect 30772 33180 31724 33236
rect 31780 33180 32844 33236
rect 32900 33180 32910 33236
rect 10668 33124 10724 33180
rect 2482 33068 2492 33124
rect 2548 33068 3500 33124
rect 3556 33068 3566 33124
rect 10668 33068 17836 33124
rect 17892 33068 17902 33124
rect 19282 33068 19292 33124
rect 19348 33068 20244 33124
rect 24882 33068 24892 33124
rect 24948 33068 28140 33124
rect 28196 33068 28206 33124
rect 28914 33068 28924 33124
rect 28980 33068 31500 33124
rect 31556 33068 31566 33124
rect 32386 33068 32396 33124
rect 32452 33068 32732 33124
rect 32788 33068 32798 33124
rect 12422 32956 12460 33012
rect 12516 32956 12526 33012
rect 12870 32956 12908 33012
rect 12964 32956 12974 33012
rect 12908 32900 12964 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 20188 32900 20244 33068
rect 29362 32956 29372 33012
rect 29428 32956 29932 33012
rect 29988 32956 29998 33012
rect 10882 32844 10892 32900
rect 10948 32844 12964 32900
rect 13430 32844 13468 32900
rect 13524 32844 14364 32900
rect 14420 32844 14430 32900
rect 19170 32844 19180 32900
rect 19236 32844 19628 32900
rect 19684 32844 19694 32900
rect 20178 32844 20188 32900
rect 20244 32844 20860 32900
rect 20916 32844 20926 32900
rect 21298 32844 21308 32900
rect 21364 32844 30604 32900
rect 30660 32844 32172 32900
rect 32228 32844 32238 32900
rect 3938 32732 3948 32788
rect 4004 32732 4732 32788
rect 4788 32732 4798 32788
rect 9650 32732 9660 32788
rect 9716 32732 9996 32788
rect 10052 32732 10062 32788
rect 12002 32732 12012 32788
rect 12068 32732 32060 32788
rect 32116 32732 32126 32788
rect 41570 32732 41580 32788
rect 41636 32732 42028 32788
rect 42084 32732 43036 32788
rect 43092 32732 43102 32788
rect 8082 32620 8092 32676
rect 8148 32620 8876 32676
rect 8932 32620 10108 32676
rect 10164 32620 10174 32676
rect 12226 32620 12236 32676
rect 12292 32620 12460 32676
rect 12516 32620 12526 32676
rect 12674 32620 12684 32676
rect 12740 32620 13132 32676
rect 13188 32620 13198 32676
rect 17714 32620 17724 32676
rect 17780 32620 22092 32676
rect 22148 32620 22158 32676
rect 27878 32620 27916 32676
rect 27972 32620 27982 32676
rect 31938 32620 31948 32676
rect 32004 32620 36428 32676
rect 36484 32620 41356 32676
rect 41412 32620 41422 32676
rect 11554 32508 11564 32564
rect 11620 32508 13468 32564
rect 13524 32508 13534 32564
rect 18956 32508 21756 32564
rect 21812 32508 21822 32564
rect 26226 32508 26236 32564
rect 26292 32508 26908 32564
rect 33954 32508 33964 32564
rect 34020 32508 34030 32564
rect 38546 32508 38556 32564
rect 38612 32508 39452 32564
rect 39508 32508 39518 32564
rect 40114 32508 40124 32564
rect 40180 32508 40908 32564
rect 40964 32508 40974 32564
rect 18956 32452 19012 32508
rect 26852 32452 26908 32508
rect 33964 32452 34020 32508
rect 13346 32396 13356 32452
rect 13412 32396 15932 32452
rect 15988 32396 15998 32452
rect 17938 32396 17948 32452
rect 18004 32396 18844 32452
rect 18900 32396 18956 32452
rect 19012 32396 19022 32452
rect 20290 32396 20300 32452
rect 20356 32396 21308 32452
rect 21364 32396 21374 32452
rect 26852 32396 29596 32452
rect 29652 32396 32396 32452
rect 32452 32396 32462 32452
rect 32946 32396 32956 32452
rect 33012 32396 33628 32452
rect 33684 32396 33694 32452
rect 33964 32396 46956 32452
rect 47012 32396 47516 32452
rect 47572 32396 48300 32452
rect 48356 32396 48366 32452
rect 20626 32172 20636 32228
rect 20692 32172 26908 32228
rect 31378 32172 31388 32228
rect 31444 32172 33740 32228
rect 33796 32172 33806 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 26852 32116 26908 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 26852 32060 32284 32116
rect 32340 32060 32350 32116
rect 1810 31948 1820 32004
rect 1876 31948 6076 32004
rect 6132 31948 6142 32004
rect 39442 31948 39452 32004
rect 39508 31948 41804 32004
rect 41860 31948 41870 32004
rect 5730 31836 5740 31892
rect 5796 31836 8428 31892
rect 8484 31836 8494 31892
rect 16370 31836 16380 31892
rect 16436 31836 18508 31892
rect 18564 31836 18574 31892
rect 22642 31836 22652 31892
rect 22708 31836 23660 31892
rect 23716 31836 23726 31892
rect 32050 31836 32060 31892
rect 32116 31836 43148 31892
rect 43204 31836 43214 31892
rect 15250 31724 15260 31780
rect 15316 31724 18060 31780
rect 18116 31724 18126 31780
rect 18274 31724 18284 31780
rect 18340 31724 18732 31780
rect 18788 31724 18798 31780
rect 19954 31724 19964 31780
rect 20020 31724 21756 31780
rect 21812 31724 21822 31780
rect 22530 31724 22540 31780
rect 22596 31724 23212 31780
rect 23268 31724 27916 31780
rect 27972 31724 27982 31780
rect 32498 31724 32508 31780
rect 32564 31724 34076 31780
rect 34132 31724 34142 31780
rect 5394 31612 5404 31668
rect 5460 31612 11564 31668
rect 11620 31612 11630 31668
rect 11890 31612 11900 31668
rect 11956 31612 13580 31668
rect 13636 31612 13646 31668
rect 17714 31612 17724 31668
rect 17780 31612 19628 31668
rect 19684 31612 19694 31668
rect 20290 31612 20300 31668
rect 20356 31612 20412 31668
rect 20468 31612 20478 31668
rect 20626 31612 20636 31668
rect 20692 31612 21868 31668
rect 21924 31612 21934 31668
rect 26852 31612 31164 31668
rect 31220 31612 39564 31668
rect 39620 31612 39630 31668
rect 26852 31556 26908 31612
rect 40012 31556 40068 31836
rect 40562 31724 40572 31780
rect 40628 31724 41132 31780
rect 41188 31724 41198 31780
rect 40226 31612 40236 31668
rect 40292 31612 40908 31668
rect 40964 31612 40974 31668
rect 2482 31500 2492 31556
rect 2548 31500 3612 31556
rect 3668 31500 3678 31556
rect 17938 31500 17948 31556
rect 18004 31500 18844 31556
rect 18900 31500 18910 31556
rect 19366 31500 19404 31556
rect 19460 31500 19470 31556
rect 19628 31500 23884 31556
rect 23940 31500 25452 31556
rect 25508 31500 26908 31556
rect 30594 31500 30604 31556
rect 30660 31500 30940 31556
rect 30996 31500 31500 31556
rect 31556 31500 31566 31556
rect 32834 31500 32844 31556
rect 32900 31500 33628 31556
rect 33684 31500 33694 31556
rect 40012 31500 40572 31556
rect 40628 31500 40638 31556
rect 41346 31500 41356 31556
rect 41412 31500 42700 31556
rect 42756 31500 42766 31556
rect 19628 31444 19684 31500
rect 15362 31388 15372 31444
rect 15428 31388 19684 31444
rect 33842 31388 33852 31444
rect 33908 31388 34524 31444
rect 34580 31388 47516 31444
rect 47572 31388 48300 31444
rect 48356 31388 48366 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 15810 31164 15820 31220
rect 15876 31164 17500 31220
rect 17556 31164 17566 31220
rect 24658 31164 24668 31220
rect 24724 31164 25452 31220
rect 25508 31164 25518 31220
rect 30818 31164 30828 31220
rect 30884 31164 31724 31220
rect 31780 31164 31790 31220
rect 40338 31164 40348 31220
rect 40404 31164 40796 31220
rect 40852 31164 40862 31220
rect 41122 31164 41132 31220
rect 41188 31164 42140 31220
rect 42196 31164 42206 31220
rect 4834 31052 4844 31108
rect 4900 31052 5740 31108
rect 5796 31052 5806 31108
rect 15474 31052 15484 31108
rect 15540 31052 16604 31108
rect 16660 31052 17388 31108
rect 17444 31052 17454 31108
rect 25218 31052 25228 31108
rect 25284 31052 26460 31108
rect 26516 31052 26908 31108
rect 3938 30940 3948 30996
rect 4004 30940 5068 30996
rect 5124 30940 5134 30996
rect 6066 30940 6076 30996
rect 6132 30940 9660 30996
rect 9716 30940 11116 30996
rect 11172 30940 11182 30996
rect 12674 30940 12684 30996
rect 12740 30940 23548 30996
rect 12562 30828 12572 30884
rect 12628 30828 14588 30884
rect 14644 30828 14654 30884
rect 18050 30828 18060 30884
rect 18116 30828 19740 30884
rect 19796 30828 19806 30884
rect 23492 30772 23548 30940
rect 26852 30772 26908 31052
rect 37426 30940 37436 30996
rect 37492 30940 38668 30996
rect 38724 30940 38734 30996
rect 33618 30828 33628 30884
rect 33684 30828 40348 30884
rect 40404 30828 41468 30884
rect 41524 30828 41534 30884
rect 23492 30716 24444 30772
rect 24500 30716 25116 30772
rect 25172 30716 25182 30772
rect 26852 30716 28476 30772
rect 28532 30716 28542 30772
rect 14802 30604 14812 30660
rect 14868 30604 15372 30660
rect 15428 30604 15438 30660
rect 19058 30604 19068 30660
rect 19124 30604 25676 30660
rect 25732 30604 25742 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 17714 30492 17724 30548
rect 17780 30492 23548 30548
rect 23604 30492 24108 30548
rect 24164 30492 24174 30548
rect 12002 30380 12012 30436
rect 12068 30380 13468 30436
rect 13524 30380 14028 30436
rect 14084 30380 14094 30436
rect 43026 30380 43036 30436
rect 43092 30380 43596 30436
rect 43652 30380 43662 30436
rect 8418 30268 8428 30324
rect 8484 30268 12572 30324
rect 12628 30268 12638 30324
rect 19404 30268 19740 30324
rect 19796 30268 19806 30324
rect 22866 30268 22876 30324
rect 22932 30268 24892 30324
rect 24948 30268 24958 30324
rect 40450 30268 40460 30324
rect 40516 30268 40796 30324
rect 40852 30268 40862 30324
rect 41906 30268 41916 30324
rect 41972 30268 43148 30324
rect 43204 30268 43214 30324
rect 19404 30212 19460 30268
rect 10658 30156 10668 30212
rect 10724 30156 11676 30212
rect 11732 30156 11742 30212
rect 19394 30156 19404 30212
rect 19460 30156 19470 30212
rect 19618 30156 19628 30212
rect 19684 30156 20076 30212
rect 20132 30156 23212 30212
rect 23268 30156 23278 30212
rect 24994 30156 25004 30212
rect 25060 30156 28812 30212
rect 28868 30156 28878 30212
rect 31938 30156 31948 30212
rect 32004 30156 32284 30212
rect 32340 30156 35532 30212
rect 35588 30156 35598 30212
rect 38098 30156 38108 30212
rect 38164 30156 39060 30212
rect 39218 30156 39228 30212
rect 39284 30156 41020 30212
rect 41076 30156 41086 30212
rect 44146 30156 44156 30212
rect 44212 30156 47180 30212
rect 47236 30156 47246 30212
rect 8754 30044 8764 30100
rect 8820 30044 12236 30100
rect 12292 30044 13916 30100
rect 13972 30044 13982 30100
rect 36306 30044 36316 30100
rect 36372 30044 38668 30100
rect 38724 30044 38734 30100
rect 39004 29988 39060 30156
rect 40786 30044 40796 30100
rect 40852 30044 41244 30100
rect 41300 30044 41310 30100
rect 42354 30044 42364 30100
rect 42420 30044 43932 30100
rect 43988 30044 43998 30100
rect 18834 29932 18844 29988
rect 18900 29932 19852 29988
rect 19908 29932 20860 29988
rect 20916 29932 24556 29988
rect 24612 29932 24622 29988
rect 25890 29932 25900 29988
rect 25956 29932 26236 29988
rect 26292 29932 26302 29988
rect 39004 29932 44044 29988
rect 44100 29932 44940 29988
rect 44996 29932 45006 29988
rect 45602 29932 45612 29988
rect 45668 29932 46732 29988
rect 46788 29932 46798 29988
rect 21746 29820 21756 29876
rect 21812 29820 22428 29876
rect 22484 29820 22494 29876
rect 27010 29820 27020 29876
rect 27076 29820 27804 29876
rect 27860 29820 27870 29876
rect 38994 29820 39004 29876
rect 39060 29820 42476 29876
rect 42532 29820 42542 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 31826 29708 31836 29764
rect 31892 29708 40908 29764
rect 40964 29708 41916 29764
rect 41972 29708 41982 29764
rect 15698 29596 15708 29652
rect 15764 29596 16380 29652
rect 16436 29596 22428 29652
rect 22484 29596 22494 29652
rect 23202 29596 23212 29652
rect 23268 29596 23884 29652
rect 23940 29596 23950 29652
rect 35970 29596 35980 29652
rect 36036 29596 36764 29652
rect 36820 29596 38668 29652
rect 38612 29540 38668 29596
rect 13906 29484 13916 29540
rect 13972 29484 17276 29540
rect 17332 29484 17342 29540
rect 18162 29484 18172 29540
rect 18228 29484 18620 29540
rect 18676 29484 18686 29540
rect 19170 29484 19180 29540
rect 19236 29484 21644 29540
rect 21700 29484 21710 29540
rect 29362 29484 29372 29540
rect 29428 29484 30156 29540
rect 30212 29484 34076 29540
rect 34132 29484 34524 29540
rect 34580 29484 34590 29540
rect 38612 29484 41244 29540
rect 41300 29484 41580 29540
rect 41636 29484 41646 29540
rect 17042 29372 17052 29428
rect 17108 29372 25228 29428
rect 25284 29372 26012 29428
rect 26068 29372 33292 29428
rect 33348 29372 33358 29428
rect 39778 29372 39788 29428
rect 39844 29372 43372 29428
rect 43428 29372 46844 29428
rect 46900 29372 48300 29428
rect 48356 29372 48366 29428
rect 17798 29260 17836 29316
rect 17892 29260 17902 29316
rect 23436 29260 29484 29316
rect 29540 29260 29550 29316
rect 30482 29260 30492 29316
rect 30548 29260 31164 29316
rect 31220 29260 31230 29316
rect 33394 29260 33404 29316
rect 33460 29260 33964 29316
rect 34020 29260 36988 29316
rect 37044 29260 37054 29316
rect 12002 29148 12012 29204
rect 12068 29148 13356 29204
rect 13412 29148 13422 29204
rect 13682 29148 13692 29204
rect 13748 29148 15260 29204
rect 15316 29148 16604 29204
rect 16660 29148 16670 29204
rect 23436 29092 23492 29260
rect 24210 29148 24220 29204
rect 24276 29148 25228 29204
rect 25284 29148 25294 29204
rect 25554 29148 25564 29204
rect 25620 29148 27468 29204
rect 27524 29148 27534 29204
rect 34188 29148 38332 29204
rect 38388 29148 38398 29204
rect 18386 29036 18396 29092
rect 18452 29036 23436 29092
rect 23492 29036 23502 29092
rect 30706 29036 30716 29092
rect 30772 29036 31836 29092
rect 31892 29036 33628 29092
rect 33684 29036 33694 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 34188 28980 34244 29148
rect 36390 29036 36428 29092
rect 36484 29036 36494 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 13458 28924 13468 28980
rect 13524 28924 34188 28980
rect 34244 28924 34254 28980
rect 18918 28812 18956 28868
rect 19012 28812 19022 28868
rect 19506 28812 19516 28868
rect 19572 28812 23548 28868
rect 23604 28812 26012 28868
rect 26068 28812 26078 28868
rect 30594 28812 30604 28868
rect 30660 28812 36204 28868
rect 36260 28812 36270 28868
rect 37398 28812 37436 28868
rect 37492 28812 37502 28868
rect 38210 28812 38220 28868
rect 38276 28812 38780 28868
rect 38836 28812 38846 28868
rect 8306 28700 8316 28756
rect 8372 28700 9884 28756
rect 9940 28700 9950 28756
rect 16940 28700 17052 28756
rect 17108 28700 17388 28756
rect 17444 28700 17454 28756
rect 21644 28700 22652 28756
rect 22708 28700 25564 28756
rect 25620 28700 25630 28756
rect 29810 28700 29820 28756
rect 29876 28700 31500 28756
rect 31556 28700 31566 28756
rect 36082 28700 36092 28756
rect 36148 28700 37100 28756
rect 37156 28700 37166 28756
rect 37324 28700 39116 28756
rect 39172 28700 39182 28756
rect 16940 28644 16996 28700
rect 21644 28644 21700 28700
rect 37324 28644 37380 28700
rect 6626 28588 6636 28644
rect 6692 28588 8204 28644
rect 8260 28588 8270 28644
rect 8978 28588 8988 28644
rect 9044 28588 9772 28644
rect 9828 28588 9838 28644
rect 14354 28588 14364 28644
rect 14420 28588 14924 28644
rect 14980 28588 14990 28644
rect 16930 28588 16940 28644
rect 16996 28588 17006 28644
rect 19282 28588 19292 28644
rect 19348 28588 19740 28644
rect 19796 28588 19806 28644
rect 20748 28588 21700 28644
rect 23650 28588 23660 28644
rect 23716 28588 25004 28644
rect 25060 28588 25070 28644
rect 29474 28588 29484 28644
rect 29540 28588 30156 28644
rect 30212 28588 30222 28644
rect 32610 28588 32620 28644
rect 32676 28588 37380 28644
rect 38658 28588 38668 28644
rect 38724 28588 38892 28644
rect 38948 28588 45500 28644
rect 45556 28588 46284 28644
rect 46340 28588 46350 28644
rect 46722 28588 46732 28644
rect 46788 28588 46956 28644
rect 47012 28588 47964 28644
rect 48020 28588 48030 28644
rect 20748 28532 20804 28588
rect 21644 28532 21700 28588
rect 8642 28476 8652 28532
rect 8708 28476 10332 28532
rect 10388 28476 16156 28532
rect 16212 28476 16222 28532
rect 20738 28476 20748 28532
rect 20804 28476 20814 28532
rect 21634 28476 21644 28532
rect 21700 28476 21710 28532
rect 24098 28476 24108 28532
rect 24164 28476 25452 28532
rect 25508 28476 25518 28532
rect 33618 28476 33628 28532
rect 33684 28476 33964 28532
rect 34020 28476 34524 28532
rect 34580 28476 35196 28532
rect 35252 28476 35262 28532
rect 39330 28476 39340 28532
rect 39396 28476 40236 28532
rect 40292 28476 41132 28532
rect 41188 28476 41198 28532
rect 16930 28364 16940 28420
rect 16996 28364 18508 28420
rect 18564 28364 18574 28420
rect 20626 28364 20636 28420
rect 20692 28364 21980 28420
rect 22036 28364 22046 28420
rect 23874 28364 23884 28420
rect 23940 28364 24668 28420
rect 24724 28364 24734 28420
rect 30370 28364 30380 28420
rect 30436 28364 31164 28420
rect 31220 28364 31230 28420
rect 14802 28252 14812 28308
rect 14868 28252 14878 28308
rect 5170 28028 5180 28084
rect 5236 28028 9660 28084
rect 9716 28028 10780 28084
rect 10836 28028 10846 28084
rect 14812 27972 14868 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 27346 28140 27356 28196
rect 27412 28140 29932 28196
rect 29988 28140 38556 28196
rect 38612 28140 38622 28196
rect 44034 28140 44044 28196
rect 44100 28140 46396 28196
rect 46452 28140 46462 28196
rect 17714 28028 17724 28084
rect 17780 28028 18620 28084
rect 18676 28028 18844 28084
rect 18900 28028 18910 28084
rect 19058 28028 19068 28084
rect 19124 28028 19404 28084
rect 19460 28028 22428 28084
rect 22484 28028 23660 28084
rect 23716 28028 24108 28084
rect 24164 28028 24332 28084
rect 24388 28028 24398 28084
rect 27010 28028 27020 28084
rect 27076 28028 31948 28084
rect 32004 28028 32014 28084
rect 32274 28028 32284 28084
rect 32340 28028 34860 28084
rect 34916 28028 34926 28084
rect 35084 28028 39228 28084
rect 39284 28028 39294 28084
rect 43026 28028 43036 28084
rect 43092 28028 45500 28084
rect 45556 28028 45566 28084
rect 32284 27972 32340 28028
rect 13570 27916 13580 27972
rect 13636 27916 14140 27972
rect 14196 27916 14206 27972
rect 14466 27916 14476 27972
rect 14532 27916 14868 27972
rect 27682 27916 27692 27972
rect 27748 27916 28028 27972
rect 28084 27916 28094 27972
rect 30594 27916 30604 27972
rect 30660 27916 32340 27972
rect 2818 27804 2828 27860
rect 2884 27804 4060 27860
rect 4116 27804 4126 27860
rect 14812 27748 14868 27916
rect 16818 27804 16828 27860
rect 16884 27804 19516 27860
rect 19572 27804 19582 27860
rect 26852 27804 27468 27860
rect 27524 27804 27534 27860
rect 26852 27748 26908 27804
rect 35084 27748 35140 28028
rect 37986 27916 37996 27972
rect 38052 27916 40908 27972
rect 40964 27916 41580 27972
rect 41636 27916 41646 27972
rect 43586 27916 43596 27972
rect 43652 27916 46060 27972
rect 46116 27916 46126 27972
rect 14812 27692 18508 27748
rect 18564 27692 18574 27748
rect 26114 27692 26124 27748
rect 26180 27692 26908 27748
rect 27570 27692 27580 27748
rect 27636 27692 35140 27748
rect 16706 27580 16716 27636
rect 16772 27580 17724 27636
rect 17780 27580 17790 27636
rect 25974 27580 26012 27636
rect 26068 27580 26078 27636
rect 30930 27580 30940 27636
rect 30996 27580 32172 27636
rect 32228 27580 35588 27636
rect 7858 27468 7868 27524
rect 7924 27468 9212 27524
rect 9268 27468 10108 27524
rect 10164 27468 10174 27524
rect 14578 27468 14588 27524
rect 14644 27468 15036 27524
rect 15092 27468 15102 27524
rect 21746 27468 21756 27524
rect 21812 27468 30044 27524
rect 30100 27468 30110 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 35532 27412 35588 27580
rect 37996 27524 38052 27916
rect 41010 27804 41020 27860
rect 41076 27804 44716 27860
rect 44772 27804 44782 27860
rect 40338 27692 40348 27748
rect 40404 27692 42700 27748
rect 42756 27692 42766 27748
rect 38882 27580 38892 27636
rect 38948 27580 39564 27636
rect 39620 27580 39630 27636
rect 37650 27468 37660 27524
rect 37716 27468 38052 27524
rect 42354 27468 42364 27524
rect 42420 27468 43484 27524
rect 43540 27468 43550 27524
rect 9314 27356 9324 27412
rect 9380 27356 9884 27412
rect 9940 27356 10780 27412
rect 10836 27356 10846 27412
rect 33506 27356 33516 27412
rect 33572 27356 33852 27412
rect 33908 27356 34188 27412
rect 34244 27356 34254 27412
rect 35532 27356 39788 27412
rect 39844 27356 39854 27412
rect 40002 27356 40012 27412
rect 40068 27356 43036 27412
rect 43092 27356 43102 27412
rect 10098 27244 10108 27300
rect 10164 27244 12348 27300
rect 12404 27244 12414 27300
rect 12562 27244 12572 27300
rect 12628 27244 22092 27300
rect 22148 27244 22540 27300
rect 22596 27244 22606 27300
rect 23202 27244 23212 27300
rect 23268 27244 24444 27300
rect 24500 27244 24510 27300
rect 25666 27244 25676 27300
rect 25732 27244 26572 27300
rect 26628 27244 26638 27300
rect 26852 27244 30940 27300
rect 30996 27244 38892 27300
rect 38948 27244 38958 27300
rect 40674 27244 40684 27300
rect 40740 27244 45836 27300
rect 45892 27244 45902 27300
rect 26852 27188 26908 27244
rect 7634 27132 7644 27188
rect 7700 27132 8204 27188
rect 8260 27132 13580 27188
rect 13636 27132 14476 27188
rect 14532 27132 14542 27188
rect 14914 27132 14924 27188
rect 14980 27132 15018 27188
rect 15092 27132 17612 27188
rect 17668 27132 17678 27188
rect 19394 27132 19404 27188
rect 19460 27132 19628 27188
rect 19684 27132 20020 27188
rect 20850 27132 20860 27188
rect 20916 27132 21756 27188
rect 21812 27132 26908 27188
rect 31798 27132 31836 27188
rect 31892 27132 31902 27188
rect 32946 27132 32956 27188
rect 33012 27132 33852 27188
rect 33908 27132 33918 27188
rect 36978 27132 36988 27188
rect 37044 27132 38444 27188
rect 38500 27132 38510 27188
rect 41458 27132 41468 27188
rect 41524 27132 42700 27188
rect 42756 27132 44156 27188
rect 44212 27132 45388 27188
rect 45444 27132 45454 27188
rect 4162 27020 4172 27076
rect 4228 27020 5628 27076
rect 5684 27020 5694 27076
rect 8082 27020 8092 27076
rect 8148 27020 9436 27076
rect 9492 27020 9502 27076
rect 12002 27020 12012 27076
rect 12068 27020 12572 27076
rect 12628 27020 12638 27076
rect 15026 27020 15036 27076
rect 15092 27020 15148 27132
rect 19964 27076 20020 27132
rect 17714 27020 17724 27076
rect 17780 27020 19740 27076
rect 19796 27020 19806 27076
rect 19964 27020 20748 27076
rect 20804 27020 20814 27076
rect 23492 27020 31276 27076
rect 31332 27020 32508 27076
rect 32564 27020 33180 27076
rect 33236 27020 33246 27076
rect 39442 27020 39452 27076
rect 39508 27020 40124 27076
rect 40180 27020 40190 27076
rect 42242 27020 42252 27076
rect 42308 27020 45612 27076
rect 45668 27020 45678 27076
rect 5628 26964 5684 27020
rect 2594 26908 2604 26964
rect 2660 26908 3836 26964
rect 3892 26908 3902 26964
rect 5628 26908 8876 26964
rect 8932 26908 9996 26964
rect 10052 26908 10062 26964
rect 11106 26908 11116 26964
rect 11172 26908 12684 26964
rect 12740 26908 15372 26964
rect 15428 26908 15438 26964
rect 17154 26908 17164 26964
rect 17220 26908 17500 26964
rect 17556 26908 18900 26964
rect 20076 26908 21308 26964
rect 21364 26908 21374 26964
rect 18844 26852 19012 26908
rect 20076 26852 20132 26908
rect 18956 26796 20132 26852
rect 20188 26796 21532 26852
rect 21588 26796 21598 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 20188 26628 20244 26796
rect 21522 26684 21532 26740
rect 21588 26684 21756 26740
rect 21812 26684 21822 26740
rect 23492 26628 23548 27020
rect 31826 26908 31836 26964
rect 31892 26908 37212 26964
rect 37268 26908 37278 26964
rect 39778 26908 39788 26964
rect 39844 26908 41244 26964
rect 41300 26908 41310 26964
rect 43362 26908 43372 26964
rect 43428 26908 43820 26964
rect 43876 26908 45276 26964
rect 45332 26908 45342 26964
rect 30818 26796 30828 26852
rect 30884 26796 31164 26852
rect 31220 26796 31230 26852
rect 39666 26796 39676 26852
rect 39732 26796 40908 26852
rect 40964 26796 40974 26852
rect 28466 26684 28476 26740
rect 28532 26684 33516 26740
rect 33572 26684 33582 26740
rect 38612 26684 40348 26740
rect 40404 26684 41916 26740
rect 41972 26684 41982 26740
rect 20178 26572 20188 26628
rect 20244 26572 20254 26628
rect 20710 26572 20748 26628
rect 20804 26572 23548 26628
rect 38612 26516 38668 26684
rect 22166 26460 22204 26516
rect 22260 26460 22270 26516
rect 30034 26460 30044 26516
rect 30100 26460 38668 26516
rect 9538 26348 9548 26404
rect 9604 26348 10108 26404
rect 10164 26348 10668 26404
rect 10724 26348 33180 26404
rect 33236 26348 33516 26404
rect 33572 26348 33582 26404
rect 35298 26348 35308 26404
rect 35364 26348 36988 26404
rect 37044 26348 37324 26404
rect 37380 26348 37390 26404
rect 5170 26236 5180 26292
rect 5236 26236 5740 26292
rect 5796 26236 8764 26292
rect 8820 26236 8830 26292
rect 12338 26236 12348 26292
rect 12404 26236 13804 26292
rect 13860 26236 13870 26292
rect 14466 26236 14476 26292
rect 14532 26236 14924 26292
rect 14980 26236 14990 26292
rect 26852 26236 27916 26292
rect 27972 26236 40236 26292
rect 40292 26236 40302 26292
rect 43026 26236 43036 26292
rect 43092 26236 44268 26292
rect 44324 26236 44334 26292
rect 9846 26124 9884 26180
rect 9940 26124 9950 26180
rect 17378 26124 17388 26180
rect 17444 26124 19292 26180
rect 19348 26124 25620 26180
rect 25564 26068 25620 26124
rect 26852 26068 26908 26236
rect 34402 26124 34412 26180
rect 34468 26124 41468 26180
rect 41524 26124 41534 26180
rect 2034 26012 2044 26068
rect 2100 26012 25228 26068
rect 25284 26012 25294 26068
rect 25564 26012 26908 26068
rect 38612 26012 47740 26068
rect 47796 26012 47806 26068
rect 9650 25900 9660 25956
rect 9716 25900 11116 25956
rect 11172 25900 11182 25956
rect 14018 25900 14028 25956
rect 14084 25900 14476 25956
rect 14532 25900 14542 25956
rect 14886 25900 14924 25956
rect 14980 25900 14990 25956
rect 18274 25900 18284 25956
rect 18340 25900 25564 25956
rect 25620 25900 25630 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 15362 25788 15372 25844
rect 15428 25788 26572 25844
rect 26628 25788 26638 25844
rect 29362 25788 29372 25844
rect 29428 25788 30044 25844
rect 30100 25788 30110 25844
rect 30790 25788 30828 25844
rect 30884 25788 30894 25844
rect 38612 25732 38668 26012
rect 40786 25900 40796 25956
rect 40852 25900 40862 25956
rect 24546 25676 24556 25732
rect 24612 25676 27132 25732
rect 27188 25676 28252 25732
rect 28308 25676 38668 25732
rect 40796 25620 40852 25900
rect 11732 25564 12012 25620
rect 12068 25564 18060 25620
rect 18116 25564 18126 25620
rect 18722 25564 18732 25620
rect 18788 25564 19740 25620
rect 19796 25564 20300 25620
rect 20356 25564 20366 25620
rect 22194 25564 22204 25620
rect 22260 25564 23100 25620
rect 23156 25564 23166 25620
rect 26898 25564 26908 25620
rect 26964 25564 27860 25620
rect 28018 25564 28028 25620
rect 28084 25564 40852 25620
rect 45378 25564 45388 25620
rect 45444 25564 46508 25620
rect 46564 25564 46574 25620
rect 9174 25452 9212 25508
rect 9268 25452 9278 25508
rect 11732 25396 11788 25564
rect 27804 25508 27860 25564
rect 12898 25452 12908 25508
rect 12964 25452 13580 25508
rect 13636 25452 13646 25508
rect 18386 25452 18396 25508
rect 18452 25452 19964 25508
rect 20020 25452 22428 25508
rect 22484 25452 23772 25508
rect 23828 25452 24500 25508
rect 26562 25452 26572 25508
rect 26628 25452 27580 25508
rect 27636 25452 27646 25508
rect 27804 25452 28140 25508
rect 28196 25452 28206 25508
rect 28578 25452 28588 25508
rect 28644 25452 29820 25508
rect 29876 25452 29886 25508
rect 30258 25452 30268 25508
rect 30324 25452 31500 25508
rect 31556 25452 31566 25508
rect 31826 25452 31836 25508
rect 31892 25452 35756 25508
rect 35812 25452 35822 25508
rect 24444 25396 24500 25452
rect 11554 25340 11564 25396
rect 11620 25340 11788 25396
rect 18834 25340 18844 25396
rect 18900 25340 19292 25396
rect 19348 25340 21308 25396
rect 21364 25340 22988 25396
rect 23044 25340 23996 25396
rect 24052 25340 24062 25396
rect 24434 25340 24444 25396
rect 24500 25340 24510 25396
rect 26226 25340 26236 25396
rect 26292 25340 31612 25396
rect 31668 25340 32732 25396
rect 32788 25340 32798 25396
rect 46946 25340 46956 25396
rect 47012 25340 48300 25396
rect 48356 25340 48366 25396
rect 8642 25228 8652 25284
rect 8708 25228 13804 25284
rect 13860 25228 14812 25284
rect 14868 25228 14878 25284
rect 16146 25228 16156 25284
rect 16212 25228 17388 25284
rect 17444 25228 17454 25284
rect 18060 25228 19180 25284
rect 19236 25228 19246 25284
rect 19842 25228 19852 25284
rect 19908 25228 21532 25284
rect 21588 25228 22204 25284
rect 22260 25228 22270 25284
rect 26114 25228 26124 25284
rect 26180 25228 27692 25284
rect 27748 25228 27758 25284
rect 27906 25228 27916 25284
rect 27972 25228 28028 25284
rect 28084 25228 28094 25284
rect 31154 25228 31164 25284
rect 31220 25228 32172 25284
rect 32228 25228 32620 25284
rect 32676 25228 32686 25284
rect 42018 25228 42028 25284
rect 42084 25228 44940 25284
rect 44996 25228 45006 25284
rect 18060 25060 18116 25228
rect 26338 25116 26348 25172
rect 26404 25116 26796 25172
rect 26852 25116 26862 25172
rect 27010 25116 27020 25172
rect 27076 25116 27468 25172
rect 27524 25116 27534 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 9874 25004 9884 25060
rect 9940 25004 10500 25060
rect 18050 25004 18060 25060
rect 18116 25004 18126 25060
rect 21494 25004 21532 25060
rect 21588 25004 21598 25060
rect 21746 25004 21756 25060
rect 21812 25004 21850 25060
rect 10444 24836 10500 25004
rect 10994 24892 11004 24948
rect 11060 24892 11340 24948
rect 11396 24892 11406 24948
rect 11890 24892 11900 24948
rect 11956 24892 12460 24948
rect 12516 24892 12526 24948
rect 13458 24892 13468 24948
rect 13524 24892 14252 24948
rect 14308 24892 14318 24948
rect 19058 24892 19068 24948
rect 19124 24892 20748 24948
rect 20804 24892 20814 24948
rect 21858 24892 21868 24948
rect 21924 24892 22204 24948
rect 22260 24892 22270 24948
rect 26786 24892 26796 24948
rect 26852 24892 28812 24948
rect 28868 24892 29148 24948
rect 29204 24892 29214 24948
rect 9090 24780 9100 24836
rect 9156 24780 9884 24836
rect 9940 24780 9950 24836
rect 10444 24780 10556 24836
rect 10612 24780 10622 24836
rect 24210 24780 24220 24836
rect 24276 24780 26348 24836
rect 26404 24780 26414 24836
rect 37874 24780 37884 24836
rect 37940 24780 38556 24836
rect 38612 24780 38622 24836
rect 8530 24668 8540 24724
rect 8596 24668 8988 24724
rect 9044 24668 9660 24724
rect 9716 24668 11340 24724
rect 11396 24668 14700 24724
rect 14756 24668 14766 24724
rect 24994 24668 25004 24724
rect 25060 24668 29148 24724
rect 29204 24668 29708 24724
rect 29764 24668 29774 24724
rect 32274 24668 32284 24724
rect 32340 24668 34524 24724
rect 34580 24668 36540 24724
rect 36596 24668 36606 24724
rect 37426 24668 37436 24724
rect 37492 24668 38780 24724
rect 38836 24668 38846 24724
rect 41122 24668 41132 24724
rect 41188 24668 42140 24724
rect 42196 24668 43036 24724
rect 43092 24668 43102 24724
rect 5618 24556 5628 24612
rect 5684 24556 8316 24612
rect 8372 24556 9492 24612
rect 12422 24556 12460 24612
rect 12516 24556 12526 24612
rect 13430 24556 13468 24612
rect 13524 24556 13534 24612
rect 27570 24556 27580 24612
rect 27636 24556 28252 24612
rect 28308 24556 31836 24612
rect 31892 24556 39340 24612
rect 39396 24556 39406 24612
rect 9436 24500 9492 24556
rect 9426 24444 9436 24500
rect 9492 24444 9502 24500
rect 14354 24444 14364 24500
rect 14420 24444 14700 24500
rect 14756 24444 14766 24500
rect 26226 24444 26236 24500
rect 26292 24444 27804 24500
rect 27860 24444 27870 24500
rect 30156 24444 31164 24500
rect 31220 24444 31230 24500
rect 32498 24444 32508 24500
rect 32564 24444 34188 24500
rect 34244 24444 34748 24500
rect 34804 24444 34814 24500
rect 34972 24444 38668 24500
rect 30156 24388 30212 24444
rect 34972 24388 35028 24444
rect 12674 24332 12684 24388
rect 12740 24332 13356 24388
rect 13412 24332 13422 24388
rect 18162 24332 18172 24388
rect 18228 24332 30212 24388
rect 30370 24332 30380 24388
rect 30436 24332 31276 24388
rect 31332 24332 31948 24388
rect 32004 24332 35028 24388
rect 36082 24332 36092 24388
rect 36148 24332 38444 24388
rect 38500 24332 38510 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 9762 24220 9772 24276
rect 9828 24220 10444 24276
rect 10500 24220 21028 24276
rect 20972 24164 21028 24220
rect 26796 24220 27468 24276
rect 27524 24220 27534 24276
rect 28354 24220 28364 24276
rect 28420 24220 29596 24276
rect 29652 24220 30044 24276
rect 30100 24220 30492 24276
rect 30548 24220 30558 24276
rect 36194 24220 36204 24276
rect 36260 24220 38332 24276
rect 38388 24220 38398 24276
rect 26796 24164 26852 24220
rect 38612 24164 38668 24444
rect 12114 24108 12124 24164
rect 12180 24108 16380 24164
rect 16436 24108 16446 24164
rect 20972 24108 26796 24164
rect 26852 24108 26862 24164
rect 27346 24108 27356 24164
rect 27412 24108 31948 24164
rect 32004 24108 36988 24164
rect 37044 24108 37054 24164
rect 38612 24108 39788 24164
rect 39844 24108 39854 24164
rect 7746 23996 7756 24052
rect 7812 23996 9884 24052
rect 9940 23996 13580 24052
rect 13636 23996 14140 24052
rect 14196 23996 15036 24052
rect 15092 23996 15102 24052
rect 32610 23996 32620 24052
rect 32676 23996 33852 24052
rect 33908 23996 33918 24052
rect 36418 23996 36428 24052
rect 36484 23996 36494 24052
rect 36614 23996 36652 24052
rect 36708 23996 36718 24052
rect 36428 23940 36484 23996
rect 4162 23884 4172 23940
rect 4228 23884 9996 23940
rect 10052 23884 10062 23940
rect 11218 23884 11228 23940
rect 11284 23884 12124 23940
rect 12180 23884 12190 23940
rect 12674 23884 12684 23940
rect 12740 23884 12908 23940
rect 12964 23884 12974 23940
rect 20178 23884 20188 23940
rect 20244 23884 20860 23940
rect 20916 23884 21644 23940
rect 21700 23884 23324 23940
rect 23380 23884 23390 23940
rect 26852 23884 27020 23940
rect 27076 23884 27086 23940
rect 29138 23884 29148 23940
rect 29204 23884 29214 23940
rect 33170 23884 33180 23940
rect 33236 23884 39452 23940
rect 39508 23884 39900 23940
rect 39956 23884 42028 23940
rect 42084 23884 42094 23940
rect 46162 23884 46172 23940
rect 46228 23884 47180 23940
rect 47236 23884 48412 23940
rect 48468 23884 48478 23940
rect 2930 23772 2940 23828
rect 2996 23772 3836 23828
rect 3892 23772 3902 23828
rect 4834 23772 4844 23828
rect 4900 23772 8988 23828
rect 9044 23772 9054 23828
rect 9314 23772 9324 23828
rect 9380 23772 9884 23828
rect 9940 23772 9950 23828
rect 15474 23772 15484 23828
rect 15540 23772 17724 23828
rect 17780 23772 17790 23828
rect 18844 23772 26796 23828
rect 26852 23772 26908 23884
rect 18844 23716 18900 23772
rect 29148 23716 29204 23884
rect 37538 23772 37548 23828
rect 37604 23772 37996 23828
rect 38052 23772 38556 23828
rect 38612 23772 38622 23828
rect 12898 23660 12908 23716
rect 12964 23660 14476 23716
rect 14532 23660 14542 23716
rect 14690 23660 14700 23716
rect 14756 23660 17164 23716
rect 17220 23660 17388 23716
rect 17444 23660 17454 23716
rect 17602 23660 17612 23716
rect 17668 23660 18900 23716
rect 22530 23660 22540 23716
rect 22596 23660 24668 23716
rect 24724 23660 24734 23716
rect 25218 23660 25228 23716
rect 25284 23660 26236 23716
rect 26292 23660 29204 23716
rect 32162 23660 32172 23716
rect 32228 23660 32396 23716
rect 32452 23660 36204 23716
rect 36260 23660 36270 23716
rect 38434 23660 38444 23716
rect 38500 23660 47292 23716
rect 47348 23660 47358 23716
rect 17612 23604 17668 23660
rect 9174 23548 9212 23604
rect 9268 23548 9278 23604
rect 16706 23548 16716 23604
rect 16772 23548 17668 23604
rect 20402 23548 20412 23604
rect 20468 23548 23324 23604
rect 23380 23548 23390 23604
rect 24322 23548 24332 23604
rect 24388 23548 36092 23604
rect 36148 23548 36158 23604
rect 39666 23548 39676 23604
rect 39732 23548 41972 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 36390 23492 36428 23548
rect 36484 23492 36494 23548
rect 41916 23492 41972 23548
rect 10210 23436 10220 23492
rect 10276 23436 10668 23492
rect 10724 23436 17948 23492
rect 18004 23436 18014 23492
rect 41906 23436 41916 23492
rect 41972 23436 43596 23492
rect 43652 23436 43662 23492
rect 9090 23324 9100 23380
rect 9156 23324 9548 23380
rect 9604 23324 9614 23380
rect 17490 23324 17500 23380
rect 17556 23324 20188 23380
rect 20244 23324 20254 23380
rect 22194 23324 22204 23380
rect 22260 23324 23100 23380
rect 23156 23324 23166 23380
rect 30034 23324 30044 23380
rect 30100 23324 31388 23380
rect 31444 23324 31454 23380
rect 32610 23324 32620 23380
rect 32676 23324 33292 23380
rect 33348 23324 34076 23380
rect 34132 23324 34142 23380
rect 38612 23324 38780 23380
rect 38836 23324 38846 23380
rect 4946 23212 4956 23268
rect 5012 23212 5852 23268
rect 5908 23212 6300 23268
rect 6356 23212 6366 23268
rect 9762 23212 9772 23268
rect 9828 23212 10892 23268
rect 10948 23212 10958 23268
rect 18162 23212 18172 23268
rect 18228 23212 20636 23268
rect 20692 23212 20702 23268
rect 28802 23212 28812 23268
rect 28868 23212 30492 23268
rect 30548 23212 30558 23268
rect 38612 23156 38668 23324
rect 41346 23212 41356 23268
rect 41412 23212 41692 23268
rect 41748 23212 44716 23268
rect 44772 23212 47628 23268
rect 47684 23212 47694 23268
rect 4722 23100 4732 23156
rect 4788 23100 5516 23156
rect 5572 23100 6412 23156
rect 6468 23100 10108 23156
rect 10164 23100 10174 23156
rect 11666 23100 11676 23156
rect 11732 23100 12124 23156
rect 12180 23100 13468 23156
rect 13524 23100 13534 23156
rect 16930 23100 16940 23156
rect 16996 23100 17388 23156
rect 17444 23100 17454 23156
rect 18946 23100 18956 23156
rect 19012 23100 19740 23156
rect 19796 23100 38668 23156
rect 40114 23100 40124 23156
rect 40180 23100 41020 23156
rect 41076 23100 41086 23156
rect 11330 22988 11340 23044
rect 11396 22988 11788 23044
rect 11844 22988 12572 23044
rect 12628 22988 25228 23044
rect 25284 22988 25294 23044
rect 27458 22988 27468 23044
rect 27524 22988 29372 23044
rect 29428 22988 31724 23044
rect 31780 22988 37884 23044
rect 37940 22988 37950 23044
rect 2594 22876 2604 22932
rect 2660 22876 5292 22932
rect 5348 22876 5358 22932
rect 26002 22876 26012 22932
rect 26068 22876 26460 22932
rect 26516 22876 26526 22932
rect 28130 22876 28140 22932
rect 28196 22876 31836 22932
rect 31892 22876 32508 22932
rect 32564 22876 36764 22932
rect 36820 22876 37324 22932
rect 37380 22876 37390 22932
rect 13122 22764 13132 22820
rect 13188 22764 13916 22820
rect 13972 22764 17500 22820
rect 17556 22764 17566 22820
rect 25218 22764 25228 22820
rect 25284 22764 34412 22820
rect 34468 22764 34478 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 27346 22652 27356 22708
rect 27412 22652 27916 22708
rect 27972 22652 27982 22708
rect 31042 22652 31052 22708
rect 31108 22652 31836 22708
rect 31892 22652 31902 22708
rect 36978 22652 36988 22708
rect 37044 22652 37996 22708
rect 38052 22652 38062 22708
rect 8194 22540 8204 22596
rect 8260 22540 9212 22596
rect 9268 22540 9996 22596
rect 10052 22540 10062 22596
rect 12786 22540 12796 22596
rect 12852 22540 24220 22596
rect 24276 22540 24286 22596
rect 1922 22428 1932 22484
rect 1988 22428 3388 22484
rect 10210 22428 10220 22484
rect 10276 22428 11564 22484
rect 11620 22428 12908 22484
rect 12964 22428 12974 22484
rect 14914 22428 14924 22484
rect 14980 22428 17388 22484
rect 17444 22428 21308 22484
rect 21364 22428 21374 22484
rect 23426 22428 23436 22484
rect 23492 22428 26572 22484
rect 26628 22428 29372 22484
rect 29428 22428 29438 22484
rect 29698 22428 29708 22484
rect 29764 22428 30044 22484
rect 30100 22428 30110 22484
rect 42018 22428 42028 22484
rect 42084 22428 43260 22484
rect 43316 22428 44492 22484
rect 44548 22428 44940 22484
rect 44996 22428 45006 22484
rect 3332 22372 3388 22428
rect 3332 22316 4956 22372
rect 5012 22316 5740 22372
rect 5796 22316 6524 22372
rect 6580 22316 6590 22372
rect 12450 22316 12460 22372
rect 12516 22316 16492 22372
rect 16548 22316 16558 22372
rect 18274 22316 18284 22372
rect 18340 22316 21980 22372
rect 22036 22316 22046 22372
rect 30370 22316 30380 22372
rect 30436 22316 33964 22372
rect 34020 22316 36204 22372
rect 36260 22316 36270 22372
rect 9650 22204 9660 22260
rect 9716 22204 10108 22260
rect 10164 22204 10174 22260
rect 14018 22204 14028 22260
rect 14084 22204 18172 22260
rect 18228 22204 18238 22260
rect 19506 22204 19516 22260
rect 19572 22204 20860 22260
rect 20916 22204 20926 22260
rect 29586 22204 29596 22260
rect 29652 22204 30716 22260
rect 30772 22204 30782 22260
rect 32722 22204 32732 22260
rect 32788 22204 33740 22260
rect 33796 22204 34860 22260
rect 34916 22204 34926 22260
rect 44034 22204 44044 22260
rect 44100 22204 45164 22260
rect 45220 22204 45230 22260
rect 5730 22092 5740 22148
rect 5796 22092 6188 22148
rect 6244 22092 6972 22148
rect 7028 22092 7038 22148
rect 16258 22092 16268 22148
rect 16324 22092 18396 22148
rect 18452 22092 18462 22148
rect 20626 22092 20636 22148
rect 20692 22092 28700 22148
rect 28756 22092 39004 22148
rect 39060 22092 39070 22148
rect 39442 22092 39452 22148
rect 39508 22092 39788 22148
rect 39844 22092 40460 22148
rect 40516 22092 41132 22148
rect 41188 22092 41198 22148
rect 44258 22092 44268 22148
rect 44324 22092 45500 22148
rect 45556 22092 45566 22148
rect 22530 21980 22540 22036
rect 22596 21980 22988 22036
rect 23044 21980 23436 22036
rect 23492 21980 27244 22036
rect 27300 21980 27804 22036
rect 27860 21980 27870 22036
rect 31714 21980 31724 22036
rect 31780 21980 33068 22036
rect 33124 21980 33134 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 9874 21868 9884 21924
rect 9940 21868 14924 21924
rect 14980 21868 14990 21924
rect 36082 21868 36092 21924
rect 36148 21868 37212 21924
rect 37268 21868 37278 21924
rect 13010 21756 13020 21812
rect 13076 21756 13580 21812
rect 13636 21756 13646 21812
rect 14354 21756 14364 21812
rect 14420 21756 17724 21812
rect 17780 21756 27132 21812
rect 27188 21756 27412 21812
rect 27570 21756 27580 21812
rect 27636 21756 30604 21812
rect 30660 21756 30670 21812
rect 32162 21756 32172 21812
rect 32228 21756 34076 21812
rect 34132 21756 34142 21812
rect 34402 21756 34412 21812
rect 34468 21756 36316 21812
rect 36372 21756 36382 21812
rect 10322 21644 10332 21700
rect 10388 21644 11116 21700
rect 11172 21644 14028 21700
rect 14084 21644 14094 21700
rect 19058 21644 19068 21700
rect 19124 21644 20300 21700
rect 20356 21644 21084 21700
rect 21140 21644 22204 21700
rect 22260 21644 23772 21700
rect 23828 21644 23838 21700
rect 24658 21644 24668 21700
rect 24724 21644 25452 21700
rect 25508 21644 26796 21700
rect 26852 21644 26908 21700
rect 26964 21644 26974 21700
rect 27356 21588 27412 21756
rect 28690 21644 28700 21700
rect 28756 21644 29708 21700
rect 29764 21644 29774 21700
rect 32274 21644 32284 21700
rect 32340 21644 32508 21700
rect 32564 21644 32574 21700
rect 36866 21644 36876 21700
rect 36932 21644 37772 21700
rect 37828 21644 38444 21700
rect 38500 21644 38510 21700
rect 39442 21644 39452 21700
rect 39508 21644 40124 21700
rect 40180 21644 40190 21700
rect 41458 21644 41468 21700
rect 41524 21644 41804 21700
rect 41860 21644 42812 21700
rect 42868 21644 42878 21700
rect 45938 21644 45948 21700
rect 46004 21644 47964 21700
rect 48020 21644 48030 21700
rect 32284 21588 32340 21644
rect 39452 21588 39508 21644
rect 4834 21532 4844 21588
rect 4900 21532 6412 21588
rect 6468 21532 9772 21588
rect 9828 21532 9838 21588
rect 26450 21532 26460 21588
rect 26516 21532 26628 21588
rect 27356 21532 28028 21588
rect 28084 21532 29596 21588
rect 29652 21532 29662 21588
rect 31490 21532 31500 21588
rect 31556 21532 32340 21588
rect 34514 21532 34524 21588
rect 34580 21532 35756 21588
rect 35812 21532 35822 21588
rect 37426 21532 37436 21588
rect 37492 21532 38668 21588
rect 38724 21532 39116 21588
rect 39172 21532 39508 21588
rect 42354 21532 42364 21588
rect 42420 21532 43484 21588
rect 43540 21532 43550 21588
rect 6962 21420 6972 21476
rect 7028 21420 7308 21476
rect 7364 21420 18508 21476
rect 18564 21420 18574 21476
rect 20486 21420 20524 21476
rect 20580 21420 20590 21476
rect 2930 21308 2940 21364
rect 2996 21308 5292 21364
rect 5348 21308 5358 21364
rect 14802 21308 14812 21364
rect 14868 21308 22876 21364
rect 22932 21308 22942 21364
rect 14466 21196 14476 21252
rect 14532 21196 18284 21252
rect 18340 21196 18350 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 26572 21140 26628 21532
rect 28354 21420 28364 21476
rect 28420 21420 29820 21476
rect 29876 21420 29886 21476
rect 36866 21420 36876 21476
rect 36932 21420 39340 21476
rect 39396 21420 39406 21476
rect 28242 21308 28252 21364
rect 28308 21308 28700 21364
rect 28756 21308 28766 21364
rect 29698 21308 29708 21364
rect 29764 21308 30828 21364
rect 30884 21308 30894 21364
rect 31714 21308 31724 21364
rect 31780 21308 32172 21364
rect 32228 21308 32238 21364
rect 35634 21308 35644 21364
rect 35700 21308 37212 21364
rect 37268 21308 39228 21364
rect 39284 21308 39294 21364
rect 38770 21196 38780 21252
rect 38836 21196 39676 21252
rect 39732 21196 39742 21252
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 13570 21084 13580 21140
rect 13636 21084 15148 21140
rect 15204 21084 15214 21140
rect 26562 21084 26572 21140
rect 26628 21084 28252 21140
rect 28308 21084 28318 21140
rect 25890 20972 25900 21028
rect 25956 20972 26236 21028
rect 26292 20972 26302 21028
rect 30146 20972 30156 21028
rect 30212 20972 30940 21028
rect 30996 20972 31006 21028
rect 32246 20972 32284 21028
rect 32340 20972 32350 21028
rect 32806 20972 32844 21028
rect 32900 20972 32910 21028
rect 33282 20972 33292 21028
rect 33348 20972 34188 21028
rect 34244 20972 34254 21028
rect 8978 20860 8988 20916
rect 9044 20860 9996 20916
rect 10052 20860 10062 20916
rect 18162 20860 18172 20916
rect 18228 20860 19516 20916
rect 19572 20860 19582 20916
rect 29250 20860 29260 20916
rect 29316 20860 31948 20916
rect 32004 20860 33516 20916
rect 33572 20860 33582 20916
rect 43138 20860 43148 20916
rect 43204 20860 43596 20916
rect 43652 20860 44044 20916
rect 44100 20860 44110 20916
rect 8194 20748 8204 20804
rect 8260 20748 12124 20804
rect 12180 20748 12190 20804
rect 12674 20748 12684 20804
rect 12740 20748 13804 20804
rect 13860 20748 14812 20804
rect 14868 20748 14878 20804
rect 18386 20748 18396 20804
rect 18452 20748 24780 20804
rect 24836 20748 24846 20804
rect 26450 20748 26460 20804
rect 26516 20748 27244 20804
rect 27300 20748 27310 20804
rect 30940 20692 30996 20860
rect 32386 20748 32396 20804
rect 32452 20748 33404 20804
rect 33460 20748 33470 20804
rect 33730 20748 33740 20804
rect 33796 20748 34636 20804
rect 34692 20748 34702 20804
rect 34962 20748 34972 20804
rect 35028 20748 38668 20804
rect 8530 20636 8540 20692
rect 8596 20636 9660 20692
rect 9716 20636 14140 20692
rect 14196 20636 14206 20692
rect 25554 20636 25564 20692
rect 25620 20636 28028 20692
rect 28084 20636 28094 20692
rect 30930 20636 30940 20692
rect 30996 20636 31006 20692
rect 31266 20636 31276 20692
rect 31332 20636 31500 20692
rect 31556 20636 31566 20692
rect 31826 20636 31836 20692
rect 31892 20636 32284 20692
rect 32340 20636 32350 20692
rect 32610 20636 32620 20692
rect 32676 20636 38444 20692
rect 38500 20636 38510 20692
rect 38612 20580 38668 20748
rect 7522 20524 7532 20580
rect 7588 20524 8428 20580
rect 8484 20524 10556 20580
rect 10612 20524 10622 20580
rect 17042 20524 17052 20580
rect 17108 20524 18396 20580
rect 18452 20524 18462 20580
rect 21746 20524 21756 20580
rect 21812 20524 22764 20580
rect 22820 20524 22830 20580
rect 22978 20524 22988 20580
rect 23044 20524 23660 20580
rect 23716 20524 23726 20580
rect 26562 20524 26572 20580
rect 26628 20524 26908 20580
rect 26964 20524 26974 20580
rect 30594 20524 30604 20580
rect 30660 20524 32844 20580
rect 32900 20524 32910 20580
rect 34514 20524 34524 20580
rect 34580 20524 37996 20580
rect 38052 20524 38062 20580
rect 38612 20524 39676 20580
rect 39732 20524 39742 20580
rect 23426 20412 23436 20468
rect 23492 20412 38668 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 38612 20356 38668 20412
rect 21522 20300 21532 20356
rect 21588 20300 22428 20356
rect 22484 20300 26124 20356
rect 26180 20300 27804 20356
rect 27860 20300 27870 20356
rect 31164 20300 31724 20356
rect 31780 20300 31790 20356
rect 38612 20300 42476 20356
rect 42532 20300 42542 20356
rect 31164 20244 31220 20300
rect 10882 20188 10892 20244
rect 10948 20188 14364 20244
rect 14420 20188 14430 20244
rect 18050 20188 18060 20244
rect 18116 20188 20412 20244
rect 20468 20188 20478 20244
rect 26674 20188 26684 20244
rect 26740 20188 31164 20244
rect 31220 20188 31230 20244
rect 33842 20188 33852 20244
rect 33908 20188 34916 20244
rect 42578 20188 42588 20244
rect 42644 20188 43484 20244
rect 43540 20188 43550 20244
rect 18060 20132 18116 20188
rect 34860 20132 34916 20188
rect 5058 20076 5068 20132
rect 5124 20076 5852 20132
rect 5908 20076 5918 20132
rect 6962 20076 6972 20132
rect 7028 20076 8988 20132
rect 9044 20076 11340 20132
rect 11396 20076 11406 20132
rect 12786 20076 12796 20132
rect 12852 20076 13356 20132
rect 13412 20076 15148 20132
rect 15204 20076 18116 20132
rect 23874 20076 23884 20132
rect 23940 20076 25116 20132
rect 25172 20076 25182 20132
rect 25330 20076 25340 20132
rect 25396 20076 26236 20132
rect 26292 20076 28028 20132
rect 28084 20076 28094 20132
rect 29362 20076 29372 20132
rect 29428 20076 29932 20132
rect 29988 20076 32172 20132
rect 32228 20076 32238 20132
rect 32386 20076 32396 20132
rect 32452 20076 32844 20132
rect 32900 20076 33516 20132
rect 33572 20076 33582 20132
rect 34850 20076 34860 20132
rect 34916 20076 34926 20132
rect 38658 20076 38668 20132
rect 38724 20076 39004 20132
rect 39060 20076 39070 20132
rect 5618 19964 5628 20020
rect 5684 19964 6524 20020
rect 6580 19964 6590 20020
rect 10434 19964 10444 20020
rect 10500 19964 11564 20020
rect 11620 19964 14700 20020
rect 14756 19964 16380 20020
rect 16436 19964 16446 20020
rect 22642 19964 22652 20020
rect 22708 19964 23436 20020
rect 23492 19964 23502 20020
rect 26898 19964 26908 20020
rect 26964 19964 27468 20020
rect 27524 19964 27534 20020
rect 27682 19964 27692 20020
rect 27748 19964 28252 20020
rect 28308 19964 28812 20020
rect 28868 19964 28878 20020
rect 29026 19964 29036 20020
rect 29092 19964 29484 20020
rect 29540 19964 30268 20020
rect 30324 19964 30334 20020
rect 33842 19964 33852 20020
rect 33908 19964 34076 20020
rect 34132 19964 34142 20020
rect 34374 19964 34412 20020
rect 34468 19964 34478 20020
rect 38098 19964 38108 20020
rect 38164 19964 38892 20020
rect 38948 19964 38958 20020
rect 43138 19964 43148 20020
rect 43204 19964 46060 20020
rect 46116 19964 46126 20020
rect 20962 19852 20972 19908
rect 21028 19852 21980 19908
rect 22036 19852 22046 19908
rect 25890 19852 25900 19908
rect 25956 19852 27132 19908
rect 27188 19852 27198 19908
rect 27570 19852 27580 19908
rect 27636 19852 29260 19908
rect 29316 19852 29326 19908
rect 30716 19852 33068 19908
rect 33124 19852 34188 19908
rect 34244 19852 34254 19908
rect 30716 19796 30772 19852
rect 24546 19740 24556 19796
rect 24612 19740 30772 19796
rect 31154 19740 31164 19796
rect 31220 19740 36204 19796
rect 36260 19740 39452 19796
rect 39508 19740 42364 19796
rect 42420 19740 42430 19796
rect 15810 19628 15820 19684
rect 15876 19628 26796 19684
rect 26852 19628 27692 19684
rect 27748 19628 27758 19684
rect 32806 19628 32844 19684
rect 32900 19628 32910 19684
rect 36530 19628 36540 19684
rect 36596 19628 37996 19684
rect 38052 19628 38062 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 4386 19404 4396 19460
rect 4452 19404 6972 19460
rect 7028 19404 7038 19460
rect 17042 19404 17052 19460
rect 17108 19404 28924 19460
rect 28980 19404 29596 19460
rect 29652 19404 29662 19460
rect 8418 19292 8428 19348
rect 8484 19292 9884 19348
rect 9940 19292 10556 19348
rect 10612 19292 10622 19348
rect 16818 19292 16828 19348
rect 16884 19292 17276 19348
rect 17332 19292 18284 19348
rect 18340 19292 18350 19348
rect 28578 19292 28588 19348
rect 28644 19292 29372 19348
rect 29428 19292 29438 19348
rect 41794 19292 41804 19348
rect 41860 19292 45052 19348
rect 45108 19292 45118 19348
rect 26338 19180 26348 19236
rect 26404 19180 30828 19236
rect 30884 19180 30894 19236
rect 36418 19180 36428 19236
rect 36484 19180 37548 19236
rect 37604 19180 38332 19236
rect 38388 19180 38398 19236
rect 38546 19180 38556 19236
rect 38612 19180 40348 19236
rect 40404 19180 42924 19236
rect 42980 19180 43596 19236
rect 43652 19180 43662 19236
rect 14354 19068 14364 19124
rect 14420 19068 17836 19124
rect 17892 19068 19964 19124
rect 20020 19068 21868 19124
rect 21924 19068 21934 19124
rect 25554 19068 25564 19124
rect 25620 19068 27356 19124
rect 27412 19068 27422 19124
rect 27654 19068 27692 19124
rect 27748 19068 27758 19124
rect 31938 19068 31948 19124
rect 32004 19068 32284 19124
rect 32340 19068 32350 19124
rect 33058 19068 33068 19124
rect 33124 19068 38444 19124
rect 38500 19068 38510 19124
rect 44034 19068 44044 19124
rect 44100 19068 45836 19124
rect 45892 19068 45902 19124
rect 4162 18956 4172 19012
rect 4228 18956 4732 19012
rect 4788 18956 5180 19012
rect 5236 18956 9212 19012
rect 9268 18956 9278 19012
rect 9436 18956 9996 19012
rect 10052 18956 13468 19012
rect 13524 18956 13916 19012
rect 13972 18956 13982 19012
rect 35298 18956 35308 19012
rect 35364 18956 35756 19012
rect 35812 18956 41020 19012
rect 41076 18956 41086 19012
rect 9436 18900 9492 18956
rect 8866 18844 8876 18900
rect 8932 18844 9492 18900
rect 26674 18844 26684 18900
rect 26740 18844 27020 18900
rect 27076 18844 27086 18900
rect 28242 18844 28252 18900
rect 28308 18844 34972 18900
rect 35028 18844 35420 18900
rect 35476 18844 35868 18900
rect 35924 18844 35934 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 28354 18732 28364 18788
rect 28420 18732 28700 18788
rect 28756 18732 28766 18788
rect 29586 18732 29596 18788
rect 29652 18732 37660 18788
rect 37716 18732 37726 18788
rect 37996 18732 41076 18788
rect 24434 18620 24444 18676
rect 24500 18620 25564 18676
rect 25620 18620 25630 18676
rect 27122 18620 27132 18676
rect 27188 18620 27692 18676
rect 27748 18620 27758 18676
rect 32498 18620 32508 18676
rect 32564 18620 33068 18676
rect 33124 18620 33134 18676
rect 37996 18564 38052 18732
rect 38434 18620 38444 18676
rect 38500 18620 38892 18676
rect 38948 18620 38958 18676
rect 41020 18564 41076 18732
rect 43026 18620 43036 18676
rect 43092 18620 46060 18676
rect 46116 18620 46126 18676
rect 15092 18508 25004 18564
rect 25060 18508 25070 18564
rect 29026 18508 29036 18564
rect 29092 18508 30940 18564
rect 30996 18508 31006 18564
rect 35970 18508 35980 18564
rect 36036 18508 37212 18564
rect 37268 18508 38052 18564
rect 39004 18508 39508 18564
rect 41010 18508 41020 18564
rect 41076 18508 41086 18564
rect 15092 18452 15148 18508
rect 39004 18452 39060 18508
rect 39452 18452 39508 18508
rect 2594 18396 2604 18452
rect 2660 18396 4060 18452
rect 4116 18396 4126 18452
rect 9314 18396 9324 18452
rect 9380 18396 10892 18452
rect 10948 18396 10958 18452
rect 11330 18396 11340 18452
rect 11396 18396 12124 18452
rect 12180 18396 12190 18452
rect 12338 18396 12348 18452
rect 12404 18396 14252 18452
rect 14308 18396 14318 18452
rect 14690 18396 14700 18452
rect 14756 18396 15148 18452
rect 15698 18396 15708 18452
rect 15764 18396 17052 18452
rect 17108 18396 17118 18452
rect 19618 18396 19628 18452
rect 19684 18396 21756 18452
rect 21812 18396 25228 18452
rect 25284 18396 25676 18452
rect 25732 18396 25742 18452
rect 26450 18396 26460 18452
rect 26516 18396 29484 18452
rect 29540 18396 29550 18452
rect 31938 18396 31948 18452
rect 32004 18396 33964 18452
rect 34020 18396 34030 18452
rect 36642 18396 36652 18452
rect 36708 18396 36988 18452
rect 37044 18396 37772 18452
rect 37828 18396 39060 18452
rect 39218 18396 39228 18452
rect 39284 18396 39294 18452
rect 39452 18396 39676 18452
rect 39732 18396 40908 18452
rect 40964 18396 40974 18452
rect 44930 18396 44940 18452
rect 44996 18396 45836 18452
rect 45892 18396 45902 18452
rect 15708 18340 15764 18396
rect 9650 18284 9660 18340
rect 9716 18284 10108 18340
rect 10164 18284 11564 18340
rect 11620 18284 11630 18340
rect 13794 18284 13804 18340
rect 13860 18284 15764 18340
rect 24770 18284 24780 18340
rect 24836 18284 28252 18340
rect 28308 18284 28318 18340
rect 36418 18284 36428 18340
rect 36484 18284 37996 18340
rect 38052 18284 38062 18340
rect 39228 18228 39284 18396
rect 40786 18284 40796 18340
rect 40852 18284 41468 18340
rect 41524 18284 41916 18340
rect 41972 18284 41982 18340
rect 44146 18284 44156 18340
rect 44212 18284 46620 18340
rect 46676 18284 47740 18340
rect 47796 18284 48300 18340
rect 48356 18284 48366 18340
rect 10770 18172 10780 18228
rect 10836 18172 14028 18228
rect 14084 18172 14094 18228
rect 24434 18172 24444 18228
rect 24500 18172 29372 18228
rect 29428 18172 31052 18228
rect 31108 18172 31118 18228
rect 38322 18172 38332 18228
rect 38388 18172 39284 18228
rect 9762 18060 9772 18116
rect 9828 18060 10444 18116
rect 10500 18060 11228 18116
rect 11284 18060 11294 18116
rect 12002 18060 12012 18116
rect 12068 18060 13020 18116
rect 13076 18060 16156 18116
rect 16212 18060 16222 18116
rect 18386 18060 18396 18116
rect 18452 18060 20860 18116
rect 20916 18060 24780 18116
rect 24836 18060 24846 18116
rect 26758 18060 26796 18116
rect 26852 18060 26862 18116
rect 37090 18060 37100 18116
rect 37156 18060 39004 18116
rect 39060 18060 39070 18116
rect 41906 18060 41916 18116
rect 41972 18060 42812 18116
rect 42868 18060 42878 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 13794 17948 13804 18004
rect 13860 17948 14700 18004
rect 14756 17948 14766 18004
rect 16594 17948 16604 18004
rect 16660 17948 22092 18004
rect 22148 17948 22158 18004
rect 23762 17948 23772 18004
rect 23828 17948 24556 18004
rect 24612 17948 34916 18004
rect 36418 17948 36428 18004
rect 36484 17948 37436 18004
rect 37492 17948 38668 18004
rect 38724 17948 40012 18004
rect 40068 17948 40078 18004
rect 34860 17892 34916 17948
rect 11106 17836 11116 17892
rect 11172 17836 11788 17892
rect 11844 17836 15820 17892
rect 15876 17836 15886 17892
rect 16034 17836 16044 17892
rect 16100 17836 16716 17892
rect 16772 17836 18956 17892
rect 19012 17836 22988 17892
rect 23044 17836 23054 17892
rect 26982 17836 27020 17892
rect 27076 17836 27086 17892
rect 28802 17836 28812 17892
rect 28868 17836 29820 17892
rect 29876 17836 29886 17892
rect 31602 17836 31612 17892
rect 31668 17836 32732 17892
rect 32788 17836 32798 17892
rect 34850 17836 34860 17892
rect 34916 17836 35084 17892
rect 35140 17836 35420 17892
rect 35476 17836 35486 17892
rect 44034 17836 44044 17892
rect 44100 17836 44548 17892
rect 44706 17836 44716 17892
rect 44772 17836 45724 17892
rect 45780 17836 45790 17892
rect 44492 17780 44548 17836
rect 12450 17724 12460 17780
rect 12516 17724 13580 17780
rect 13636 17724 13646 17780
rect 14242 17724 14252 17780
rect 14308 17724 16604 17780
rect 16660 17724 16670 17780
rect 17042 17724 17052 17780
rect 17108 17724 19180 17780
rect 19236 17724 21588 17780
rect 27234 17724 27244 17780
rect 27300 17724 27468 17780
rect 27524 17724 27534 17780
rect 34514 17724 34524 17780
rect 34580 17724 34748 17780
rect 34804 17724 34814 17780
rect 35970 17724 35980 17780
rect 36036 17724 37212 17780
rect 37268 17724 37278 17780
rect 43810 17724 43820 17780
rect 43876 17724 44268 17780
rect 44324 17724 44334 17780
rect 44492 17724 45052 17780
rect 45108 17724 46284 17780
rect 46340 17724 46350 17780
rect 21532 17668 21588 17724
rect 4946 17612 4956 17668
rect 5012 17612 6524 17668
rect 6580 17612 8764 17668
rect 8820 17612 8830 17668
rect 9874 17612 9884 17668
rect 9940 17612 11340 17668
rect 11396 17612 11406 17668
rect 11666 17612 11676 17668
rect 11732 17612 11742 17668
rect 14802 17612 14812 17668
rect 14868 17612 16156 17668
rect 16212 17612 17388 17668
rect 17444 17612 17454 17668
rect 18274 17612 18284 17668
rect 18340 17612 19292 17668
rect 19348 17612 19358 17668
rect 21522 17612 21532 17668
rect 21588 17612 24108 17668
rect 24164 17612 24174 17668
rect 24658 17612 24668 17668
rect 24724 17612 29316 17668
rect 29474 17612 29484 17668
rect 29540 17612 37436 17668
rect 37492 17612 37502 17668
rect 38098 17612 38108 17668
rect 38164 17612 38556 17668
rect 38612 17612 39004 17668
rect 39060 17612 39070 17668
rect 39330 17612 39340 17668
rect 39396 17612 41132 17668
rect 41188 17612 41916 17668
rect 41972 17612 41982 17668
rect 11676 17556 11732 17612
rect 29260 17556 29316 17612
rect 2482 17500 2492 17556
rect 2548 17500 3836 17556
rect 3892 17500 3902 17556
rect 4610 17500 4620 17556
rect 4676 17500 6076 17556
rect 6132 17500 6748 17556
rect 6804 17500 6814 17556
rect 11106 17500 11116 17556
rect 11172 17500 11732 17556
rect 12450 17500 12460 17556
rect 12516 17500 13804 17556
rect 13860 17500 13870 17556
rect 21858 17500 21868 17556
rect 21924 17500 22092 17556
rect 22148 17500 22158 17556
rect 26786 17500 26796 17556
rect 26852 17500 27692 17556
rect 27748 17500 27758 17556
rect 29260 17500 35308 17556
rect 35746 17500 35756 17556
rect 35812 17500 36988 17556
rect 37044 17500 37054 17556
rect 35252 17444 35308 17500
rect 7858 17388 7868 17444
rect 7924 17388 13468 17444
rect 13524 17388 13534 17444
rect 15474 17388 15484 17444
rect 15540 17388 16156 17444
rect 16212 17388 20076 17444
rect 20132 17388 20142 17444
rect 26450 17388 26460 17444
rect 26516 17388 27020 17444
rect 27076 17388 27468 17444
rect 27524 17388 27534 17444
rect 30034 17388 30044 17444
rect 30100 17388 30940 17444
rect 30996 17388 31006 17444
rect 31154 17388 31164 17444
rect 31220 17388 31724 17444
rect 31780 17388 31790 17444
rect 35252 17388 36764 17444
rect 36820 17388 36830 17444
rect 10098 17276 10108 17332
rect 10164 17276 10948 17332
rect 17490 17276 17500 17332
rect 17556 17276 18732 17332
rect 18788 17276 19628 17332
rect 19684 17276 19694 17332
rect 26674 17276 26684 17332
rect 26740 17276 29932 17332
rect 29988 17276 33068 17332
rect 33124 17276 33134 17332
rect 33506 17276 33516 17332
rect 33572 17276 36708 17332
rect 39218 17276 39228 17332
rect 39284 17276 40012 17332
rect 40068 17276 41020 17332
rect 41076 17276 42364 17332
rect 42420 17276 42430 17332
rect 10892 17220 10948 17276
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 36652 17220 36708 17276
rect 10882 17164 10892 17220
rect 10948 17164 12012 17220
rect 12068 17164 13468 17220
rect 13524 17164 14588 17220
rect 14644 17164 14654 17220
rect 17602 17164 17612 17220
rect 17668 17164 19348 17220
rect 22530 17164 22540 17220
rect 22596 17164 34636 17220
rect 34692 17164 35980 17220
rect 36036 17164 36046 17220
rect 36642 17164 36652 17220
rect 36708 17164 36718 17220
rect 37426 17164 37436 17220
rect 37492 17164 41356 17220
rect 41412 17164 41422 17220
rect 19292 17108 19348 17164
rect 15362 17052 15372 17108
rect 15428 17052 16772 17108
rect 18274 17052 18284 17108
rect 18340 17052 19068 17108
rect 19124 17052 19134 17108
rect 19292 17052 19852 17108
rect 19908 17052 26908 17108
rect 27010 17052 27020 17108
rect 27076 17052 29932 17108
rect 29988 17052 32172 17108
rect 32228 17052 34076 17108
rect 34132 17052 34142 17108
rect 37650 17052 37660 17108
rect 37716 17052 38220 17108
rect 38276 17052 40908 17108
rect 40964 17052 40974 17108
rect 16716 16996 16772 17052
rect 26852 16996 26908 17052
rect 4162 16940 4172 16996
rect 4228 16940 7084 16996
rect 7140 16940 8988 16996
rect 9044 16940 10332 16996
rect 10388 16940 10398 16996
rect 11890 16940 11900 16996
rect 11956 16940 12684 16996
rect 12740 16940 12750 16996
rect 14578 16940 14588 16996
rect 14644 16940 16044 16996
rect 16100 16940 16110 16996
rect 16706 16940 16716 16996
rect 16772 16940 18060 16996
rect 18116 16940 18126 16996
rect 21298 16940 21308 16996
rect 21364 16940 21980 16996
rect 22036 16940 23772 16996
rect 23828 16940 25228 16996
rect 25284 16940 25294 16996
rect 26852 16940 33516 16996
rect 33572 16940 33582 16996
rect 33730 16940 33740 16996
rect 33796 16940 34300 16996
rect 34356 16940 34748 16996
rect 34804 16940 34814 16996
rect 35970 16940 35980 16996
rect 36036 16940 36876 16996
rect 36932 16940 36942 16996
rect 37090 16940 37100 16996
rect 37156 16940 39228 16996
rect 39284 16940 39294 16996
rect 39442 16940 39452 16996
rect 39508 16940 40572 16996
rect 40628 16940 40638 16996
rect 4946 16828 4956 16884
rect 5012 16828 9324 16884
rect 9380 16828 9390 16884
rect 9874 16828 9884 16884
rect 9940 16828 10444 16884
rect 10500 16828 10510 16884
rect 16594 16828 16604 16884
rect 16660 16828 17836 16884
rect 17892 16828 17902 16884
rect 18274 16828 18284 16884
rect 18340 16828 19068 16884
rect 19124 16828 19134 16884
rect 20636 16828 21756 16884
rect 21812 16828 22428 16884
rect 22484 16828 24668 16884
rect 24724 16828 24734 16884
rect 27318 16828 27356 16884
rect 27412 16828 27422 16884
rect 28018 16828 28028 16884
rect 28084 16828 28700 16884
rect 28756 16828 28766 16884
rect 36754 16828 36764 16884
rect 36820 16828 37884 16884
rect 37940 16828 37950 16884
rect 38612 16828 39340 16884
rect 39396 16828 39406 16884
rect 43586 16828 43596 16884
rect 43652 16828 45724 16884
rect 45780 16828 46732 16884
rect 46788 16828 46798 16884
rect 8866 16716 8876 16772
rect 8932 16716 9660 16772
rect 9716 16716 9726 16772
rect 19282 16716 19292 16772
rect 19348 16716 20076 16772
rect 20132 16716 20142 16772
rect 20636 16660 20692 16828
rect 38612 16772 38668 16828
rect 20850 16716 20860 16772
rect 20916 16716 21644 16772
rect 21700 16716 21710 16772
rect 22194 16716 22204 16772
rect 22260 16716 22876 16772
rect 22932 16716 25676 16772
rect 25732 16716 25742 16772
rect 27206 16716 27244 16772
rect 27300 16716 27310 16772
rect 30930 16716 30940 16772
rect 30996 16716 31276 16772
rect 31332 16716 31342 16772
rect 34850 16716 34860 16772
rect 34916 16716 35756 16772
rect 35812 16716 36204 16772
rect 36260 16716 36652 16772
rect 36708 16716 36718 16772
rect 36866 16716 36876 16772
rect 36932 16716 37828 16772
rect 38434 16716 38444 16772
rect 38500 16716 38668 16772
rect 41570 16716 41580 16772
rect 41636 16716 44716 16772
rect 44772 16716 44782 16772
rect 47282 16716 47292 16772
rect 47348 16716 47740 16772
rect 47796 16716 47806 16772
rect 8754 16604 8764 16660
rect 8820 16604 12124 16660
rect 12180 16604 12190 16660
rect 16146 16604 16156 16660
rect 16212 16604 18508 16660
rect 18564 16604 18574 16660
rect 20626 16604 20636 16660
rect 20692 16604 20702 16660
rect 22978 16604 22988 16660
rect 23044 16604 23996 16660
rect 24052 16604 24062 16660
rect 29922 16604 29932 16660
rect 29988 16604 30492 16660
rect 30548 16604 30558 16660
rect 32162 16604 32172 16660
rect 32228 16604 33516 16660
rect 33572 16604 35532 16660
rect 35588 16604 35598 16660
rect 36642 16604 36652 16660
rect 36708 16604 37324 16660
rect 37380 16604 37390 16660
rect 37772 16548 37828 16716
rect 38210 16604 38220 16660
rect 38276 16604 39788 16660
rect 39844 16604 39854 16660
rect 43138 16604 43148 16660
rect 43204 16604 44604 16660
rect 44660 16604 44670 16660
rect 17602 16492 17612 16548
rect 17668 16492 21476 16548
rect 37772 16492 38780 16548
rect 38836 16492 38846 16548
rect 39330 16492 39340 16548
rect 39396 16492 39900 16548
rect 39956 16492 39966 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 21420 16436 21476 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 16706 16380 16716 16436
rect 16772 16380 18620 16436
rect 18676 16380 19516 16436
rect 19572 16380 19582 16436
rect 21410 16380 21420 16436
rect 21476 16380 22428 16436
rect 22484 16380 22494 16436
rect 23874 16380 23884 16436
rect 23940 16380 32788 16436
rect 37090 16380 37100 16436
rect 37156 16380 37166 16436
rect 32732 16324 32788 16380
rect 37100 16324 37156 16380
rect 17714 16268 17724 16324
rect 17780 16268 31108 16324
rect 32732 16268 37156 16324
rect 16258 16156 16268 16212
rect 16324 16156 22988 16212
rect 23044 16156 23054 16212
rect 27906 16156 27916 16212
rect 27972 16156 28364 16212
rect 28420 16156 28924 16212
rect 28980 16156 28990 16212
rect 31052 16100 31108 16268
rect 41346 16156 41356 16212
rect 41412 16156 41692 16212
rect 41748 16156 41758 16212
rect 46050 16156 46060 16212
rect 46116 16156 48300 16212
rect 48356 16156 48366 16212
rect 7074 16044 7084 16100
rect 7140 16044 8540 16100
rect 8596 16044 8606 16100
rect 9650 16044 9660 16100
rect 9716 16044 10780 16100
rect 10836 16044 10846 16100
rect 15362 16044 15372 16100
rect 15428 16044 17612 16100
rect 17668 16044 17678 16100
rect 20402 16044 20412 16100
rect 20468 16044 21756 16100
rect 21812 16044 21822 16100
rect 28242 16044 28252 16100
rect 28308 16044 29484 16100
rect 29540 16044 29550 16100
rect 31052 16044 36316 16100
rect 36372 16044 36382 16100
rect 17938 15932 17948 15988
rect 18004 15932 18956 15988
rect 19012 15932 19022 15988
rect 19618 15932 19628 15988
rect 19684 15932 23548 15988
rect 23604 15932 23614 15988
rect 31154 15932 31164 15988
rect 31220 15932 34300 15988
rect 34356 15932 34366 15988
rect 36054 15932 36092 15988
rect 36148 15932 36158 15988
rect 36978 15932 36988 15988
rect 37044 15932 37082 15988
rect 42690 15932 42700 15988
rect 42756 15932 43820 15988
rect 43876 15932 44828 15988
rect 44884 15932 45500 15988
rect 45556 15932 45566 15988
rect 2482 15820 2492 15876
rect 2548 15820 3836 15876
rect 3892 15820 3902 15876
rect 9426 15820 9436 15876
rect 9492 15820 10556 15876
rect 10612 15820 11564 15876
rect 11620 15820 11630 15876
rect 20178 15820 20188 15876
rect 20244 15820 21980 15876
rect 22036 15820 22046 15876
rect 26982 15820 27020 15876
rect 27076 15820 27086 15876
rect 33170 15820 33180 15876
rect 33236 15820 36540 15876
rect 36596 15820 36606 15876
rect 44594 15820 44604 15876
rect 44660 15820 45052 15876
rect 45108 15820 45118 15876
rect 15810 15708 15820 15764
rect 15876 15708 15886 15764
rect 30930 15708 30940 15764
rect 30996 15708 37100 15764
rect 37156 15708 38556 15764
rect 38612 15708 38622 15764
rect 15820 15540 15876 15708
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 27122 15596 27132 15652
rect 27188 15596 29932 15652
rect 29988 15596 29998 15652
rect 31266 15596 31276 15652
rect 31332 15596 32284 15652
rect 32340 15596 32350 15652
rect 32610 15596 32620 15652
rect 32676 15596 33180 15652
rect 33236 15596 33246 15652
rect 35410 15596 35420 15652
rect 35476 15596 41468 15652
rect 41524 15596 41534 15652
rect 15250 15484 15260 15540
rect 15316 15484 15596 15540
rect 15652 15484 16492 15540
rect 16548 15484 16558 15540
rect 19506 15484 19516 15540
rect 19572 15484 21196 15540
rect 21252 15484 21262 15540
rect 22194 15484 22204 15540
rect 22260 15484 22270 15540
rect 28578 15484 28588 15540
rect 28644 15484 37548 15540
rect 37604 15484 37614 15540
rect 37986 15484 37996 15540
rect 38052 15484 38780 15540
rect 38836 15484 38846 15540
rect 46610 15484 46620 15540
rect 46676 15484 47292 15540
rect 47348 15484 47358 15540
rect 22204 15428 22260 15484
rect 37996 15428 38052 15484
rect 8418 15372 8428 15428
rect 8484 15372 9660 15428
rect 9716 15372 9726 15428
rect 12786 15372 12796 15428
rect 12852 15372 21420 15428
rect 21476 15372 22260 15428
rect 25862 15372 25900 15428
rect 25956 15372 25966 15428
rect 37174 15372 37212 15428
rect 37268 15372 37278 15428
rect 37426 15372 37436 15428
rect 37492 15372 38052 15428
rect 11666 15260 11676 15316
rect 11732 15260 14364 15316
rect 14420 15260 14924 15316
rect 14980 15260 14990 15316
rect 21970 15260 21980 15316
rect 22036 15260 22316 15316
rect 22372 15260 22382 15316
rect 23538 15260 23548 15316
rect 23604 15260 24556 15316
rect 24612 15260 27244 15316
rect 27300 15260 27310 15316
rect 31938 15260 31948 15316
rect 32004 15260 32284 15316
rect 32340 15260 33404 15316
rect 33460 15260 33470 15316
rect 34626 15260 34636 15316
rect 34692 15260 35644 15316
rect 35700 15260 35710 15316
rect 36642 15260 36652 15316
rect 36708 15260 36718 15316
rect 37538 15260 37548 15316
rect 37604 15260 37884 15316
rect 37940 15260 37950 15316
rect 36652 15204 36708 15260
rect 16034 15148 16044 15204
rect 16100 15148 19740 15204
rect 19796 15148 19806 15204
rect 20962 15148 20972 15204
rect 21028 15148 21532 15204
rect 21588 15148 22204 15204
rect 22260 15148 22270 15204
rect 24658 15148 24668 15204
rect 24724 15148 25452 15204
rect 25508 15148 25518 15204
rect 27570 15148 27580 15204
rect 27636 15148 28252 15204
rect 28308 15148 28318 15204
rect 34066 15148 34076 15204
rect 34132 15148 36708 15204
rect 37426 15148 37436 15204
rect 37492 15148 38332 15204
rect 38388 15148 38892 15204
rect 38948 15148 38958 15204
rect 4610 15036 4620 15092
rect 4676 15036 5740 15092
rect 5796 15036 5806 15092
rect 6066 15036 6076 15092
rect 6132 15036 7756 15092
rect 7812 15036 10108 15092
rect 10164 15036 11564 15092
rect 11620 15036 11630 15092
rect 13122 15036 13132 15092
rect 13188 15036 44268 15092
rect 44324 15036 44334 15092
rect 17154 14924 17164 14980
rect 17220 14924 25340 14980
rect 25396 14924 25406 14980
rect 27906 14924 27916 14980
rect 27972 14924 30492 14980
rect 30548 14924 33964 14980
rect 34020 14924 34030 14980
rect 35634 14924 35644 14980
rect 35700 14924 36092 14980
rect 36148 14924 36158 14980
rect 37846 14924 37884 14980
rect 37940 14924 37950 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 7410 14812 7420 14868
rect 7476 14812 8204 14868
rect 8260 14812 8270 14868
rect 20066 14812 20076 14868
rect 20132 14812 25228 14868
rect 25284 14812 26124 14868
rect 26180 14812 26190 14868
rect 33730 14812 33740 14868
rect 33796 14812 34972 14868
rect 35028 14812 35038 14868
rect 36166 14812 36204 14868
rect 36260 14812 39564 14868
rect 39620 14812 39630 14868
rect 5170 14700 5180 14756
rect 5236 14700 6076 14756
rect 6132 14700 10332 14756
rect 10388 14700 10398 14756
rect 19842 14700 19852 14756
rect 19908 14700 20636 14756
rect 20692 14700 20702 14756
rect 27122 14700 27132 14756
rect 27188 14700 27692 14756
rect 27748 14700 27758 14756
rect 34850 14700 34860 14756
rect 34916 14700 36988 14756
rect 37044 14700 37054 14756
rect 8418 14588 8428 14644
rect 8484 14588 11004 14644
rect 11060 14588 12236 14644
rect 12292 14588 12302 14644
rect 14690 14588 14700 14644
rect 14756 14588 17276 14644
rect 17332 14588 17342 14644
rect 20850 14588 20860 14644
rect 20916 14588 21756 14644
rect 21812 14588 22540 14644
rect 22596 14588 22606 14644
rect 23202 14588 23212 14644
rect 23268 14588 27468 14644
rect 27524 14588 27534 14644
rect 30930 14588 30940 14644
rect 30996 14588 35644 14644
rect 35700 14588 38556 14644
rect 38612 14588 38622 14644
rect 7634 14476 7644 14532
rect 7700 14476 8540 14532
rect 8596 14476 8606 14532
rect 17154 14476 17164 14532
rect 17220 14476 17724 14532
rect 17780 14476 20300 14532
rect 20356 14476 21308 14532
rect 21364 14476 21374 14532
rect 21532 14476 23548 14532
rect 23604 14476 23614 14532
rect 31378 14476 31388 14532
rect 31444 14476 31948 14532
rect 32004 14476 32014 14532
rect 32274 14476 32284 14532
rect 32340 14476 33404 14532
rect 33460 14476 33470 14532
rect 35942 14476 35980 14532
rect 36036 14476 36046 14532
rect 21532 14420 21588 14476
rect 17042 14364 17052 14420
rect 17108 14364 17388 14420
rect 17444 14364 21588 14420
rect 22978 14364 22988 14420
rect 23044 14364 23996 14420
rect 24052 14364 25004 14420
rect 25060 14364 25070 14420
rect 31042 14364 31052 14420
rect 31108 14364 31500 14420
rect 31556 14364 31566 14420
rect 33954 14364 33964 14420
rect 34020 14364 35196 14420
rect 35252 14364 36092 14420
rect 36148 14364 36158 14420
rect 3602 14252 3612 14308
rect 3668 14252 5068 14308
rect 5124 14252 5964 14308
rect 6020 14252 6972 14308
rect 7028 14252 11116 14308
rect 11172 14252 11340 14308
rect 11396 14252 14364 14308
rect 14420 14252 14430 14308
rect 16034 14252 16044 14308
rect 16100 14252 16604 14308
rect 16660 14252 16670 14308
rect 20178 14252 20188 14308
rect 20244 14252 21084 14308
rect 21140 14252 22092 14308
rect 22148 14252 22158 14308
rect 24658 14252 24668 14308
rect 24724 14252 25564 14308
rect 25620 14252 28588 14308
rect 28644 14252 28654 14308
rect 25666 14140 25676 14196
rect 25732 14140 29708 14196
rect 29764 14140 29774 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 28354 14028 28364 14084
rect 28420 14028 30380 14084
rect 30436 14028 30940 14084
rect 30996 14028 31006 14084
rect 37174 14028 37212 14084
rect 37268 14028 37278 14084
rect 12002 13916 12012 13972
rect 12068 13916 15708 13972
rect 15764 13916 15774 13972
rect 19170 13916 19180 13972
rect 19236 13916 21308 13972
rect 21364 13916 21374 13972
rect 29810 13916 29820 13972
rect 29876 13916 34524 13972
rect 34580 13916 34972 13972
rect 35028 13916 35038 13972
rect 38434 13916 38444 13972
rect 38500 13916 40796 13972
rect 40852 13916 41132 13972
rect 41188 13916 41692 13972
rect 41748 13916 41758 13972
rect 45154 13916 45164 13972
rect 45220 13916 46508 13972
rect 46564 13916 46574 13972
rect 6290 13804 6300 13860
rect 6356 13804 7980 13860
rect 8036 13804 8046 13860
rect 15250 13804 15260 13860
rect 15316 13804 16268 13860
rect 16324 13804 16334 13860
rect 28466 13804 28476 13860
rect 28532 13804 34860 13860
rect 34916 13804 35532 13860
rect 35588 13804 35598 13860
rect 1698 13692 1708 13748
rect 1764 13692 3612 13748
rect 3668 13692 3678 13748
rect 6850 13692 6860 13748
rect 6916 13692 7756 13748
rect 7812 13692 9884 13748
rect 9940 13692 9950 13748
rect 16146 13692 16156 13748
rect 16212 13692 17612 13748
rect 17668 13692 17678 13748
rect 20738 13692 20748 13748
rect 20804 13692 21420 13748
rect 21476 13692 22988 13748
rect 23044 13692 23054 13748
rect 28578 13692 28588 13748
rect 28644 13692 29484 13748
rect 29540 13692 29550 13748
rect 30146 13692 30156 13748
rect 30212 13692 30492 13748
rect 30548 13692 30558 13748
rect 32722 13692 32732 13748
rect 32788 13692 34076 13748
rect 34132 13692 34188 13748
rect 34244 13692 34254 13748
rect 36082 13692 36092 13748
rect 36148 13692 36316 13748
rect 36372 13692 36382 13748
rect 37314 13692 37324 13748
rect 37380 13692 38220 13748
rect 38276 13692 38668 13748
rect 45826 13692 45836 13748
rect 45892 13692 47404 13748
rect 47460 13692 47740 13748
rect 47796 13692 48300 13748
rect 48356 13692 48366 13748
rect 15026 13580 15036 13636
rect 15092 13524 15148 13636
rect 15474 13580 15484 13636
rect 15540 13580 17500 13636
rect 17556 13580 17566 13636
rect 24322 13580 24332 13636
rect 24388 13580 28364 13636
rect 28420 13580 28430 13636
rect 31154 13580 31164 13636
rect 31220 13580 31612 13636
rect 31668 13580 33180 13636
rect 33236 13580 33246 13636
rect 33618 13580 33628 13636
rect 33684 13580 36540 13636
rect 36596 13580 37548 13636
rect 37604 13580 37614 13636
rect 38612 13580 38668 13692
rect 38724 13580 38734 13636
rect 4956 13468 9212 13524
rect 9268 13468 9278 13524
rect 15092 13468 15260 13524
rect 15316 13468 15708 13524
rect 15764 13468 15774 13524
rect 17826 13468 17836 13524
rect 17892 13468 19068 13524
rect 19124 13468 20188 13524
rect 20244 13468 20254 13524
rect 26450 13468 26460 13524
rect 26516 13468 27132 13524
rect 27188 13468 33292 13524
rect 33348 13468 33358 13524
rect 34972 13468 35308 13524
rect 35364 13468 35374 13524
rect 4956 13412 5012 13468
rect 4946 13356 4956 13412
rect 5012 13356 5022 13412
rect 5730 13356 5740 13412
rect 5796 13356 6748 13412
rect 6804 13356 20524 13412
rect 20580 13356 23548 13412
rect 25778 13356 25788 13412
rect 25844 13356 30604 13412
rect 30660 13356 30670 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 14242 13244 14252 13300
rect 14308 13244 16044 13300
rect 16100 13244 16110 13300
rect 23492 13188 23548 13356
rect 34972 13300 35028 13468
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 28354 13244 28364 13300
rect 28420 13244 29148 13300
rect 29204 13244 35028 13300
rect 23492 13132 23772 13188
rect 23828 13132 23838 13188
rect 27906 13132 27916 13188
rect 27972 13132 28252 13188
rect 28308 13132 28318 13188
rect 29362 13132 29372 13188
rect 29428 13132 30716 13188
rect 30772 13132 30782 13188
rect 14354 13020 14364 13076
rect 14420 13020 14812 13076
rect 14868 13020 16380 13076
rect 16436 13020 16446 13076
rect 21186 13020 21196 13076
rect 21252 13020 21644 13076
rect 21700 13020 24108 13076
rect 24164 13020 24174 13076
rect 26898 13020 26908 13076
rect 26964 13020 30660 13076
rect 33170 13020 33180 13076
rect 33236 13020 33852 13076
rect 33908 13020 33918 13076
rect 35186 13020 35196 13076
rect 35252 13020 35756 13076
rect 35812 13020 37996 13076
rect 38052 13020 38062 13076
rect 30604 12964 30660 13020
rect 4946 12908 4956 12964
rect 5012 12908 6188 12964
rect 6244 12908 6254 12964
rect 15810 12908 15820 12964
rect 15876 12908 16940 12964
rect 16996 12908 17388 12964
rect 17444 12908 17454 12964
rect 27346 12908 27356 12964
rect 27412 12908 29596 12964
rect 29652 12908 29662 12964
rect 30604 12908 30716 12964
rect 30772 12908 33516 12964
rect 33572 12908 34972 12964
rect 35028 12908 35038 12964
rect 29596 12852 29652 12908
rect 2594 12796 2604 12852
rect 2660 12796 3836 12852
rect 3892 12796 3902 12852
rect 8754 12796 8764 12852
rect 8820 12796 11228 12852
rect 11284 12796 11294 12852
rect 15922 12796 15932 12852
rect 15988 12796 16492 12852
rect 16548 12796 17836 12852
rect 17892 12796 17902 12852
rect 25442 12796 25452 12852
rect 25508 12796 29372 12852
rect 29428 12796 29438 12852
rect 29596 12796 34188 12852
rect 34244 12796 34254 12852
rect 34402 12796 34412 12852
rect 34468 12796 34860 12852
rect 34916 12796 35868 12852
rect 35924 12796 36428 12852
rect 36484 12796 37436 12852
rect 37492 12796 37502 12852
rect 37874 12796 37884 12852
rect 37940 12796 38668 12852
rect 38724 12796 38734 12852
rect 34188 12740 34244 12796
rect 8866 12684 8876 12740
rect 8932 12684 12124 12740
rect 12180 12684 12190 12740
rect 14130 12684 14140 12740
rect 14196 12684 16156 12740
rect 16212 12684 16222 12740
rect 23874 12684 23884 12740
rect 23940 12684 25004 12740
rect 25060 12684 25070 12740
rect 26114 12684 26124 12740
rect 26180 12684 26236 12740
rect 26292 12684 26302 12740
rect 27682 12684 27692 12740
rect 27748 12684 29260 12740
rect 29316 12684 29326 12740
rect 30370 12684 30380 12740
rect 30436 12684 32620 12740
rect 32676 12684 32686 12740
rect 34188 12684 34524 12740
rect 34580 12684 34590 12740
rect 41122 12684 41132 12740
rect 41188 12684 44940 12740
rect 44996 12684 45006 12740
rect 15138 12572 15148 12628
rect 15204 12572 18620 12628
rect 18676 12572 18686 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 25004 12516 25060 12684
rect 26786 12572 26796 12628
rect 26852 12572 36316 12628
rect 36372 12572 36382 12628
rect 15922 12460 15932 12516
rect 15988 12460 16492 12516
rect 16548 12460 16558 12516
rect 25004 12460 27020 12516
rect 27076 12460 28364 12516
rect 28420 12460 28430 12516
rect 29250 12460 29260 12516
rect 29316 12460 33628 12516
rect 33684 12460 33694 12516
rect 34038 12460 34076 12516
rect 34132 12460 34142 12516
rect 34374 12460 34412 12516
rect 34468 12460 34478 12516
rect 3602 12348 3612 12404
rect 3668 12348 4172 12404
rect 4228 12348 5292 12404
rect 5348 12348 7308 12404
rect 7364 12348 7374 12404
rect 15026 12348 15036 12404
rect 15092 12348 17724 12404
rect 17780 12348 17790 12404
rect 25890 12348 25900 12404
rect 25956 12348 27356 12404
rect 27412 12348 28420 12404
rect 33282 12348 33292 12404
rect 33348 12348 36092 12404
rect 36148 12348 37324 12404
rect 37380 12348 39228 12404
rect 39284 12348 39294 12404
rect 42578 12348 42588 12404
rect 42644 12348 44828 12404
rect 44884 12348 44894 12404
rect 28364 12292 28420 12348
rect 16258 12236 16268 12292
rect 16324 12236 21980 12292
rect 22036 12236 22316 12292
rect 22372 12236 22382 12292
rect 24210 12236 24220 12292
rect 24276 12236 26460 12292
rect 26516 12236 26796 12292
rect 26852 12236 26862 12292
rect 27682 12236 27692 12292
rect 27748 12236 28140 12292
rect 28196 12236 28206 12292
rect 28354 12236 28364 12292
rect 28420 12236 28430 12292
rect 31042 12236 31052 12292
rect 31108 12236 31500 12292
rect 31556 12236 32396 12292
rect 32452 12236 33068 12292
rect 33124 12236 33134 12292
rect 12338 12124 12348 12180
rect 12404 12124 23884 12180
rect 23940 12124 23950 12180
rect 27346 12124 27356 12180
rect 27412 12124 29148 12180
rect 29204 12124 29214 12180
rect 29586 12124 29596 12180
rect 29652 12124 32508 12180
rect 32564 12124 34300 12180
rect 34356 12124 34366 12180
rect 34514 12124 34524 12180
rect 34580 12124 37548 12180
rect 37604 12124 37614 12180
rect 14690 12012 14700 12068
rect 14756 12012 15596 12068
rect 15652 12012 15662 12068
rect 17938 12012 17948 12068
rect 18004 12012 18620 12068
rect 18676 12012 18686 12068
rect 22082 12012 22092 12068
rect 22148 12012 23548 12068
rect 23604 12012 23614 12068
rect 29810 12012 29820 12068
rect 29876 12012 31612 12068
rect 31668 12012 31948 12068
rect 32004 12012 32014 12068
rect 38770 12012 38780 12068
rect 38836 12012 40124 12068
rect 40180 12012 40190 12068
rect 43586 12012 43596 12068
rect 43652 12012 45276 12068
rect 45332 12012 45342 12068
rect 14354 11900 14364 11956
rect 14420 11900 14430 11956
rect 20290 11900 20300 11956
rect 20356 11900 20748 11956
rect 20804 11900 20814 11956
rect 22642 11900 22652 11956
rect 22708 11900 22718 11956
rect 34822 11900 34860 11956
rect 34916 11900 34926 11956
rect 35186 11900 35196 11956
rect 35252 11900 36092 11956
rect 36148 11900 36158 11956
rect 14130 11788 14140 11844
rect 14196 11788 14308 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 7970 11676 7980 11732
rect 8036 11676 8764 11732
rect 8820 11676 8830 11732
rect 14252 11620 14308 11788
rect 14364 11732 14420 11900
rect 22652 11732 22708 11900
rect 44370 11788 44380 11844
rect 44436 11788 46284 11844
rect 46340 11788 46956 11844
rect 47012 11788 47022 11844
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 14364 11676 16044 11732
rect 16100 11676 16110 11732
rect 21074 11676 21084 11732
rect 21140 11676 21756 11732
rect 21812 11676 23324 11732
rect 23380 11676 23390 11732
rect 27906 11676 27916 11732
rect 27972 11676 29932 11732
rect 29988 11676 29998 11732
rect 31714 11676 31724 11732
rect 31780 11676 31948 11732
rect 32004 11676 32508 11732
rect 32564 11676 32574 11732
rect 14252 11564 14756 11620
rect 15026 11564 15036 11620
rect 15092 11564 15372 11620
rect 15428 11564 15438 11620
rect 21858 11564 21868 11620
rect 21924 11564 22876 11620
rect 22932 11564 22942 11620
rect 34626 11564 34636 11620
rect 34692 11564 34972 11620
rect 35028 11564 35038 11620
rect 14700 11508 14756 11564
rect 12898 11452 12908 11508
rect 12964 11452 13916 11508
rect 13972 11452 14308 11508
rect 14690 11452 14700 11508
rect 14756 11452 14766 11508
rect 18050 11452 18060 11508
rect 18116 11452 18956 11508
rect 19012 11452 19022 11508
rect 30258 11452 30268 11508
rect 30324 11452 35420 11508
rect 35476 11452 35486 11508
rect 14252 11396 14308 11452
rect 14242 11340 14252 11396
rect 14308 11340 14318 11396
rect 17826 11340 17836 11396
rect 17892 11340 18732 11396
rect 18788 11340 19068 11396
rect 19124 11340 19134 11396
rect 27794 11340 27804 11396
rect 27860 11340 30604 11396
rect 30660 11340 30828 11396
rect 30884 11340 30894 11396
rect 37202 11340 37212 11396
rect 37268 11340 38108 11396
rect 38164 11340 38174 11396
rect 41010 11340 41020 11396
rect 41076 11340 41916 11396
rect 41972 11340 41982 11396
rect 23202 11228 23212 11284
rect 23268 11228 24332 11284
rect 24388 11228 24398 11284
rect 4946 11116 4956 11172
rect 5012 11116 7868 11172
rect 7924 11116 7934 11172
rect 18946 11116 18956 11172
rect 19012 11116 21196 11172
rect 21252 11116 21262 11172
rect 37986 11116 37996 11172
rect 38052 11116 39452 11172
rect 39508 11116 39518 11172
rect 14914 11004 14924 11060
rect 14980 11004 15260 11060
rect 15316 11004 15326 11060
rect 20962 11004 20972 11060
rect 21028 11004 22316 11060
rect 22372 11004 22382 11060
rect 23762 11004 23772 11060
rect 23828 11004 34524 11060
rect 34580 11004 34590 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 9314 10892 9324 10948
rect 9380 10892 19684 10948
rect 20178 10892 20188 10948
rect 20244 10892 20748 10948
rect 20804 10892 20814 10948
rect 34626 10892 34636 10948
rect 34692 10892 35084 10948
rect 35140 10892 39340 10948
rect 39396 10892 39406 10948
rect 19628 10836 19684 10892
rect 14130 10780 14140 10836
rect 14196 10780 14812 10836
rect 14868 10780 15260 10836
rect 15316 10780 15326 10836
rect 16146 10780 16156 10836
rect 16212 10780 18956 10836
rect 19012 10780 19022 10836
rect 19628 10780 35532 10836
rect 35588 10780 35598 10836
rect 38098 10780 38108 10836
rect 38164 10780 41132 10836
rect 41188 10780 41198 10836
rect 45266 10780 45276 10836
rect 45332 10780 45724 10836
rect 45780 10780 45790 10836
rect 37314 10668 37324 10724
rect 37380 10668 38780 10724
rect 38836 10668 38846 10724
rect 45938 10668 45948 10724
rect 46004 10668 47292 10724
rect 47348 10668 47358 10724
rect 8642 10556 8652 10612
rect 8708 10556 9660 10612
rect 9716 10556 11452 10612
rect 11508 10556 11518 10612
rect 19058 10556 19068 10612
rect 19124 10556 19516 10612
rect 19572 10556 19582 10612
rect 19730 10556 19740 10612
rect 19796 10556 21084 10612
rect 21140 10556 21150 10612
rect 29474 10556 29484 10612
rect 29540 10556 31052 10612
rect 31108 10556 31118 10612
rect 37762 10556 37772 10612
rect 37828 10556 39788 10612
rect 39844 10556 39854 10612
rect 19516 10500 19572 10556
rect 12450 10444 12460 10500
rect 12516 10444 13132 10500
rect 13188 10444 13198 10500
rect 19516 10444 21980 10500
rect 22036 10444 22876 10500
rect 22932 10444 22942 10500
rect 27794 10444 27804 10500
rect 27860 10444 28140 10500
rect 28196 10444 28206 10500
rect 38434 10444 38444 10500
rect 38500 10444 40796 10500
rect 40852 10444 42140 10500
rect 42196 10444 44940 10500
rect 44996 10444 45500 10500
rect 45556 10444 45566 10500
rect 10882 10332 10892 10388
rect 10948 10332 12908 10388
rect 12964 10332 12974 10388
rect 13570 10332 13580 10388
rect 13636 10332 15820 10388
rect 15876 10332 28476 10388
rect 28532 10332 28542 10388
rect 43474 10332 43484 10388
rect 43540 10332 46844 10388
rect 46900 10332 46910 10388
rect 13122 10220 13132 10276
rect 13188 10220 30828 10276
rect 30884 10220 30894 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 20626 10108 20636 10164
rect 20692 10108 21532 10164
rect 21588 10108 21598 10164
rect 26226 10108 26236 10164
rect 26292 10108 31892 10164
rect 31836 10052 31892 10108
rect 16258 9996 16268 10052
rect 16324 9996 18172 10052
rect 18228 9996 19180 10052
rect 19236 9996 19246 10052
rect 21298 9996 21308 10052
rect 21364 9996 21644 10052
rect 21700 9996 21710 10052
rect 26674 9996 26684 10052
rect 26740 9996 28140 10052
rect 28196 9996 28206 10052
rect 31836 9996 33068 10052
rect 33124 9996 34860 10052
rect 34916 9996 34926 10052
rect 35084 9996 35868 10052
rect 35924 9996 36988 10052
rect 37044 9996 37054 10052
rect 37202 9996 37212 10052
rect 37268 9996 37996 10052
rect 38052 9996 38062 10052
rect 35084 9940 35140 9996
rect 11442 9884 11452 9940
rect 11508 9884 12684 9940
rect 12740 9884 12750 9940
rect 18834 9884 18844 9940
rect 18900 9884 22484 9940
rect 22642 9884 22652 9940
rect 22708 9884 24892 9940
rect 24948 9884 24958 9940
rect 31042 9884 31052 9940
rect 31108 9884 31836 9940
rect 31892 9884 35140 9940
rect 35746 9884 35756 9940
rect 35812 9884 36092 9940
rect 36148 9884 39116 9940
rect 39172 9884 39182 9940
rect 46498 9884 46508 9940
rect 46564 9884 48300 9940
rect 48356 9884 48366 9940
rect 22428 9828 22484 9884
rect 12562 9772 12572 9828
rect 12628 9772 13580 9828
rect 13636 9772 13646 9828
rect 20738 9772 20748 9828
rect 20804 9772 21644 9828
rect 21700 9772 21710 9828
rect 22428 9772 24220 9828
rect 24276 9772 25788 9828
rect 25844 9772 25854 9828
rect 31378 9772 31388 9828
rect 31444 9772 33852 9828
rect 33908 9772 33918 9828
rect 35522 9772 35532 9828
rect 35588 9772 38668 9828
rect 38612 9716 38668 9772
rect 2482 9660 2492 9716
rect 2548 9660 3500 9716
rect 3556 9660 3566 9716
rect 6402 9660 6412 9716
rect 6468 9660 7644 9716
rect 7700 9660 7710 9716
rect 8194 9660 8204 9716
rect 8260 9660 8540 9716
rect 8596 9660 8606 9716
rect 17490 9660 17500 9716
rect 17556 9660 17836 9716
rect 17892 9660 19292 9716
rect 19348 9660 26908 9716
rect 26964 9660 26974 9716
rect 32050 9660 32060 9716
rect 32116 9660 32844 9716
rect 32900 9660 34076 9716
rect 34132 9660 35644 9716
rect 35700 9660 35710 9716
rect 38612 9660 39004 9716
rect 39060 9660 39070 9716
rect 40786 9660 40796 9716
rect 40852 9660 41916 9716
rect 41972 9660 41982 9716
rect 10994 9548 11004 9604
rect 11060 9548 12348 9604
rect 12404 9548 13468 9604
rect 13524 9548 13534 9604
rect 15250 9548 15260 9604
rect 15316 9548 16604 9604
rect 16660 9548 16670 9604
rect 19842 9548 19852 9604
rect 19908 9548 21308 9604
rect 21364 9548 21374 9604
rect 29474 9548 29484 9604
rect 29540 9548 30716 9604
rect 30772 9548 30782 9604
rect 32610 9548 32620 9604
rect 32676 9548 34636 9604
rect 34692 9548 37212 9604
rect 37268 9548 38108 9604
rect 38164 9548 38174 9604
rect 38108 9492 38164 9548
rect 14914 9436 14924 9492
rect 14980 9436 16044 9492
rect 16100 9436 16110 9492
rect 17612 9436 18172 9492
rect 18228 9436 18238 9492
rect 28130 9436 28140 9492
rect 28196 9436 28364 9492
rect 28420 9436 32284 9492
rect 32340 9436 34300 9492
rect 34356 9436 34366 9492
rect 38108 9436 39676 9492
rect 39732 9436 39742 9492
rect 17612 9268 17668 9436
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 18274 9324 18284 9380
rect 18340 9324 18844 9380
rect 18900 9324 18910 9380
rect 20738 9324 20748 9380
rect 20804 9324 21644 9380
rect 21700 9324 21710 9380
rect 29362 9324 29372 9380
rect 29428 9324 35532 9380
rect 35588 9324 35598 9380
rect 16258 9212 16268 9268
rect 16324 9212 16334 9268
rect 17154 9212 17164 9268
rect 17220 9212 17612 9268
rect 17668 9212 17678 9268
rect 18610 9212 18620 9268
rect 18676 9212 18686 9268
rect 19394 9212 19404 9268
rect 19460 9212 20188 9268
rect 20244 9212 21532 9268
rect 21588 9212 21598 9268
rect 30034 9212 30044 9268
rect 30100 9212 30380 9268
rect 30436 9212 30446 9268
rect 39442 9212 39452 9268
rect 39508 9212 41244 9268
rect 41300 9212 41310 9268
rect 4386 9100 4396 9156
rect 4452 9100 7084 9156
rect 7140 9100 7150 9156
rect 6626 8988 6636 9044
rect 6692 8988 7420 9044
rect 7476 8988 7486 9044
rect 8306 8988 8316 9044
rect 8372 8988 9436 9044
rect 9492 8988 9502 9044
rect 16268 8932 16324 9212
rect 18620 9156 18676 9212
rect 18620 9100 18956 9156
rect 19012 9100 19852 9156
rect 19908 9100 19918 9156
rect 21186 9100 21196 9156
rect 21252 9100 21644 9156
rect 21700 9100 21710 9156
rect 23874 9100 23884 9156
rect 23940 9100 24668 9156
rect 24724 9100 25228 9156
rect 25284 9100 25294 9156
rect 28130 9100 28140 9156
rect 28196 9100 37212 9156
rect 37268 9100 37278 9156
rect 17266 8988 17276 9044
rect 17332 8988 18396 9044
rect 18452 8988 18462 9044
rect 19170 8988 19180 9044
rect 19236 8988 22988 9044
rect 23044 8988 23054 9044
rect 26852 8988 27580 9044
rect 27636 8988 29148 9044
rect 29204 8988 29214 9044
rect 30706 8988 30716 9044
rect 30772 8988 33404 9044
rect 33460 8988 33470 9044
rect 15362 8876 15372 8932
rect 15428 8876 16324 8932
rect 16818 8876 16828 8932
rect 16884 8876 18844 8932
rect 18900 8876 18910 8932
rect 21298 8876 21308 8932
rect 21364 8876 22204 8932
rect 22260 8876 23772 8932
rect 23828 8876 24556 8932
rect 24612 8876 24622 8932
rect 26852 8820 26908 8988
rect 32274 8876 32284 8932
rect 32340 8876 33068 8932
rect 33124 8876 33134 8932
rect 37314 8876 37324 8932
rect 37380 8876 38108 8932
rect 38164 8876 38174 8932
rect 38770 8876 38780 8932
rect 38836 8876 40796 8932
rect 40852 8876 40862 8932
rect 2482 8764 2492 8820
rect 2548 8764 3388 8820
rect 3444 8764 3454 8820
rect 17938 8764 17948 8820
rect 18004 8764 18284 8820
rect 18340 8764 18350 8820
rect 18498 8764 18508 8820
rect 18564 8764 19292 8820
rect 19348 8764 19358 8820
rect 23650 8764 23660 8820
rect 23716 8764 26908 8820
rect 28466 8764 28476 8820
rect 28532 8764 29260 8820
rect 29316 8764 35420 8820
rect 35476 8764 35486 8820
rect 9650 8652 9660 8708
rect 9716 8652 25228 8708
rect 25284 8652 25294 8708
rect 36418 8652 36428 8708
rect 36484 8652 38108 8708
rect 38164 8652 38174 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 11890 8540 11900 8596
rect 11956 8540 12908 8596
rect 12964 8540 31052 8596
rect 31108 8540 31118 8596
rect 16482 8428 16492 8484
rect 16548 8428 17276 8484
rect 17332 8428 17342 8484
rect 21634 8428 21644 8484
rect 21700 8428 28140 8484
rect 28196 8428 28206 8484
rect 28466 8428 28476 8484
rect 28532 8428 30324 8484
rect 33282 8428 33292 8484
rect 33348 8428 34076 8484
rect 34132 8428 34142 8484
rect 34402 8428 34412 8484
rect 34468 8428 38668 8484
rect 30268 8372 30324 8428
rect 38612 8372 38668 8428
rect 13682 8316 13692 8372
rect 13748 8316 14812 8372
rect 14868 8316 14878 8372
rect 15474 8316 15484 8372
rect 15540 8316 16044 8372
rect 16100 8316 16380 8372
rect 16436 8316 16446 8372
rect 18722 8316 18732 8372
rect 18788 8316 25676 8372
rect 25732 8316 25742 8372
rect 25890 8316 25900 8372
rect 25956 8316 27132 8372
rect 27188 8316 27804 8372
rect 27860 8316 29708 8372
rect 29764 8316 29774 8372
rect 30268 8316 32172 8372
rect 32228 8316 32238 8372
rect 38612 8316 43820 8372
rect 43876 8316 43886 8372
rect 14364 8148 14420 8316
rect 14578 8204 14588 8260
rect 14644 8204 17556 8260
rect 19506 8204 19516 8260
rect 19572 8204 20524 8260
rect 20580 8204 20590 8260
rect 34738 8204 34748 8260
rect 34804 8204 35756 8260
rect 35812 8204 37660 8260
rect 37716 8204 37726 8260
rect 41682 8204 41692 8260
rect 41748 8204 45388 8260
rect 45444 8204 45454 8260
rect 17500 8148 17556 8204
rect 10770 8092 10780 8148
rect 10836 8092 12236 8148
rect 12292 8092 12572 8148
rect 12628 8092 12638 8148
rect 14364 8092 15260 8148
rect 15316 8092 15326 8148
rect 17500 8092 20972 8148
rect 21028 8092 23660 8148
rect 23716 8092 23726 8148
rect 25218 8092 25228 8148
rect 25284 8092 35196 8148
rect 35252 8092 36092 8148
rect 36148 8092 36158 8148
rect 37538 8092 37548 8148
rect 37604 8092 40572 8148
rect 40628 8092 42364 8148
rect 42420 8092 43148 8148
rect 43204 8092 43214 8148
rect 16482 7980 16492 8036
rect 16548 7980 20412 8036
rect 20468 7980 22652 8036
rect 22708 7980 22718 8036
rect 28802 7980 28812 8036
rect 28868 7980 29932 8036
rect 29988 7980 29998 8036
rect 37202 7980 37212 8036
rect 37268 7980 37884 8036
rect 37940 7980 37950 8036
rect 12786 7868 12796 7924
rect 12852 7868 15148 7924
rect 17042 7868 17052 7924
rect 17108 7868 18060 7924
rect 18116 7868 18126 7924
rect 22754 7868 22764 7924
rect 22820 7868 24724 7924
rect 7410 7756 7420 7812
rect 7476 7756 13580 7812
rect 13636 7756 14028 7812
rect 14084 7756 14094 7812
rect 15092 7700 15148 7868
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 24668 7812 24724 7868
rect 20188 7756 23716 7812
rect 24668 7756 37212 7812
rect 37268 7756 38836 7812
rect 20188 7700 20244 7756
rect 23660 7700 23716 7756
rect 1698 7644 1708 7700
rect 1764 7644 3388 7700
rect 4274 7644 4284 7700
rect 4340 7644 7532 7700
rect 7588 7644 7598 7700
rect 8194 7644 8204 7700
rect 8260 7644 9324 7700
rect 9380 7644 9390 7700
rect 15092 7644 16380 7700
rect 16436 7644 16446 7700
rect 16706 7644 16716 7700
rect 16772 7644 20244 7700
rect 21298 7644 21308 7700
rect 21364 7644 23436 7700
rect 23492 7644 23502 7700
rect 23660 7644 30940 7700
rect 30996 7644 31006 7700
rect 32498 7644 32508 7700
rect 32564 7644 34972 7700
rect 35028 7644 35038 7700
rect 35522 7644 35532 7700
rect 35588 7644 36652 7700
rect 36708 7644 37884 7700
rect 37940 7644 37950 7700
rect 3332 7364 3388 7644
rect 38780 7588 38836 7756
rect 17714 7532 17724 7588
rect 17780 7532 18284 7588
rect 18340 7532 18350 7588
rect 19618 7532 19628 7588
rect 19684 7532 24220 7588
rect 24276 7532 25676 7588
rect 25732 7532 25742 7588
rect 29698 7532 29708 7588
rect 29764 7532 34076 7588
rect 34132 7532 34142 7588
rect 38770 7532 38780 7588
rect 38836 7532 42476 7588
rect 42532 7532 44268 7588
rect 44324 7532 44334 7588
rect 45042 7532 45052 7588
rect 45108 7532 46956 7588
rect 47012 7532 47628 7588
rect 47684 7532 48300 7588
rect 48356 7532 48366 7588
rect 10434 7420 10444 7476
rect 10500 7420 11788 7476
rect 11844 7420 11854 7476
rect 13906 7420 13916 7476
rect 13972 7420 15876 7476
rect 18834 7420 18844 7476
rect 18900 7420 20748 7476
rect 20804 7420 20814 7476
rect 24994 7420 25004 7476
rect 25060 7420 26460 7476
rect 26516 7420 26526 7476
rect 26898 7420 26908 7476
rect 26964 7420 27468 7476
rect 27524 7420 32508 7476
rect 32564 7420 32574 7476
rect 43138 7420 43148 7476
rect 43204 7420 45500 7476
rect 45556 7420 45566 7476
rect 3332 7308 4732 7364
rect 4788 7308 5180 7364
rect 5236 7308 6076 7364
rect 6132 7308 7196 7364
rect 7252 7308 8540 7364
rect 8596 7308 8988 7364
rect 9044 7308 9772 7364
rect 9828 7308 9838 7364
rect 15820 7252 15876 7420
rect 16034 7308 16044 7364
rect 16100 7308 17276 7364
rect 17332 7308 17342 7364
rect 20402 7308 20412 7364
rect 20468 7308 22092 7364
rect 22148 7308 22158 7364
rect 11554 7196 11564 7252
rect 11620 7196 12124 7252
rect 12180 7196 12572 7252
rect 12628 7196 12638 7252
rect 15810 7196 15820 7252
rect 15876 7196 18060 7252
rect 18116 7196 21084 7252
rect 21140 7196 21150 7252
rect 23202 7196 23212 7252
rect 23268 7196 25564 7252
rect 25620 7196 25630 7252
rect 40226 7196 40236 7252
rect 40292 7196 41580 7252
rect 41636 7196 41646 7252
rect 14914 7084 14924 7140
rect 14980 7084 15372 7140
rect 15428 7084 16716 7140
rect 16772 7084 16782 7140
rect 18386 7084 18396 7140
rect 18452 7084 21420 7140
rect 21476 7084 21486 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 8978 6972 8988 7028
rect 9044 6972 12460 7028
rect 12516 6972 12526 7028
rect 12674 6972 12684 7028
rect 12740 6972 19012 7028
rect 25778 6972 25788 7028
rect 25844 6972 26908 7028
rect 26964 6972 26974 7028
rect 10210 6860 10220 6916
rect 10276 6860 15148 6916
rect 15474 6860 15484 6916
rect 15540 6860 18732 6916
rect 18788 6860 18798 6916
rect 8194 6748 8204 6804
rect 8260 6748 8540 6804
rect 8596 6748 8606 6804
rect 11778 6748 11788 6804
rect 11844 6748 14588 6804
rect 14644 6748 14654 6804
rect 15092 6692 15148 6860
rect 18956 6804 19012 6972
rect 18946 6748 18956 6804
rect 19012 6748 19022 6804
rect 23314 6748 23324 6804
rect 23380 6748 29764 6804
rect 43138 6748 43148 6804
rect 43204 6748 46844 6804
rect 46900 6748 46910 6804
rect 29708 6692 29764 6748
rect 9874 6636 9884 6692
rect 9940 6636 10668 6692
rect 10724 6636 10734 6692
rect 11330 6636 11340 6692
rect 11396 6636 14140 6692
rect 14196 6636 14206 6692
rect 15092 6636 17444 6692
rect 18610 6636 18620 6692
rect 18676 6636 20188 6692
rect 20244 6636 20254 6692
rect 20738 6636 20748 6692
rect 20804 6636 26124 6692
rect 26180 6636 26190 6692
rect 26450 6636 26460 6692
rect 26516 6636 26796 6692
rect 26852 6636 28084 6692
rect 28354 6636 28364 6692
rect 28420 6636 29148 6692
rect 29204 6636 29214 6692
rect 29708 6636 32620 6692
rect 32676 6636 32686 6692
rect 36082 6636 36092 6692
rect 36148 6636 37548 6692
rect 37604 6636 37614 6692
rect 42354 6636 42364 6692
rect 42420 6636 43708 6692
rect 43764 6636 43774 6692
rect 44818 6636 44828 6692
rect 44884 6636 45052 6692
rect 45108 6636 47180 6692
rect 47236 6636 48188 6692
rect 48244 6636 48254 6692
rect 6738 6524 6748 6580
rect 6804 6524 7532 6580
rect 7588 6524 7598 6580
rect 9650 6524 9660 6580
rect 9716 6524 14476 6580
rect 14532 6524 14542 6580
rect 14700 6524 15036 6580
rect 15092 6524 17164 6580
rect 17220 6524 17230 6580
rect 2482 6412 2492 6468
rect 2548 6412 3612 6468
rect 3668 6412 3678 6468
rect 7074 6412 7084 6468
rect 7140 6412 12236 6468
rect 12292 6412 12302 6468
rect 14700 6356 14756 6524
rect 17388 6468 17444 6636
rect 28028 6580 28084 6636
rect 18386 6524 18396 6580
rect 18452 6524 20300 6580
rect 20356 6524 20366 6580
rect 23538 6524 23548 6580
rect 23604 6524 25004 6580
rect 25060 6524 25070 6580
rect 26338 6524 26348 6580
rect 26404 6524 27804 6580
rect 27860 6524 27870 6580
rect 28028 6524 29260 6580
rect 29316 6524 29326 6580
rect 36306 6524 36316 6580
rect 36372 6524 37100 6580
rect 37156 6524 37166 6580
rect 45938 6524 45948 6580
rect 46004 6524 47516 6580
rect 47572 6524 48300 6580
rect 48356 6524 48366 6580
rect 17388 6412 22092 6468
rect 22148 6412 22158 6468
rect 23762 6412 23772 6468
rect 23828 6412 25228 6468
rect 25284 6412 26908 6468
rect 28018 6412 28028 6468
rect 28084 6412 29820 6468
rect 29876 6412 29886 6468
rect 33506 6412 33516 6468
rect 33572 6412 35196 6468
rect 35252 6412 35262 6468
rect 35970 6412 35980 6468
rect 36036 6412 38668 6468
rect 38724 6412 39788 6468
rect 39844 6412 39854 6468
rect 26852 6356 26908 6412
rect 9986 6300 9996 6356
rect 10052 6300 14756 6356
rect 15138 6300 15148 6356
rect 15204 6300 19180 6356
rect 19236 6300 19246 6356
rect 20178 6300 20188 6356
rect 20244 6300 23212 6356
rect 23268 6300 23884 6356
rect 23940 6300 23950 6356
rect 24098 6300 24108 6356
rect 24164 6300 25340 6356
rect 25396 6300 25406 6356
rect 26852 6300 32060 6356
rect 32116 6300 38668 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 23884 6244 23940 6300
rect 38612 6244 38668 6300
rect 8754 6188 8764 6244
rect 8820 6188 9212 6244
rect 9268 6188 18732 6244
rect 18788 6188 18798 6244
rect 23884 6188 24668 6244
rect 24724 6188 24734 6244
rect 38612 6188 39004 6244
rect 39060 6188 39070 6244
rect 4722 6076 4732 6132
rect 4788 6076 5180 6132
rect 5236 6076 5246 6132
rect 8978 6076 8988 6132
rect 9044 6076 11004 6132
rect 11060 6076 11070 6132
rect 16930 6076 16940 6132
rect 16996 6076 17724 6132
rect 17780 6076 20356 6132
rect 22530 6076 22540 6132
rect 22596 6076 23996 6132
rect 24052 6076 24062 6132
rect 24434 6076 24444 6132
rect 24500 6076 25452 6132
rect 25508 6076 25518 6132
rect 26852 6076 32172 6132
rect 32228 6076 36988 6132
rect 37044 6076 37054 6132
rect 43250 6076 43260 6132
rect 43316 6076 44156 6132
rect 44212 6076 44940 6132
rect 44996 6076 45006 6132
rect 20300 6020 20356 6076
rect 24444 6020 24500 6076
rect 15026 5964 15036 6020
rect 15092 5964 19068 6020
rect 19124 5964 19134 6020
rect 20300 5964 24500 6020
rect 8866 5852 8876 5908
rect 8932 5852 9884 5908
rect 9940 5852 11004 5908
rect 11060 5852 11070 5908
rect 18722 5852 18732 5908
rect 18788 5852 20636 5908
rect 20692 5852 20702 5908
rect 25778 5852 25788 5908
rect 25844 5852 26740 5908
rect 26684 5796 26740 5852
rect 26852 5796 26908 6076
rect 28242 5964 28252 6020
rect 28308 5964 31052 6020
rect 31108 5964 31118 6020
rect 38546 5964 38556 6020
rect 38612 5964 39676 6020
rect 39732 5964 42028 6020
rect 42084 5964 42924 6020
rect 42980 5964 42990 6020
rect 31938 5852 31948 5908
rect 32004 5852 32508 5908
rect 32564 5852 34076 5908
rect 34132 5852 34142 5908
rect 14354 5740 14364 5796
rect 14420 5740 15484 5796
rect 15540 5740 19740 5796
rect 19796 5740 20748 5796
rect 20804 5740 21196 5796
rect 21252 5740 21756 5796
rect 21812 5740 21822 5796
rect 24546 5740 24556 5796
rect 24612 5740 26012 5796
rect 26068 5740 26078 5796
rect 26674 5740 26684 5796
rect 26740 5740 26908 5796
rect 3042 5628 3052 5684
rect 3108 5628 3724 5684
rect 3780 5628 3790 5684
rect 11778 5628 11788 5684
rect 11844 5628 17388 5684
rect 17444 5628 17454 5684
rect 19282 5628 19292 5684
rect 19348 5628 25228 5684
rect 25284 5628 25294 5684
rect 28802 5628 28812 5684
rect 28868 5628 31724 5684
rect 31780 5628 31790 5684
rect 9762 5516 9772 5572
rect 9828 5516 15596 5572
rect 15652 5516 15662 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 10658 5404 10668 5460
rect 10724 5404 16268 5460
rect 16324 5404 16334 5460
rect 3714 5292 3724 5348
rect 3780 5292 4732 5348
rect 4788 5292 4798 5348
rect 10434 5292 10444 5348
rect 10500 5292 12348 5348
rect 12404 5292 12414 5348
rect 37090 5292 37100 5348
rect 37156 5292 37996 5348
rect 38052 5292 38062 5348
rect 3490 5180 3500 5236
rect 3556 5180 7588 5236
rect 14802 5180 14812 5236
rect 14868 5180 18732 5236
rect 18788 5180 18798 5236
rect 28354 5180 28364 5236
rect 28420 5180 30044 5236
rect 30100 5180 30110 5236
rect 34066 5180 34076 5236
rect 34132 5180 34636 5236
rect 34692 5180 35532 5236
rect 35588 5180 35598 5236
rect 7532 5124 7588 5180
rect 1922 5068 1932 5124
rect 1988 5068 3836 5124
rect 3892 5068 3902 5124
rect 7522 5068 7532 5124
rect 7588 5068 10444 5124
rect 10500 5068 10510 5124
rect 12898 5068 12908 5124
rect 12964 5068 13860 5124
rect 14354 5068 14364 5124
rect 14420 5068 16380 5124
rect 16436 5068 16446 5124
rect 19282 5068 19292 5124
rect 19348 5068 21420 5124
rect 21476 5068 21486 5124
rect 22418 5068 22428 5124
rect 22484 5068 27580 5124
rect 27636 5068 27646 5124
rect 28578 5068 28588 5124
rect 28644 5068 29260 5124
rect 29316 5068 29326 5124
rect 30156 5068 30828 5124
rect 30884 5068 33628 5124
rect 33684 5068 35084 5124
rect 35140 5068 35150 5124
rect 38434 5068 38444 5124
rect 38500 5068 42140 5124
rect 42196 5068 42206 5124
rect 2706 4956 2716 5012
rect 2772 4956 7420 5012
rect 7476 4956 7486 5012
rect 11890 4956 11900 5012
rect 11956 4956 13580 5012
rect 13636 4956 13646 5012
rect 13804 4900 13860 5068
rect 30156 5012 30212 5068
rect 18498 4956 18508 5012
rect 18564 4956 23212 5012
rect 23268 4956 24780 5012
rect 24836 4956 24846 5012
rect 26852 4956 29596 5012
rect 29652 4956 30212 5012
rect 38770 4956 38780 5012
rect 38836 4956 39452 5012
rect 39508 4956 39518 5012
rect 26852 4900 26908 4956
rect 7634 4844 7644 4900
rect 7700 4844 13468 4900
rect 13524 4844 13534 4900
rect 13804 4844 26908 4900
rect 31378 4844 31388 4900
rect 31444 4844 33740 4900
rect 33796 4844 33806 4900
rect 25218 4732 25228 4788
rect 25284 4732 33292 4788
rect 33348 4732 33358 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 5730 4508 5740 4564
rect 5796 4508 11788 4564
rect 11844 4508 11854 4564
rect 15092 4508 26908 4564
rect 15092 4452 15148 4508
rect 10546 4396 10556 4452
rect 10612 4396 15148 4452
rect 17490 4396 17500 4452
rect 17556 4396 20188 4452
rect 20244 4396 20972 4452
rect 21028 4396 21038 4452
rect 24882 4396 24892 4452
rect 24948 4396 26236 4452
rect 26292 4396 26302 4452
rect 8194 4284 8204 4340
rect 8260 4284 10220 4340
rect 10276 4284 11228 4340
rect 11284 4284 11294 4340
rect 21522 4284 21532 4340
rect 21588 4284 25900 4340
rect 25956 4284 25966 4340
rect 26852 4284 26908 4508
rect 32274 4396 32284 4452
rect 32340 4396 34860 4452
rect 34916 4396 34926 4452
rect 39106 4396 39116 4452
rect 39172 4396 40012 4452
rect 40068 4396 40078 4452
rect 40338 4396 40348 4452
rect 40404 4396 43260 4452
rect 43316 4396 43326 4452
rect 26964 4284 26974 4340
rect 41010 4284 41020 4340
rect 41076 4284 43820 4340
rect 43876 4284 43886 4340
rect 25900 4228 25956 4284
rect 24658 4172 24668 4228
rect 24724 4172 25676 4228
rect 25732 4172 25742 4228
rect 25900 4172 28364 4228
rect 28420 4172 28430 4228
rect 19954 4060 19964 4116
rect 20020 4060 25340 4116
rect 25396 4060 25406 4116
rect 26674 4060 26684 4116
rect 26740 4060 27916 4116
rect 27972 4060 27982 4116
rect 28914 4060 28924 4116
rect 28980 4060 30044 4116
rect 30100 4060 30110 4116
rect 33394 4060 33404 4116
rect 33460 4060 35308 4116
rect 35364 4060 35374 4116
rect 7186 3948 7196 4004
rect 7252 3948 14476 4004
rect 14532 3948 14542 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 5506 3836 5516 3892
rect 5572 3836 11116 3892
rect 11172 3836 11182 3892
rect 11340 3836 15372 3892
rect 15428 3836 15438 3892
rect 31154 3836 31164 3892
rect 31220 3836 34412 3892
rect 34468 3836 34478 3892
rect 11340 3780 11396 3836
rect 3266 3724 3276 3780
rect 3332 3724 3724 3780
rect 3780 3724 5628 3780
rect 5684 3724 5694 3780
rect 6962 3724 6972 3780
rect 7028 3724 11396 3780
rect 14130 3724 14140 3780
rect 14196 3724 16828 3780
rect 16884 3724 16894 3780
rect 17378 3724 17388 3780
rect 17444 3724 20748 3780
rect 20804 3724 20814 3780
rect 21074 3724 21084 3780
rect 21140 3724 22092 3780
rect 22148 3724 24556 3780
rect 24612 3724 24622 3780
rect 3154 3612 3164 3668
rect 3220 3612 4284 3668
rect 4340 3612 4350 3668
rect 8306 3612 8316 3668
rect 8372 3612 9324 3668
rect 9380 3612 9390 3668
rect 13234 3612 13244 3668
rect 13300 3612 15708 3668
rect 15764 3612 15774 3668
rect 27794 3612 27804 3668
rect 27860 3612 29372 3668
rect 29428 3612 29438 3668
rect 34514 3612 34524 3668
rect 34580 3612 36988 3668
rect 37044 3612 37054 3668
rect 37874 3612 37884 3668
rect 37940 3612 40796 3668
rect 40852 3612 40862 3668
rect 42354 3612 42364 3668
rect 42420 3612 44604 3668
rect 44660 3612 44670 3668
rect 3378 3500 3388 3556
rect 3444 3500 5964 3556
rect 6020 3500 6030 3556
rect 7868 3500 21420 3556
rect 21476 3500 21486 3556
rect 29138 3500 29148 3556
rect 29204 3500 31276 3556
rect 31332 3500 31342 3556
rect 33964 3500 36428 3556
rect 36484 3500 36494 3556
rect 37090 3500 37100 3556
rect 37156 3500 39788 3556
rect 39844 3500 39854 3556
rect 42466 3500 42476 3556
rect 42532 3500 43596 3556
rect 43652 3500 43662 3556
rect 7868 3444 7924 3500
rect 4050 3388 4060 3444
rect 4116 3388 6188 3444
rect 6244 3388 6254 3444
rect 7858 3388 7868 3444
rect 7924 3388 7934 3444
rect 12450 3388 12460 3444
rect 12516 3388 13580 3444
rect 13636 3388 13646 3444
rect 20178 3388 20188 3444
rect 20244 3388 25228 3444
rect 25284 3388 25294 3444
rect 30034 3388 30044 3444
rect 30100 3388 33740 3444
rect 33796 3388 33806 3444
rect 33964 3332 34020 3500
rect 43474 3388 43484 3444
rect 43540 3388 46508 3444
rect 46564 3388 46574 3444
rect 4386 3276 4396 3332
rect 4452 3276 34020 3332
rect 36754 3276 36764 3332
rect 36820 3276 38892 3332
rect 38948 3276 38958 3332
rect 40114 3276 40124 3332
rect 40180 3276 42700 3332
rect 42756 3276 42766 3332
rect 45714 3276 45724 3332
rect 45780 3276 47404 3332
rect 47460 3276 47470 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 7746 2940 7756 2996
rect 7812 2940 38444 2996
rect 38500 2940 38510 2996
<< via3 >>
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 17836 41244 17892 41300
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 19068 38780 19124 38836
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 17836 38220 17892 38276
rect 20188 37996 20244 38052
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 29820 37212 29876 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19068 36652 19124 36708
rect 29372 36316 29428 36372
rect 29932 36316 29988 36372
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 19628 35980 19684 36036
rect 20188 35980 20244 36036
rect 29820 35420 29876 35476
rect 19628 35308 19684 35364
rect 28476 35308 28532 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 26012 35196 26068 35252
rect 29932 35084 29988 35140
rect 12236 34972 12292 35028
rect 19628 34860 19684 34916
rect 27804 34748 27860 34804
rect 30828 34524 30884 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 28476 34412 28532 34468
rect 29372 34300 29428 34356
rect 17836 33964 17892 34020
rect 27804 33964 27860 34020
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 20300 33292 20356 33348
rect 12460 32956 12516 33012
rect 12908 32956 12964 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 13468 32844 13524 32900
rect 12236 32620 12292 32676
rect 27916 32620 27972 32676
rect 18956 32396 19012 32452
rect 20300 32396 20356 32452
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 27916 31724 27972 31780
rect 20300 31612 20356 31668
rect 19404 31500 19460 31556
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19628 30156 19684 30212
rect 25900 29932 25956 29988
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 17836 29260 17892 29316
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 36428 29036 36484 29092
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 13468 28924 13524 28980
rect 18956 28812 19012 28868
rect 37436 28812 37492 28868
rect 9884 28700 9940 28756
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 26012 27580 26068 27636
rect 21756 27468 21812 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 9884 27356 9940 27412
rect 14924 27132 14980 27188
rect 19404 27132 19460 27188
rect 31836 27132 31892 27188
rect 20748 27020 20804 27076
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 21532 26684 21588 26740
rect 20748 26572 20804 26628
rect 22204 26460 22260 26516
rect 27916 26236 27972 26292
rect 9884 26124 9940 26180
rect 14924 25900 14980 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 30828 25788 30884 25844
rect 9212 25452 9268 25508
rect 27916 25228 27972 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 21532 25004 21588 25060
rect 21756 25004 21812 25060
rect 22204 24892 22260 24948
rect 12460 24556 12516 24612
rect 13468 24556 13524 24612
rect 31948 24332 32004 24388
rect 36092 24332 36148 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 36204 24220 36260 24276
rect 9884 23996 9940 24052
rect 36652 23996 36708 24052
rect 12908 23884 12964 23940
rect 9884 23772 9940 23828
rect 26796 23772 26852 23828
rect 25228 23660 25284 23716
rect 26236 23660 26292 23716
rect 36204 23660 36260 23716
rect 9212 23548 9268 23604
rect 36092 23548 36148 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 36428 23492 36484 23548
rect 25228 22988 25284 23044
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 27356 22652 27412 22708
rect 36988 22652 37044 22708
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 20524 21420 20580 21476
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 32284 20972 32340 21028
rect 32844 20972 32900 21028
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 34412 19964 34468 20020
rect 32844 19628 32900 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 27692 19068 27748 19124
rect 32284 19068 32340 19124
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 26796 18060 26852 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 27020 17836 27076 17892
rect 34860 17836 34916 17892
rect 27244 17724 27300 17780
rect 35980 17724 36036 17780
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 27020 17052 27076 17108
rect 27356 16828 27412 16884
rect 37884 16828 37940 16884
rect 27244 16716 27300 16772
rect 36204 16716 36260 16772
rect 36652 16716 36708 16772
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 36092 15932 36148 15988
rect 36988 15932 37044 15988
rect 27020 15820 27076 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 25900 15372 25956 15428
rect 37212 15372 37268 15428
rect 35644 15260 35700 15316
rect 35644 14924 35700 14980
rect 37884 14924 37940 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 36204 14812 36260 14868
rect 35980 14476 36036 14532
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 37212 14028 37268 14084
rect 34076 13692 34132 13748
rect 36092 13692 36148 13748
rect 20524 13356 20580 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 26236 12684 26292 12740
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 34076 12460 34132 12516
rect 34412 12460 34468 12516
rect 37324 12348 37380 12404
rect 27692 12236 27748 12292
rect 34860 11900 34916 11956
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 49420 4768 50236
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 19808 50204 20128 50236
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 17836 41300 17892 41310
rect 17836 38276 17892 41244
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 17836 38210 17892 38220
rect 19068 38836 19124 38846
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 19068 36708 19124 38780
rect 19068 36642 19124 36652
rect 19808 37660 20128 39172
rect 35168 49420 35488 50236
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 19628 36036 19684 36046
rect 19628 35364 19684 35980
rect 19628 35298 19684 35308
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 12236 35028 12292 35038
rect 12236 32676 12292 34972
rect 19628 34916 19684 34926
rect 17836 34020 17892 34030
rect 12236 32610 12292 32620
rect 12460 33012 12516 33022
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 9884 28756 9940 28766
rect 9884 27412 9940 28700
rect 9884 27346 9940 27356
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 9884 26180 9940 26190
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 9212 25508 9268 25518
rect 9212 23604 9268 25452
rect 9884 24052 9940 26124
rect 12460 24612 12516 32956
rect 12460 24546 12516 24556
rect 12908 33012 12964 33022
rect 9884 23828 9940 23996
rect 12908 23940 12964 32956
rect 13468 32900 13524 32910
rect 13468 28980 13524 32844
rect 17836 29316 17892 33964
rect 17836 29250 17892 29260
rect 18956 32452 19012 32462
rect 13468 24612 13524 28924
rect 18956 28868 19012 32396
rect 18956 28802 19012 28812
rect 19404 31556 19460 31566
rect 14924 27188 14980 27198
rect 14924 25956 14980 27132
rect 19404 27188 19460 31500
rect 19628 30212 19684 34860
rect 19628 30146 19684 30156
rect 19808 34524 20128 36036
rect 20188 38052 20244 38062
rect 20188 36036 20244 37996
rect 29820 37268 29876 37278
rect 20188 35970 20244 35980
rect 29372 36372 29428 36382
rect 28476 35364 28532 35374
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 26012 35252 26068 35262
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 20300 33348 20356 33358
rect 20300 32452 20356 33292
rect 20300 31668 20356 32396
rect 20300 31602 20356 31612
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19404 27122 19460 27132
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 14924 25890 14980 25900
rect 19808 26684 20128 28196
rect 25900 29988 25956 29998
rect 21756 27524 21812 27534
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 13468 24546 13524 24556
rect 19808 25116 20128 26628
rect 20748 27076 20804 27086
rect 20748 26628 20804 27020
rect 20748 26562 20804 26572
rect 21532 26740 21588 26750
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 12908 23874 12964 23884
rect 9884 23762 9940 23772
rect 9212 23538 9268 23548
rect 19808 23548 20128 25060
rect 21532 25060 21588 26684
rect 21532 24994 21588 25004
rect 21756 25060 21812 27468
rect 21756 24994 21812 25004
rect 22204 26516 22260 26526
rect 22204 24948 22260 26460
rect 22204 24882 22260 24892
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 25228 23716 25284 23726
rect 25228 23044 25284 23660
rect 25228 22978 25284 22988
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 20524 21476 20580 21486
rect 20524 13412 20580 21420
rect 25900 15428 25956 29932
rect 26012 27636 26068 35196
rect 27804 34804 27860 34814
rect 27804 34020 27860 34748
rect 28476 34468 28532 35308
rect 28476 34402 28532 34412
rect 29372 34356 29428 36316
rect 29820 35476 29876 37212
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 29820 35410 29876 35420
rect 29932 36372 29988 36382
rect 29932 35140 29988 36316
rect 29932 35074 29988 35084
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 29372 34290 29428 34300
rect 30828 34580 30884 34590
rect 27804 33954 27860 33964
rect 27916 32676 27972 32686
rect 27916 31780 27972 32620
rect 27916 31714 27972 31724
rect 26012 27570 26068 27580
rect 27916 26292 27972 26302
rect 27916 25284 27972 26236
rect 30828 25844 30884 34524
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 31836 27188 31892 27198
rect 31836 26908 31892 27132
rect 31836 26852 32004 26908
rect 30828 25778 30884 25788
rect 27916 25218 27972 25228
rect 31948 24388 32004 26852
rect 31948 24322 32004 24332
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 36428 29092 36484 29102
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 26796 23828 26852 23838
rect 25900 15362 25956 15372
rect 26236 23716 26292 23726
rect 20524 13346 20580 13356
rect 26236 12740 26292 23660
rect 26796 18116 26852 23772
rect 35168 22764 35488 24276
rect 36092 24388 36148 24398
rect 36092 23604 36148 24332
rect 36204 24276 36260 24286
rect 36204 23716 36260 24220
rect 36204 23650 36260 23660
rect 36092 23538 36148 23548
rect 36428 23548 36484 29036
rect 37436 28868 37492 28878
rect 37436 26908 37492 28812
rect 37324 26852 37492 26908
rect 36428 23482 36484 23492
rect 36652 24052 36708 24062
rect 26796 18050 26852 18060
rect 27356 22708 27412 22718
rect 27020 17892 27076 17902
rect 27020 17108 27076 17836
rect 27020 15876 27076 17052
rect 27244 17780 27300 17790
rect 27244 16772 27300 17724
rect 27356 16884 27412 22652
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 32284 21028 32340 21038
rect 27356 16818 27412 16828
rect 27692 19124 27748 19134
rect 27244 16706 27300 16716
rect 27020 15810 27076 15820
rect 26236 12674 26292 12684
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 27692 12292 27748 19068
rect 32284 19124 32340 20972
rect 32844 21028 32900 21038
rect 32844 19684 32900 20972
rect 32844 19618 32900 19628
rect 34412 20020 34468 20030
rect 32284 19058 32340 19068
rect 34076 13748 34132 13758
rect 34076 12516 34132 13692
rect 34076 12450 34132 12460
rect 34412 12516 34468 19964
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 34412 12450 34468 12460
rect 34860 17892 34916 17902
rect 27692 12226 27748 12236
rect 34860 11956 34916 17836
rect 34860 11890 34916 11900
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35980 17780 36036 17790
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35644 15316 35700 15326
rect 35644 14980 35700 15260
rect 35644 14914 35700 14924
rect 35168 13356 35488 14868
rect 35980 14532 36036 17724
rect 36204 16772 36260 16782
rect 35980 14466 36036 14476
rect 36092 15988 36148 15998
rect 36092 13748 36148 15932
rect 36204 14868 36260 16716
rect 36652 16772 36708 23996
rect 36652 16706 36708 16716
rect 36988 22708 37044 22718
rect 36988 15988 37044 22652
rect 36988 15922 37044 15932
rect 36204 14802 36260 14812
rect 37212 15428 37268 15438
rect 37212 14084 37268 15372
rect 37212 14018 37268 14028
rect 36092 13682 36148 13692
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 11788 35488 13300
rect 37324 12404 37380 26852
rect 37884 16884 37940 16894
rect 37884 14980 37940 16828
rect 37884 14914 37940 14924
rect 37324 12338 37380 12348
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0935_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6496 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0936_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0937_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34048 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0938_
timestamp 1698431365
transform -1 0 35616 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0939_
timestamp 1698431365
transform 1 0 35168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _0940_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34384 0 -1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0941_
timestamp 1698431365
transform 1 0 35616 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0942_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0943_
timestamp 1698431365
transform -1 0 29232 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0944_
timestamp 1698431365
transform 1 0 28560 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0945_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31696 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0946_
timestamp 1698431365
transform -1 0 34832 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0947_
timestamp 1698431365
transform -1 0 35952 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0948_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33824 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0949_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32928 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0950_
timestamp 1698431365
transform 1 0 33264 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0951_
timestamp 1698431365
transform 1 0 34720 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0952_
timestamp 1698431365
transform 1 0 34832 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0953_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36288 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0954_
timestamp 1698431365
transform -1 0 17024 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0955_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16688 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0956_
timestamp 1698431365
transform -1 0 39648 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0957_
timestamp 1698431365
transform 1 0 41776 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0958_
timestamp 1698431365
transform 1 0 34720 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0959_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0960_
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0961_
timestamp 1698431365
transform -1 0 41216 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0962_
timestamp 1698431365
transform 1 0 34832 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0963_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41664 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0964_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38080 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0965_
timestamp 1698431365
transform 1 0 36176 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0966_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0967_
timestamp 1698431365
transform -1 0 27888 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0968_
timestamp 1698431365
transform -1 0 27552 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0969_
timestamp 1698431365
transform 1 0 27104 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0970_
timestamp 1698431365
transform -1 0 30800 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0971_
timestamp 1698431365
transform -1 0 30576 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0972_
timestamp 1698431365
transform 1 0 22176 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _0973_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0974_
timestamp 1698431365
transform 1 0 30688 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0975_
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0976_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29568 0 -1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0977_
timestamp 1698431365
transform -1 0 36288 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0978_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0979_
timestamp 1698431365
transform -1 0 27552 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0980_
timestamp 1698431365
transform -1 0 35952 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0981_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29904 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0982_
timestamp 1698431365
transform -1 0 28672 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0983_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30128 0 -1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0984_
timestamp 1698431365
transform 1 0 31472 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0985_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0986_
timestamp 1698431365
transform 1 0 34384 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0987_
timestamp 1698431365
transform 1 0 28224 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0988_
timestamp 1698431365
transform -1 0 28784 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0989_
timestamp 1698431365
transform 1 0 28000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0990_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28784 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0991_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29232 0 1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0992_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31584 0 1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0993_
timestamp 1698431365
transform -1 0 32704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0994_
timestamp 1698431365
transform 1 0 37184 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0995_
timestamp 1698431365
transform -1 0 39088 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0996_
timestamp 1698431365
transform -1 0 27664 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0997_
timestamp 1698431365
transform 1 0 29456 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0998_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0999_
timestamp 1698431365
transform -1 0 32704 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1000_
timestamp 1698431365
transform -1 0 27552 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1001_
timestamp 1698431365
transform 1 0 38080 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1002_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31360 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1003_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27440 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1004_
timestamp 1698431365
transform -1 0 30800 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1005_
timestamp 1698431365
transform 1 0 29344 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1006_
timestamp 1698431365
transform -1 0 32032 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1007_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31696 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1008_
timestamp 1698431365
transform -1 0 34272 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1009_
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1010_
timestamp 1698431365
transform -1 0 30128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1011_
timestamp 1698431365
transform -1 0 35392 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1012_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31472 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1013_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29680 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1014_
timestamp 1698431365
transform 1 0 32704 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1015_
timestamp 1698431365
transform -1 0 41104 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1016_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38864 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1017_
timestamp 1698431365
transform 1 0 34832 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1018_
timestamp 1698431365
transform -1 0 37296 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1019_
timestamp 1698431365
transform 1 0 35392 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1020_
timestamp 1698431365
transform -1 0 37184 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1021_
timestamp 1698431365
transform 1 0 39760 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1022_
timestamp 1698431365
transform 1 0 35728 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1023_
timestamp 1698431365
transform -1 0 37744 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1024_
timestamp 1698431365
transform 1 0 35728 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1025_
timestamp 1698431365
transform -1 0 39760 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1026_
timestamp 1698431365
transform 1 0 34496 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1027_
timestamp 1698431365
transform -1 0 35840 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1028_
timestamp 1698431365
transform 1 0 39088 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1029_
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1030_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1031_
timestamp 1698431365
transform 1 0 37968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1032_
timestamp 1698431365
transform -1 0 33936 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1033_
timestamp 1698431365
transform 1 0 31136 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1034_
timestamp 1698431365
transform 1 0 32144 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1035_
timestamp 1698431365
transform 1 0 31248 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1036_
timestamp 1698431365
transform 1 0 32144 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1037_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1038_
timestamp 1698431365
transform -1 0 34720 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1039_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34832 0 -1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1040_
timestamp 1698431365
transform 1 0 31584 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1041_
timestamp 1698431365
transform 1 0 34048 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1042_
timestamp 1698431365
transform -1 0 31360 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1043_
timestamp 1698431365
transform 1 0 21504 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1044_
timestamp 1698431365
transform -1 0 29792 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1045_
timestamp 1698431365
transform -1 0 28784 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1046_
timestamp 1698431365
transform -1 0 34720 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1047_
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1048_
timestamp 1698431365
transform 1 0 25648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1049_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25760 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1050_
timestamp 1698431365
transform -1 0 31136 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1051_
timestamp 1698431365
transform -1 0 27552 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1052_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1053_
timestamp 1698431365
transform -1 0 25760 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1054_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25648 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1055_
timestamp 1698431365
transform -1 0 35952 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1056_
timestamp 1698431365
transform 1 0 31248 0 1 14112
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1057_
timestamp 1698431365
transform 1 0 32592 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1058_
timestamp 1698431365
transform -1 0 32032 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1059_
timestamp 1698431365
transform 1 0 32032 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1060_
timestamp 1698431365
transform 1 0 30688 0 1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1061_
timestamp 1698431365
transform -1 0 35616 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1062_
timestamp 1698431365
transform -1 0 34384 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1063_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1064_
timestamp 1698431365
transform -1 0 37968 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1065_
timestamp 1698431365
transform 1 0 36400 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1066_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1067_
timestamp 1698431365
transform 1 0 36848 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1068_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38192 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1069_
timestamp 1698431365
transform -1 0 38192 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1070_
timestamp 1698431365
transform -1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1071_
timestamp 1698431365
transform -1 0 30576 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1072_
timestamp 1698431365
transform -1 0 29904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1073_
timestamp 1698431365
transform -1 0 24640 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1074_
timestamp 1698431365
transform -1 0 29904 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1075_
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1076_
timestamp 1698431365
transform 1 0 30016 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1077_
timestamp 1698431365
transform 1 0 29904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1078_
timestamp 1698431365
transform 1 0 30016 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1079_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30464 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1080_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1081_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34496 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1082_
timestamp 1698431365
transform -1 0 32704 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1083_
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1084_
timestamp 1698431365
transform -1 0 29568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1085_
timestamp 1698431365
transform -1 0 12096 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1086_
timestamp 1698431365
transform -1 0 10640 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1087_
timestamp 1698431365
transform -1 0 18704 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1088_
timestamp 1698431365
transform -1 0 18480 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1089_
timestamp 1698431365
transform 1 0 30128 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1090_
timestamp 1698431365
transform 1 0 30912 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1091_
timestamp 1698431365
transform -1 0 34048 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1092_
timestamp 1698431365
transform -1 0 33936 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1093_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31360 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1094_
timestamp 1698431365
transform -1 0 34496 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1095_
timestamp 1698431365
transform 1 0 35952 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1096_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1097_
timestamp 1698431365
transform 1 0 35952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1098_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35952 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1099_
timestamp 1698431365
transform -1 0 33824 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1100_
timestamp 1698431365
transform 1 0 30688 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1101_
timestamp 1698431365
transform -1 0 30240 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1102_
timestamp 1698431365
transform 1 0 30352 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1103_
timestamp 1698431365
transform -1 0 32368 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1104_
timestamp 1698431365
transform 1 0 30800 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1105_
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1106_
timestamp 1698431365
transform 1 0 10416 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1107_
timestamp 1698431365
transform 1 0 9744 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1108_
timestamp 1698431365
transform 1 0 12208 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1109_
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1110_
timestamp 1698431365
transform -1 0 13328 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1111_
timestamp 1698431365
transform -1 0 11536 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1112_
timestamp 1698431365
transform -1 0 11424 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1113_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28448 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1114_
timestamp 1698431365
transform -1 0 28224 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1115_
timestamp 1698431365
transform 1 0 26880 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1116_
timestamp 1698431365
transform -1 0 28224 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1117_
timestamp 1698431365
transform -1 0 24752 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1118_
timestamp 1698431365
transform -1 0 24528 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1119_
timestamp 1698431365
transform -1 0 22176 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1120_
timestamp 1698431365
transform 1 0 14112 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1121_
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1122_
timestamp 1698431365
transform -1 0 16464 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1123_
timestamp 1698431365
transform 1 0 19936 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1124_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1125_
timestamp 1698431365
transform 1 0 21952 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1126_
timestamp 1698431365
transform -1 0 22176 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1127_
timestamp 1698431365
transform -1 0 21504 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1128_
timestamp 1698431365
transform 1 0 21504 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1129_
timestamp 1698431365
transform -1 0 25760 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1130_
timestamp 1698431365
transform -1 0 23296 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1131_
timestamp 1698431365
transform -1 0 25312 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1132_
timestamp 1698431365
transform 1 0 27664 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1133_
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1134_
timestamp 1698431365
transform 1 0 22288 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1135_
timestamp 1698431365
transform 1 0 22624 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1136_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1137_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22176 0 1 15680
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1138_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1139_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25872 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1140_
timestamp 1698431365
transform -1 0 18144 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1141_
timestamp 1698431365
transform -1 0 15680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1142_
timestamp 1698431365
transform -1 0 10192 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1143_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1144_
timestamp 1698431365
transform 1 0 7392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1145_
timestamp 1698431365
transform -1 0 19824 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1146_
timestamp 1698431365
transform -1 0 18704 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1147_
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1148_
timestamp 1698431365
transform 1 0 16464 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1149_
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1150_
timestamp 1698431365
transform 1 0 20608 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1151_
timestamp 1698431365
transform -1 0 22848 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1152_
timestamp 1698431365
transform 1 0 27440 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1153_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1154_
timestamp 1698431365
transform 1 0 35392 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1155_
timestamp 1698431365
transform -1 0 30688 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1156_
timestamp 1698431365
transform -1 0 28784 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1157_
timestamp 1698431365
transform -1 0 27664 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1158_
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1159_
timestamp 1698431365
transform -1 0 18256 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1160_
timestamp 1698431365
transform -1 0 30576 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1161_
timestamp 1698431365
transform 1 0 30464 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1162_
timestamp 1698431365
transform 1 0 23072 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1163_
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1164_
timestamp 1698431365
transform -1 0 24976 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1165_
timestamp 1698431365
transform -1 0 24752 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1166_
timestamp 1698431365
transform 1 0 31808 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1167_
timestamp 1698431365
transform -1 0 25760 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1168_
timestamp 1698431365
transform -1 0 23744 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1169_
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1170_
timestamp 1698431365
transform 1 0 23744 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1171_
timestamp 1698431365
transform -1 0 11984 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1172_
timestamp 1698431365
transform 1 0 9744 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1173_
timestamp 1698431365
transform -1 0 21056 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1174_
timestamp 1698431365
transform -1 0 31136 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1175_
timestamp 1698431365
transform -1 0 20832 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1176_
timestamp 1698431365
transform 1 0 19376 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1177_
timestamp 1698431365
transform -1 0 19824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1178_
timestamp 1698431365
transform 1 0 19264 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1179_
timestamp 1698431365
transform 1 0 18480 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1180_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1181_
timestamp 1698431365
transform -1 0 38192 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1182_
timestamp 1698431365
transform -1 0 38192 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1183_
timestamp 1698431365
transform -1 0 30464 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1184_
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1185_
timestamp 1698431365
transform 1 0 23968 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1186_
timestamp 1698431365
transform -1 0 14784 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1187_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26320 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1188_
timestamp 1698431365
transform 1 0 22736 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1189_
timestamp 1698431365
transform -1 0 26880 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1190_
timestamp 1698431365
transform -1 0 12656 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1191_
timestamp 1698431365
transform -1 0 25200 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1192_
timestamp 1698431365
transform 1 0 25200 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1193_
timestamp 1698431365
transform 1 0 25648 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1194_
timestamp 1698431365
transform -1 0 28336 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1195_
timestamp 1698431365
transform -1 0 30240 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1196_
timestamp 1698431365
transform -1 0 35840 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1197_
timestamp 1698431365
transform 1 0 34384 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1198_
timestamp 1698431365
transform -1 0 29680 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1199_
timestamp 1698431365
transform -1 0 28560 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1200_
timestamp 1698431365
transform -1 0 28672 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1201_
timestamp 1698431365
transform -1 0 28224 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1202_
timestamp 1698431365
transform -1 0 26880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1203_
timestamp 1698431365
transform -1 0 26768 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1204_
timestamp 1698431365
transform 1 0 25760 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1205_
timestamp 1698431365
transform 1 0 32032 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1206_
timestamp 1698431365
transform 1 0 34048 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1207_
timestamp 1698431365
transform 1 0 32928 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1208_
timestamp 1698431365
transform -1 0 23632 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1209_
timestamp 1698431365
transform 1 0 28224 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1210_
timestamp 1698431365
transform 1 0 28896 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1211_
timestamp 1698431365
transform 1 0 29568 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1212_
timestamp 1698431365
transform -1 0 34048 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1213_
timestamp 1698431365
transform -1 0 34048 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1214_
timestamp 1698431365
transform -1 0 31248 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1215_
timestamp 1698431365
transform 1 0 33936 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1216_
timestamp 1698431365
transform -1 0 32704 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1217_
timestamp 1698431365
transform 1 0 31808 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1218_
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1219_
timestamp 1698431365
transform 1 0 41440 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1220_
timestamp 1698431365
transform -1 0 44240 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1221_
timestamp 1698431365
transform -1 0 44464 0 -1 21952
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1222_
timestamp 1698431365
transform 1 0 38528 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1223_
timestamp 1698431365
transform 1 0 45584 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1224_
timestamp 1698431365
transform -1 0 31696 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1225_
timestamp 1698431365
transform -1 0 41440 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1226_
timestamp 1698431365
transform 1 0 42448 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1227_
timestamp 1698431365
transform 1 0 11984 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1228_
timestamp 1698431365
transform 1 0 44016 0 -1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1229_
timestamp 1698431365
transform 1 0 31136 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1230_
timestamp 1698431365
transform 1 0 41440 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1231_
timestamp 1698431365
transform 1 0 41328 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1232_
timestamp 1698431365
transform 1 0 40768 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1233_
timestamp 1698431365
transform -1 0 28560 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1234_
timestamp 1698431365
transform -1 0 45248 0 -1 28224
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1235_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1236_
timestamp 1698431365
transform -1 0 31248 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1237_
timestamp 1698431365
transform 1 0 25760 0 1 31360
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1238_
timestamp 1698431365
transform -1 0 18928 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1239_
timestamp 1698431365
transform 1 0 31360 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1240_
timestamp 1698431365
transform 1 0 42336 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1241_
timestamp 1698431365
transform 1 0 15120 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1242_
timestamp 1698431365
transform 1 0 19600 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1243_
timestamp 1698431365
transform 1 0 19264 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1244_
timestamp 1698431365
transform 1 0 19600 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1245_
timestamp 1698431365
transform -1 0 19152 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1246_
timestamp 1698431365
transform -1 0 30464 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1247_
timestamp 1698431365
transform 1 0 23184 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1248_
timestamp 1698431365
transform 1 0 18144 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1249_
timestamp 1698431365
transform 1 0 15904 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1250_
timestamp 1698431365
transform 1 0 19152 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1251_
timestamp 1698431365
transform 1 0 18592 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1252_
timestamp 1698431365
transform 1 0 23968 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1253_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1254_
timestamp 1698431365
transform 1 0 10192 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1255_
timestamp 1698431365
transform -1 0 14000 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1256_
timestamp 1698431365
transform -1 0 13104 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1257_
timestamp 1698431365
transform -1 0 12656 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1258_
timestamp 1698431365
transform 1 0 10640 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1259_
timestamp 1698431365
transform 1 0 9968 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1260_
timestamp 1698431365
transform -1 0 13440 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1261_
timestamp 1698431365
transform -1 0 12656 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1262_
timestamp 1698431365
transform 1 0 11424 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1263_
timestamp 1698431365
transform 1 0 18480 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1264_
timestamp 1698431365
transform -1 0 11088 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1265_
timestamp 1698431365
transform 1 0 13440 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1266_
timestamp 1698431365
transform -1 0 13104 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1267_
timestamp 1698431365
transform -1 0 15344 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1268_
timestamp 1698431365
transform -1 0 27216 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1269_
timestamp 1698431365
transform -1 0 22400 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1270_
timestamp 1698431365
transform 1 0 21616 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1271_
timestamp 1698431365
transform 1 0 18816 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1272_
timestamp 1698431365
transform -1 0 22736 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1273_
timestamp 1698431365
transform 1 0 20272 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1274_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1275_
timestamp 1698431365
transform 1 0 29680 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1276_
timestamp 1698431365
transform 1 0 29568 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1277_
timestamp 1698431365
transform 1 0 33824 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1278_
timestamp 1698431365
transform -1 0 29792 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1279_
timestamp 1698431365
transform 1 0 29792 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1280_
timestamp 1698431365
transform 1 0 31584 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1281_
timestamp 1698431365
transform 1 0 39424 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1282_
timestamp 1698431365
transform -1 0 42784 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1283_
timestamp 1698431365
transform 1 0 40544 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1284_
timestamp 1698431365
transform 1 0 40544 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1285_
timestamp 1698431365
transform -1 0 43456 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1286_
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1287_
timestamp 1698431365
transform -1 0 42672 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1288_
timestamp 1698431365
transform -1 0 42672 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1289_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42560 0 1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1290_
timestamp 1698431365
transform -1 0 28784 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1291_
timestamp 1698431365
transform 1 0 25312 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1292_
timestamp 1698431365
transform 1 0 26208 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1293_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1294_
timestamp 1698431365
transform 1 0 35392 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1295_
timestamp 1698431365
transform 1 0 36960 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1296_
timestamp 1698431365
transform -1 0 36624 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1297_
timestamp 1698431365
transform 1 0 42672 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1298_
timestamp 1698431365
transform -1 0 34608 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1299_
timestamp 1698431365
transform 1 0 34384 0 1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1300_
timestamp 1698431365
transform 1 0 30128 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1301_
timestamp 1698431365
transform -1 0 10192 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1302_
timestamp 1698431365
transform 1 0 8400 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1303_
timestamp 1698431365
transform -1 0 14000 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1304_
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1305_
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1306_
timestamp 1698431365
transform -1 0 11984 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1307_
timestamp 1698431365
transform 1 0 8176 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1308_
timestamp 1698431365
transform 1 0 9072 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1309_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9296 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1310_
timestamp 1698431365
transform -1 0 29904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1311_
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1312_
timestamp 1698431365
transform 1 0 11760 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1313_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1314_
timestamp 1698431365
transform 1 0 11200 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1315_
timestamp 1698431365
transform 1 0 9520 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1316_
timestamp 1698431365
transform 1 0 10192 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1317_
timestamp 1698431365
transform -1 0 12768 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1318_
timestamp 1698431365
transform 1 0 11424 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1319_
timestamp 1698431365
transform 1 0 13664 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1320_
timestamp 1698431365
transform 1 0 9856 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1321_
timestamp 1698431365
transform 1 0 9856 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1322_
timestamp 1698431365
transform 1 0 10864 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1323_
timestamp 1698431365
transform 1 0 9632 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1324_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32816 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1325_
timestamp 1698431365
transform 1 0 10528 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1326_
timestamp 1698431365
transform 1 0 10416 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1327_
timestamp 1698431365
transform 1 0 9296 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform 1 0 9968 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1329_
timestamp 1698431365
transform 1 0 10528 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1330_
timestamp 1698431365
transform -1 0 10304 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1331_
timestamp 1698431365
transform 1 0 9632 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1332_
timestamp 1698431365
transform 1 0 8848 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1333_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10416 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1334_
timestamp 1698431365
transform 1 0 9296 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1335_
timestamp 1698431365
transform 1 0 10528 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1336_
timestamp 1698431365
transform 1 0 10304 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1337_
timestamp 1698431365
transform 1 0 9856 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1338_
timestamp 1698431365
transform 1 0 10640 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1339_
timestamp 1698431365
transform 1 0 10416 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1340_
timestamp 1698431365
transform 1 0 11312 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1341_
timestamp 1698431365
transform -1 0 5712 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1342_
timestamp 1698431365
transform 1 0 11424 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1343_
timestamp 1698431365
transform 1 0 12208 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1344_
timestamp 1698431365
transform 1 0 13104 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1345_
timestamp 1698431365
transform 1 0 16016 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1346_
timestamp 1698431365
transform 1 0 13440 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1347_
timestamp 1698431365
transform -1 0 15456 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1348_
timestamp 1698431365
transform -1 0 14560 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1349_
timestamp 1698431365
transform 1 0 13440 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1350_
timestamp 1698431365
transform 1 0 16912 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1351_
timestamp 1698431365
transform 1 0 16464 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1352_
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1353_
timestamp 1698431365
transform -1 0 22400 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1354_
timestamp 1698431365
transform 1 0 19488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1355_
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1356_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1357_
timestamp 1698431365
transform 1 0 22848 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1358_
timestamp 1698431365
transform -1 0 24752 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1359_
timestamp 1698431365
transform -1 0 24864 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1360_
timestamp 1698431365
transform 1 0 22400 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1361_
timestamp 1698431365
transform 1 0 22960 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1362_
timestamp 1698431365
transform 1 0 26320 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1363_
timestamp 1698431365
transform -1 0 27664 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1364_
timestamp 1698431365
transform 1 0 34496 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1365_
timestamp 1698431365
transform -1 0 29344 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1366_
timestamp 1698431365
transform -1 0 28112 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1367_
timestamp 1698431365
transform -1 0 25648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1368_
timestamp 1698431365
transform -1 0 26656 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1369_
timestamp 1698431365
transform 1 0 39424 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1370_
timestamp 1698431365
transform 1 0 38752 0 1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1371_
timestamp 1698431365
transform -1 0 27552 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1372_
timestamp 1698431365
transform 1 0 26432 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1373_
timestamp 1698431365
transform -1 0 34272 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1374_
timestamp 1698431365
transform -1 0 34160 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1375_
timestamp 1698431365
transform 1 0 41328 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1376_
timestamp 1698431365
transform -1 0 33376 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1377_
timestamp 1698431365
transform 1 0 32480 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1378_
timestamp 1698431365
transform 1 0 43344 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1379_
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1380_
timestamp 1698431365
transform 1 0 45248 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1381_
timestamp 1698431365
transform -1 0 42336 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1382_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1383_
timestamp 1698431365
transform -1 0 41888 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1384_
timestamp 1698431365
transform 1 0 42784 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1385_
timestamp 1698431365
transform -1 0 39984 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1386_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1387_
timestamp 1698431365
transform -1 0 28672 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1388_
timestamp 1698431365
transform 1 0 25200 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1389_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1390_
timestamp 1698431365
transform 1 0 24640 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1391_
timestamp 1698431365
transform -1 0 26320 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1392_
timestamp 1698431365
transform 1 0 24864 0 1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1393_
timestamp 1698431365
transform 1 0 19152 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1394_
timestamp 1698431365
transform -1 0 24864 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1395_
timestamp 1698431365
transform 1 0 25648 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1396_
timestamp 1698431365
transform -1 0 29456 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1397_
timestamp 1698431365
transform 1 0 27664 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1398_
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1399_
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1400_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1401_
timestamp 1698431365
transform 1 0 26544 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1402_
timestamp 1698431365
transform 1 0 27664 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1403_
timestamp 1698431365
transform -1 0 29456 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1404_
timestamp 1698431365
transform 1 0 31136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1405_
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1406_
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1407_
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1408_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1409_
timestamp 1698431365
transform 1 0 19712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1410_
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1411_
timestamp 1698431365
transform 1 0 17808 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1412_
timestamp 1698431365
transform -1 0 19600 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1413_
timestamp 1698431365
transform -1 0 33600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1414__1
timestamp 1698431365
transform -1 0 36064 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1415_
timestamp 1698431365
transform 1 0 13888 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1416_
timestamp 1698431365
transform 1 0 14560 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1417_
timestamp 1698431365
transform -1 0 16912 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1418_
timestamp 1698431365
transform 1 0 12432 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1419_
timestamp 1698431365
transform 1 0 20608 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1420_
timestamp 1698431365
transform 1 0 26320 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1421_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1422_
timestamp 1698431365
transform -1 0 28784 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1423_
timestamp 1698431365
transform 1 0 26320 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1424_
timestamp 1698431365
transform 1 0 25312 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1425_
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1426_
timestamp 1698431365
transform -1 0 17696 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1427_
timestamp 1698431365
transform 1 0 15792 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1428_
timestamp 1698431365
transform 1 0 17584 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1429_
timestamp 1698431365
transform 1 0 17472 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1430_
timestamp 1698431365
transform 1 0 14448 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1431_
timestamp 1698431365
transform 1 0 15680 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1432_
timestamp 1698431365
transform -1 0 17248 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1433_
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1434_
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1435_
timestamp 1698431365
transform -1 0 20832 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1436_
timestamp 1698431365
transform -1 0 19600 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1437_
timestamp 1698431365
transform -1 0 20944 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1438_
timestamp 1698431365
transform -1 0 21616 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1439_
timestamp 1698431365
transform -1 0 21952 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1440_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18480 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1441_
timestamp 1698431365
transform -1 0 19712 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1442_
timestamp 1698431365
transform 1 0 18816 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1443_
timestamp 1698431365
transform 1 0 22736 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1444_
timestamp 1698431365
transform 1 0 20832 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1445_
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1446_
timestamp 1698431365
transform -1 0 22624 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1447_
timestamp 1698431365
transform -1 0 22176 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1448_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1449_
timestamp 1698431365
transform 1 0 22512 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1450_
timestamp 1698431365
transform 1 0 20160 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1451_
timestamp 1698431365
transform -1 0 20272 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1452_
timestamp 1698431365
transform 1 0 20944 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1453_
timestamp 1698431365
transform -1 0 22736 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1454_
timestamp 1698431365
transform 1 0 22288 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1455_
timestamp 1698431365
transform 1 0 17584 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1456_
timestamp 1698431365
transform 1 0 20272 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1457_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22176 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1458_
timestamp 1698431365
transform -1 0 20832 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1459_
timestamp 1698431365
transform -1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1460_
timestamp 1698431365
transform -1 0 24528 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1461_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1462_
timestamp 1698431365
transform -1 0 17584 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1463_
timestamp 1698431365
transform -1 0 16352 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1464_
timestamp 1698431365
transform -1 0 17136 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1465_
timestamp 1698431365
transform 1 0 19152 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1466_
timestamp 1698431365
transform 1 0 13440 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1467_
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1468_
timestamp 1698431365
transform -1 0 21392 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1469_
timestamp 1698431365
transform 1 0 17248 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1470_
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1471_
timestamp 1698431365
transform 1 0 14672 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1472_
timestamp 1698431365
transform -1 0 15456 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1473_
timestamp 1698431365
transform -1 0 14672 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1474_
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1475_
timestamp 1698431365
transform 1 0 15232 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1476_
timestamp 1698431365
transform 1 0 15568 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1477_
timestamp 1698431365
transform 1 0 15680 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1478_
timestamp 1698431365
transform 1 0 18704 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1479_
timestamp 1698431365
transform 1 0 22848 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1480_
timestamp 1698431365
transform 1 0 16016 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1481_
timestamp 1698431365
transform -1 0 18592 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1482_
timestamp 1698431365
transform 1 0 17024 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1483_
timestamp 1698431365
transform 1 0 18368 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1484_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1485_
timestamp 1698431365
transform 1 0 17248 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1486_
timestamp 1698431365
transform 1 0 18256 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1487_
timestamp 1698431365
transform -1 0 20496 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1488_
timestamp 1698431365
transform -1 0 19600 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1489_
timestamp 1698431365
transform -1 0 15680 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1490_
timestamp 1698431365
transform -1 0 15568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1491_
timestamp 1698431365
transform -1 0 17136 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1492_
timestamp 1698431365
transform -1 0 14560 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1493_
timestamp 1698431365
transform -1 0 20944 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1494_
timestamp 1698431365
transform -1 0 20832 0 -1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1495_
timestamp 1698431365
transform -1 0 19712 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1496_
timestamp 1698431365
transform -1 0 16352 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1497_
timestamp 1698431365
transform 1 0 19488 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1498_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16240 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1499_
timestamp 1698431365
transform 1 0 14112 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1500_
timestamp 1698431365
transform 1 0 14224 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1501_
timestamp 1698431365
transform 1 0 12656 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1502_
timestamp 1698431365
transform -1 0 11088 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1503_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 -1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1504_
timestamp 1698431365
transform -1 0 27216 0 1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1505_
timestamp 1698431365
transform -1 0 23072 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1506_
timestamp 1698431365
transform 1 0 15456 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1507_
timestamp 1698431365
transform 1 0 7728 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1508_
timestamp 1698431365
transform -1 0 6944 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1509_
timestamp 1698431365
transform 1 0 7952 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1510_
timestamp 1698431365
transform -1 0 7952 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1511_
timestamp 1698431365
transform -1 0 23408 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1512_
timestamp 1698431365
transform -1 0 18480 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1513_
timestamp 1698431365
transform -1 0 11312 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1514_
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1515_
timestamp 1698431365
transform 1 0 9520 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1516_
timestamp 1698431365
transform 1 0 6496 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1517_
timestamp 1698431365
transform -1 0 6944 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1518_
timestamp 1698431365
transform 1 0 6272 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1519_
timestamp 1698431365
transform -1 0 6160 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1520_
timestamp 1698431365
transform 1 0 8400 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1521_
timestamp 1698431365
transform -1 0 8624 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1522_
timestamp 1698431365
transform -1 0 12320 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1523_
timestamp 1698431365
transform 1 0 9968 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1524_
timestamp 1698431365
transform -1 0 10080 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1525_
timestamp 1698431365
transform 1 0 11424 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1526_
timestamp 1698431365
transform -1 0 11424 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1527_
timestamp 1698431365
transform -1 0 17920 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1528_
timestamp 1698431365
transform -1 0 15120 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1529_
timestamp 1698431365
transform 1 0 22736 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1530_
timestamp 1698431365
transform -1 0 18592 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1531_
timestamp 1698431365
transform -1 0 14896 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1532_
timestamp 1698431365
transform -1 0 15120 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1533_
timestamp 1698431365
transform 1 0 15008 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1534_
timestamp 1698431365
transform -1 0 16576 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1535_
timestamp 1698431365
transform 1 0 16240 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1536_
timestamp 1698431365
transform 1 0 15344 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1537_
timestamp 1698431365
transform -1 0 17136 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1538_
timestamp 1698431365
transform 1 0 16016 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1539_
timestamp 1698431365
transform -1 0 15904 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1540_
timestamp 1698431365
transform -1 0 16800 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1541_
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1542_
timestamp 1698431365
transform 1 0 11760 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1543_
timestamp 1698431365
transform 1 0 13440 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1544_
timestamp 1698431365
transform 1 0 13440 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1545_
timestamp 1698431365
transform -1 0 16016 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1546_
timestamp 1698431365
transform 1 0 14224 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1547_
timestamp 1698431365
transform 1 0 17360 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1548_
timestamp 1698431365
transform 1 0 16464 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1549_
timestamp 1698431365
transform 1 0 17808 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1550_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1551_
timestamp 1698431365
transform -1 0 17920 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1552_
timestamp 1698431365
transform 1 0 17024 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1553_
timestamp 1698431365
transform -1 0 16800 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1554_
timestamp 1698431365
transform 1 0 18704 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1555_
timestamp 1698431365
transform -1 0 18704 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1556_
timestamp 1698431365
transform 1 0 20720 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1557_
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1558_
timestamp 1698431365
transform 1 0 27440 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1559_
timestamp 1698431365
transform 1 0 30128 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1560_
timestamp 1698431365
transform 1 0 27104 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1561_
timestamp 1698431365
transform 1 0 27328 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1562_
timestamp 1698431365
transform 1 0 28448 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1563_
timestamp 1698431365
transform 1 0 27776 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1564_
timestamp 1698431365
transform 1 0 30912 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1565_
timestamp 1698431365
transform 1 0 31024 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1566_
timestamp 1698431365
transform -1 0 35504 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1567_
timestamp 1698431365
transform -1 0 36176 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1568_
timestamp 1698431365
transform -1 0 40096 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1569_
timestamp 1698431365
transform 1 0 37520 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1570_
timestamp 1698431365
transform -1 0 38304 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1571_
timestamp 1698431365
transform -1 0 39200 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1572_
timestamp 1698431365
transform 1 0 39424 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1573_
timestamp 1698431365
transform 1 0 37744 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1574_
timestamp 1698431365
transform 1 0 37072 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1575_
timestamp 1698431365
transform 1 0 38528 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1576_
timestamp 1698431365
transform -1 0 38528 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1577_
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1578_
timestamp 1698431365
transform 1 0 38864 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1579_
timestamp 1698431365
transform -1 0 40320 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1580_
timestamp 1698431365
transform 1 0 42000 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1581_
timestamp 1698431365
transform 1 0 42112 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1582_
timestamp 1698431365
transform 1 0 42448 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1583_
timestamp 1698431365
transform 1 0 42672 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1584_
timestamp 1698431365
transform 1 0 42224 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1585_
timestamp 1698431365
transform -1 0 43344 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1586_
timestamp 1698431365
transform -1 0 30800 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1587_
timestamp 1698431365
transform 1 0 31024 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1588_
timestamp 1698431365
transform 1 0 31696 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1589_
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1590_
timestamp 1698431365
transform 1 0 32368 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1591_
timestamp 1698431365
transform 1 0 29680 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1592_
timestamp 1698431365
transform -1 0 30016 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1593_
timestamp 1698431365
transform 1 0 27104 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1594_
timestamp 1698431365
transform 1 0 26544 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1595_
timestamp 1698431365
transform 1 0 26992 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1596_
timestamp 1698431365
transform -1 0 27440 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1597_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1598_
timestamp 1698431365
transform -1 0 24640 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1599_
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1600_
timestamp 1698431365
transform -1 0 25200 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1601_
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1602_
timestamp 1698431365
transform -1 0 25760 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1603_
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1604_
timestamp 1698431365
transform -1 0 24640 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1605_
timestamp 1698431365
transform 1 0 18368 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1606_
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1607_
timestamp 1698431365
transform 1 0 18368 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1608_
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1609_
timestamp 1698431365
transform 1 0 18368 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1610_
timestamp 1698431365
transform 1 0 19488 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1611_
timestamp 1698431365
transform -1 0 18592 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1612_
timestamp 1698431365
transform -1 0 19488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1613_
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1614_
timestamp 1698431365
transform 1 0 22176 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1615_
timestamp 1698431365
transform -1 0 20944 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1616_
timestamp 1698431365
transform 1 0 19376 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1617_
timestamp 1698431365
transform 1 0 26992 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1618_
timestamp 1698431365
transform 1 0 21280 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1619_
timestamp 1698431365
transform -1 0 21056 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1620_
timestamp 1698431365
transform 1 0 22288 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1621_
timestamp 1698431365
transform -1 0 22512 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1622_
timestamp 1698431365
transform -1 0 23968 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1623_
timestamp 1698431365
transform 1 0 22848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1624_
timestamp 1698431365
transform -1 0 25760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1625_
timestamp 1698431365
transform 1 0 23408 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1626_
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1627_
timestamp 1698431365
transform -1 0 27328 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1628_
timestamp 1698431365
transform 1 0 27888 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1629_
timestamp 1698431365
transform -1 0 28448 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1630_
timestamp 1698431365
transform 1 0 34384 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1631_
timestamp 1698431365
transform 1 0 30464 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1632_
timestamp 1698431365
transform -1 0 31584 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1633_
timestamp 1698431365
transform 1 0 31024 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1634_
timestamp 1698431365
transform 1 0 30352 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1635_
timestamp 1698431365
transform 1 0 32816 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1636_
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1637_
timestamp 1698431365
transform 1 0 34720 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1638_
timestamp 1698431365
transform 1 0 35168 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1639_
timestamp 1698431365
transform 1 0 35168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1640_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1641_
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1642_
timestamp 1698431365
transform 1 0 38528 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1643_
timestamp 1698431365
transform 1 0 39088 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1644_
timestamp 1698431365
transform 1 0 40880 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1645_
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1646_
timestamp 1698431365
transform 1 0 42784 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1647_
timestamp 1698431365
transform 1 0 42672 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1648_
timestamp 1698431365
transform -1 0 22736 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1649_
timestamp 1698431365
transform 1 0 23632 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1650_
timestamp 1698431365
transform -1 0 47488 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1651_
timestamp 1698431365
transform 1 0 42560 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1652_
timestamp 1698431365
transform -1 0 43344 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1653_
timestamp 1698431365
transform 1 0 42672 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1654_
timestamp 1698431365
transform -1 0 43008 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1655_
timestamp 1698431365
transform 1 0 44912 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1656_
timestamp 1698431365
transform 1 0 45360 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1657_
timestamp 1698431365
transform 1 0 45472 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1658_
timestamp 1698431365
transform 1 0 44464 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1659_
timestamp 1698431365
transform -1 0 48272 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1660_
timestamp 1698431365
transform -1 0 48384 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1661_
timestamp 1698431365
transform -1 0 48496 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1662_
timestamp 1698431365
transform 1 0 46592 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1663_
timestamp 1698431365
transform -1 0 46928 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1664_
timestamp 1698431365
transform 1 0 46592 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1665_
timestamp 1698431365
transform -1 0 46592 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1666_
timestamp 1698431365
transform 1 0 24304 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1667_
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1668_
timestamp 1698431365
transform 1 0 26432 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1669_
timestamp 1698431365
transform 1 0 25872 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1670_
timestamp 1698431365
transform 1 0 45696 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1671_
timestamp 1698431365
transform -1 0 46368 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1672_
timestamp 1698431365
transform 1 0 46592 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1673_
timestamp 1698431365
transform 1 0 42784 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1674_
timestamp 1698431365
transform 1 0 43456 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1675_
timestamp 1698431365
transform 1 0 42784 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1676_
timestamp 1698431365
transform 1 0 43232 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1677_
timestamp 1698431365
transform 1 0 46368 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1678_
timestamp 1698431365
transform -1 0 46704 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1679_
timestamp 1698431365
transform 1 0 46368 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1680_
timestamp 1698431365
transform -1 0 46816 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1681_
timestamp 1698431365
transform -1 0 47600 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1682_
timestamp 1698431365
transform 1 0 46592 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1683_
timestamp 1698431365
transform -1 0 46816 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1684_
timestamp 1698431365
transform -1 0 48048 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1685_
timestamp 1698431365
transform -1 0 47824 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1686_
timestamp 1698431365
transform -1 0 47152 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1687_
timestamp 1698431365
transform -1 0 43680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1688_
timestamp 1698431365
transform 1 0 43008 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1689_
timestamp 1698431365
transform -1 0 42784 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1690_
timestamp 1698431365
transform -1 0 20384 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1691_
timestamp 1698431365
transform 1 0 38976 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1692_
timestamp 1698431365
transform 1 0 43344 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1693_
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1694_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1695_
timestamp 1698431365
transform 1 0 39872 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1696_
timestamp 1698431365
transform 1 0 42448 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1697_
timestamp 1698431365
transform 1 0 41776 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1698_
timestamp 1698431365
transform 1 0 45248 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1699_
timestamp 1698431365
transform -1 0 43232 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1700_
timestamp 1698431365
transform 1 0 37968 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1701_
timestamp 1698431365
transform 1 0 37520 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1702_
timestamp 1698431365
transform 1 0 36960 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1703_
timestamp 1698431365
transform -1 0 37072 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1704_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1705_
timestamp 1698431365
transform 1 0 37744 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1706_
timestamp 1698431365
transform 1 0 37408 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1707_
timestamp 1698431365
transform 1 0 34944 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1708_
timestamp 1698431365
transform -1 0 35616 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1709_
timestamp 1698431365
transform 1 0 21840 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1710_
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1711_
timestamp 1698431365
transform -1 0 20720 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1712_
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1713_
timestamp 1698431365
transform -1 0 20384 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1714_
timestamp 1698431365
transform 1 0 21392 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1715_
timestamp 1698431365
transform 1 0 20272 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1716_
timestamp 1698431365
transform 1 0 21504 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1717_
timestamp 1698431365
transform 1 0 20272 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1698431365
transform -1 0 22624 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1719_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1720_
timestamp 1698431365
transform -1 0 21840 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1721_
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1722_
timestamp 1698431365
transform -1 0 14672 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1723_
timestamp 1698431365
transform -1 0 12208 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1724_
timestamp 1698431365
transform 1 0 15232 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1725_
timestamp 1698431365
transform 1 0 14336 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1726_
timestamp 1698431365
transform -1 0 10640 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1727_
timestamp 1698431365
transform -1 0 15344 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1728_
timestamp 1698431365
transform 1 0 14672 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1729_
timestamp 1698431365
transform 1 0 13776 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1730_
timestamp 1698431365
transform -1 0 18144 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1731_
timestamp 1698431365
transform 1 0 13104 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1732_
timestamp 1698431365
transform -1 0 12096 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1733_
timestamp 1698431365
transform -1 0 14336 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1734_
timestamp 1698431365
transform 1 0 12768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1735_
timestamp 1698431365
transform -1 0 14000 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1736_
timestamp 1698431365
transform 1 0 12208 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1737_
timestamp 1698431365
transform 1 0 11424 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1738_
timestamp 1698431365
transform -1 0 10864 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1739_
timestamp 1698431365
transform 1 0 7840 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1740_
timestamp 1698431365
transform -1 0 7392 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1741_
timestamp 1698431365
transform 1 0 7504 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1742_
timestamp 1698431365
transform -1 0 7504 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1743_
timestamp 1698431365
transform -1 0 19264 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1744_
timestamp 1698431365
transform -1 0 6496 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1745_
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1746_
timestamp 1698431365
transform -1 0 3024 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1747_
timestamp 1698431365
transform 1 0 3584 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1748_
timestamp 1698431365
transform -1 0 3808 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1749_
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1750_
timestamp 1698431365
transform -1 0 2800 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1751_
timestamp 1698431365
transform 1 0 3920 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1752_
timestamp 1698431365
transform -1 0 2912 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1753_
timestamp 1698431365
transform -1 0 5936 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1754_
timestamp 1698431365
transform 1 0 3248 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1755_
timestamp 1698431365
transform -1 0 2688 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1756_
timestamp 1698431365
transform 1 0 3360 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1757_
timestamp 1698431365
transform -1 0 2688 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1758_
timestamp 1698431365
transform 1 0 3808 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1759_
timestamp 1698431365
transform -1 0 3024 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1760_
timestamp 1698431365
transform -1 0 9968 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1761_
timestamp 1698431365
transform 1 0 7952 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1762_
timestamp 1698431365
transform 1 0 8512 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1763_
timestamp 1698431365
transform -1 0 9744 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1764_
timestamp 1698431365
transform 1 0 3584 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1765_
timestamp 1698431365
transform -1 0 2800 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1766_
timestamp 1698431365
transform 1 0 5600 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1767_
timestamp 1698431365
transform 1 0 3584 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1768_
timestamp 1698431365
transform -1 0 3136 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1769_
timestamp 1698431365
transform -1 0 9296 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1770_
timestamp 1698431365
transform 1 0 7840 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1771_
timestamp 1698431365
transform -1 0 8848 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1772_
timestamp 1698431365
transform 1 0 7840 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1773_
timestamp 1698431365
transform 1 0 5040 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1774_
timestamp 1698431365
transform -1 0 2800 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1775_
timestamp 1698431365
transform 1 0 5040 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1776_
timestamp 1698431365
transform -1 0 3136 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1777_
timestamp 1698431365
transform 1 0 5824 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1778_
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1779_
timestamp 1698431365
transform -1 0 7056 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1780_
timestamp 1698431365
transform 1 0 3808 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1781_
timestamp 1698431365
transform -1 0 2800 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1782_
timestamp 1698431365
transform 1 0 3584 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1783_
timestamp 1698431365
transform -1 0 2688 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1784_
timestamp 1698431365
transform 1 0 5936 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1785_
timestamp 1698431365
transform 1 0 6272 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1786_
timestamp 1698431365
transform 1 0 3584 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1787_
timestamp 1698431365
transform -1 0 2688 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1788_
timestamp 1698431365
transform -1 0 21280 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1789_
timestamp 1698431365
transform -1 0 5824 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1790_
timestamp 1698431365
transform 1 0 3248 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1791_
timestamp 1698431365
transform -1 0 2688 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1792_
timestamp 1698431365
transform 1 0 3136 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1793_
timestamp 1698431365
transform -1 0 2688 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1794_
timestamp 1698431365
transform 1 0 3360 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1795_
timestamp 1698431365
transform -1 0 2688 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1796_
timestamp 1698431365
transform 1 0 3584 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1797_
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1798_
timestamp 1698431365
transform 1 0 5600 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1799_
timestamp 1698431365
transform 1 0 3584 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1800_
timestamp 1698431365
transform -1 0 2800 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1801_
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1802_
timestamp 1698431365
transform -1 0 4816 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1803_
timestamp 1698431365
transform 1 0 7168 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1804_
timestamp 1698431365
transform 1 0 7168 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1805_
timestamp 1698431365
transform 1 0 7392 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1806_
timestamp 1698431365
transform 1 0 7728 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1807_
timestamp 1698431365
transform 1 0 34608 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1808_
timestamp 1698431365
transform 1 0 7392 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1809_
timestamp 1698431365
transform -1 0 6608 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1810_
timestamp 1698431365
transform 1 0 7168 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1811_
timestamp 1698431365
transform -1 0 6832 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1812_
timestamp 1698431365
transform 1 0 7280 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1813_
timestamp 1698431365
transform -1 0 6944 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1814_
timestamp 1698431365
transform 1 0 34944 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1815_
timestamp 1698431365
transform 1 0 33264 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1816_
timestamp 1698431365
transform 1 0 37856 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1817_
timestamp 1698431365
transform 1 0 37408 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1818_
timestamp 1698431365
transform -1 0 37968 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1819_
timestamp 1698431365
transform 1 0 38864 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1820_
timestamp 1698431365
transform 1 0 39872 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1821_
timestamp 1698431365
transform 1 0 40992 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1822_
timestamp 1698431365
transform -1 0 41888 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1823_
timestamp 1698431365
transform -1 0 44352 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1824_
timestamp 1698431365
transform 1 0 43456 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1825_
timestamp 1698431365
transform 1 0 46256 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1826_
timestamp 1698431365
transform -1 0 46480 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1827_
timestamp 1698431365
transform 1 0 46368 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1828_
timestamp 1698431365
transform -1 0 46368 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1829_
timestamp 1698431365
transform -1 0 35280 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1830_
timestamp 1698431365
transform -1 0 32704 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1831_
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1832_
timestamp 1698431365
transform -1 0 34496 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1833_
timestamp 1698431365
transform -1 0 30240 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1834_
timestamp 1698431365
transform 1 0 30240 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1835_
timestamp 1698431365
transform 1 0 30240 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1836_
timestamp 1698431365
transform 1 0 33824 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1837_
timestamp 1698431365
transform 1 0 34160 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1838_
timestamp 1698431365
transform 1 0 32256 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1839_
timestamp 1698431365
transform 1 0 33264 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1840_
timestamp 1698431365
transform -1 0 33824 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1841_
timestamp 1698431365
transform -1 0 32928 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1842_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1843_
timestamp 1698431365
transform 1 0 29680 0 1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1844_
timestamp 1698431365
transform -1 0 32704 0 -1 9408
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1845_
timestamp 1698431365
transform 1 0 11536 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1846_
timestamp 1698431365
transform -1 0 10640 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1847_
timestamp 1698431365
transform -1 0 14112 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1848_
timestamp 1698431365
transform -1 0 12992 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1849_
timestamp 1698431365
transform -1 0 7280 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1850_
timestamp 1698431365
transform 1 0 22848 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1851_
timestamp 1698431365
transform -1 0 13104 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1852_
timestamp 1698431365
transform 1 0 10192 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1853_
timestamp 1698431365
transform 1 0 29456 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1854_
timestamp 1698431365
transform 1 0 30352 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1855_
timestamp 1698431365
transform 1 0 30688 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1856_
timestamp 1698431365
transform 1 0 33600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1857_
timestamp 1698431365
transform -1 0 15904 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1858_
timestamp 1698431365
transform 1 0 17920 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1859_
timestamp 1698431365
transform 1 0 20048 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1860_
timestamp 1698431365
transform 1 0 21392 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1861_
timestamp 1698431365
transform -1 0 37520 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1862_
timestamp 1698431365
transform -1 0 33600 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1863_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1864_
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1865_
timestamp 1698431365
transform 1 0 32256 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1866_
timestamp 1698431365
transform 1 0 38640 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1867_
timestamp 1698431365
transform 1 0 37184 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1868_
timestamp 1698431365
transform 1 0 36848 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1869_
timestamp 1698431365
transform 1 0 37744 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1870_
timestamp 1698431365
transform 1 0 39648 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1871_
timestamp 1698431365
transform 1 0 37072 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1872_
timestamp 1698431365
transform 1 0 37968 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1873_
timestamp 1698431365
transform -1 0 37632 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1874_
timestamp 1698431365
transform 1 0 38304 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1875_
timestamp 1698431365
transform 1 0 38976 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1876_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1877_
timestamp 1698431365
transform 1 0 37184 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1878_
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1879_
timestamp 1698431365
transform -1 0 37744 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1880_
timestamp 1698431365
transform -1 0 39984 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1881_
timestamp 1698431365
transform 1 0 36960 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1882_
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1883_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8624 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1884_
timestamp 1698431365
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1885_
timestamp 1698431365
transform 1 0 23408 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1886_
timestamp 1698431365
transform 1 0 23968 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1887_
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1888_
timestamp 1698431365
transform 1 0 11088 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1889_
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1890_
timestamp 1698431365
transform 1 0 11424 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1891_
timestamp 1698431365
transform 1 0 31696 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1892_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1893_
timestamp 1698431365
transform 1 0 17920 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1894_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1895_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 -1 36064
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1896_
timestamp 1698431365
transform 1 0 5824 0 -1 39200
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1897_
timestamp 1698431365
transform 1 0 9296 0 1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1898_
timestamp 1698431365
transform 1 0 5824 0 -1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1899_
timestamp 1698431365
transform 1 0 4480 0 -1 43904
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1900_
timestamp 1698431365
transform 1 0 7280 0 1 43904
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1901_
timestamp 1698431365
transform 1 0 8064 0 1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1902_
timestamp 1698431365
transform 1 0 9744 0 1 47040
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1903_
timestamp 1698431365
transform 1 0 12544 0 -1 39200
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1904_
timestamp 1698431365
transform 1 0 13664 0 -1 34496
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1905_
timestamp 1698431365
transform 1 0 15344 0 1 36064
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1906_
timestamp 1698431365
transform 1 0 15232 0 1 42336
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1907_
timestamp 1698431365
transform 1 0 12432 0 -1 43904
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1908_
timestamp 1698431365
transform 1 0 13104 0 -1 47040
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1909_
timestamp 1698431365
transform 1 0 12096 0 -1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1910_
timestamp 1698431365
transform 1 0 16016 0 1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1911_
timestamp 1698431365
transform 1 0 16016 0 1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1912_
timestamp 1698431365
transform 1 0 14224 0 1 48608
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1913_
timestamp 1698431365
transform 1 0 17584 0 1 48608
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1914_
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1915_
timestamp 1698431365
transform 1 0 26768 0 -1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1916_
timestamp 1698431365
transform 1 0 27552 0 -1 42336
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1917_
timestamp 1698431365
transform 1 0 30464 0 1 43904
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1918_
timestamp 1698431365
transform 1 0 34272 0 -1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1919_
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1920_
timestamp 1698431365
transform 1 0 39200 0 1 47040
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1921_
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1922_
timestamp 1698431365
transform 1 0 37520 0 1 42336
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1923_
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1924_
timestamp 1698431365
transform 1 0 41888 0 -1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1925_
timestamp 1698431365
transform 1 0 42560 0 -1 42336
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1926_
timestamp 1698431365
transform 1 0 42000 0 -1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1927_
timestamp 1698431365
transform 1 0 32368 0 1 47040
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1928_
timestamp 1698431365
transform 1 0 32592 0 1 48608
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1929_
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1930_
timestamp 1698431365
transform -1 0 28784 0 1 48608
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1931_
timestamp 1698431365
transform 1 0 23184 0 1 47040
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1932_
timestamp 1698431365
transform 1 0 23296 0 1 43904
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1933_
timestamp 1698431365
transform 1 0 23744 0 1 42336
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1934_
timestamp 1698431365
transform 1 0 23296 0 1 39200
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1935_
timestamp 1698431365
transform 1 0 16688 0 1 39200
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1936_
timestamp 1698431365
transform 1 0 15008 0 1 31360
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1937_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1938_
timestamp 1698431365
transform 1 0 18816 0 -1 28224
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1939_
timestamp 1698431365
transform 1 0 19600 0 -1 31360
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1940_
timestamp 1698431365
transform 1 0 21280 0 -1 34496
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1941_
timestamp 1698431365
transform 1 0 21504 0 -1 26656
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1942_
timestamp 1698431365
transform 1 0 24304 0 1 28224
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1943_
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1944_
timestamp 1698431365
transform 1 0 27104 0 -1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1945_
timestamp 1698431365
transform 1 0 29344 0 1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1946_
timestamp 1698431365
transform 1 0 30688 0 1 37632
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1947_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1948_
timestamp 1698431365
transform -1 0 39648 0 -1 42336
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1949_
timestamp 1698431365
transform -1 0 39088 0 -1 39200
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1950_
timestamp 1698431365
transform -1 0 40544 0 -1 37632
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1951_
timestamp 1698431365
transform 1 0 40544 0 1 37632
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1952_
timestamp 1698431365
transform 1 0 43344 0 -1 37632
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1953_
timestamp 1698431365
transform 1 0 41104 0 1 17248
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1954_
timestamp 1698431365
transform 1 0 41664 0 -1 15680
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1955_
timestamp 1698431365
transform 1 0 45136 0 1 15680
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1956_
timestamp 1698431365
transform 1 0 45136 0 -1 18816
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1957_
timestamp 1698431365
transform 1 0 45136 0 1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1958_
timestamp 1698431365
transform 1 0 45136 0 -1 23520
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1959_
timestamp 1698431365
transform 1 0 45136 0 -1 26656
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1960_
timestamp 1698431365
transform 1 0 23296 0 1 23520
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1961_
timestamp 1698431365
transform 1 0 26768 0 -1 28224
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1962_
timestamp 1698431365
transform 1 0 45136 0 -1 29792
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1963_
timestamp 1698431365
transform -1 0 45584 0 -1 31360
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1964_
timestamp 1698431365
transform 1 0 43008 0 -1 34496
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1965_
timestamp 1698431365
transform 1 0 45136 0 1 32928
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1966_
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1967_
timestamp 1698431365
transform 1 0 45136 0 1 12544
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1968_
timestamp 1698431365
transform 1 0 45136 0 1 9408
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1969_
timestamp 1698431365
transform 1 0 42112 0 -1 10976
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1970_
timestamp 1698431365
transform 1 0 41104 0 1 12544
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1971_
timestamp 1698431365
transform 1 0 44464 0 -1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1972_
timestamp 1698431365
transform 1 0 39648 0 1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1973_
timestamp 1698431365
transform 1 0 42000 0 -1 25088
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1974_
timestamp 1698431365
transform 1 0 41776 0 -1 29792
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1975_
timestamp 1698431365
transform -1 0 39536 0 -1 31360
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1976_
timestamp 1698431365
transform -1 0 38640 0 -1 32928
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1977_
timestamp 1698431365
transform -1 0 41440 0 1 34496
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1978_
timestamp 1698431365
transform 1 0 34272 0 -1 36064
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1979_
timestamp 1698431365
transform 1 0 19152 0 -1 42336
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1980_
timestamp 1698431365
transform 1 0 18928 0 -1 43904
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1981_
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1982_
timestamp 1698431365
transform 1 0 20048 0 -1 39200
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1983_
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1984_
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1985_
timestamp 1698431365
transform 1 0 13664 0 -1 23520
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1986_
timestamp 1698431365
transform 1 0 13440 0 1 26656
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1987_
timestamp 1698431365
transform 1 0 10640 0 -1 28224
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1988_
timestamp 1698431365
transform 1 0 12880 0 -1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1989_
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1990_
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1991_
timestamp 1698431365
transform 1 0 5712 0 -1 31360
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1992_
timestamp 1698431365
transform 1 0 5824 0 1 32928
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1993_
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1994_
timestamp 1698431365
transform 1 0 2352 0 -1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1995_
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1996_
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1997_
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1998_
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1999_
timestamp 1698431365
transform 1 0 1680 0 1 28224
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2000_
timestamp 1698431365
transform 1 0 5824 0 -1 28224
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2001_
timestamp 1698431365
transform -1 0 8848 0 1 26656
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2002_
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2003_
timestamp 1698431365
transform 1 0 1792 0 -1 25088
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2004_
timestamp 1698431365
transform 1 0 6496 0 1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2005_
timestamp 1698431365
transform -1 0 8736 0 -1 25088
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2006_
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2007_
timestamp 1698431365
transform 1 0 1680 0 -1 21952
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2008_
timestamp 1698431365
transform 1 0 5824 0 -1 20384
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2009_
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2010_
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2011_
timestamp 1698431365
transform 1 0 5824 0 -1 17248
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2012_
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2013_
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2014_
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2015_
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2016_
timestamp 1698431365
transform 1 0 1680 0 -1 4704
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2017_
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2018_
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2019_
timestamp 1698431365
transform 1 0 7840 0 1 14112
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2020_
timestamp 1698431365
transform 1 0 7840 0 1 10976
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2021_
timestamp 1698431365
transform 1 0 5040 0 -1 10976
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2022_
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2023_
timestamp 1698431365
transform 1 0 5488 0 -1 6272
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2024_
timestamp 1698431365
transform 1 0 33936 0 -1 6272
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2025_
timestamp 1698431365
transform 1 0 36400 0 -1 4704
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2026_
timestamp 1698431365
transform -1 0 44128 0 -1 4704
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2027_
timestamp 1698431365
transform 1 0 40544 0 1 6272
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2028_
timestamp 1698431365
transform 1 0 44128 0 -1 4704
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2029_
timestamp 1698431365
transform 1 0 45136 0 1 7840
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2030_
timestamp 1698431365
transform 1 0 45136 0 1 4704
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2031_
timestamp 1698431365
transform 1 0 8848 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2032_
timestamp 1698431365
transform 1 0 5936 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2033_
timestamp 1698431365
transform 1 0 21616 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2034_
timestamp 1698431365
transform 1 0 15344 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2035_
timestamp 1698431365
transform -1 0 32704 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2036_
timestamp 1698431365
transform -1 0 34832 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2037_
timestamp 1698431365
transform 1 0 10864 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2038_
timestamp 1698431365
transform 1 0 19600 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2039_
timestamp 1698431365
transform 1 0 32032 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2040_
timestamp 1698431365
transform -1 0 39200 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2041_
timestamp 1698431365
transform -1 0 40096 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2042_
timestamp 1698431365
transform 1 0 32928 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2043_
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2044_
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2045_
timestamp 1698431365
transform -1 0 42224 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2046_
timestamp 1698431365
transform -1 0 42112 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2047_
timestamp 1698431365
transform -1 0 38528 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2048_
timestamp 1698431365
transform -1 0 41104 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2059_
timestamp 1698431365
transform 1 0 42000 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__A1 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__I
timestamp 1698431365
transform 1 0 17024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0970__I
timestamp 1698431365
transform -1 0 31024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__A1
timestamp 1698431365
transform 1 0 21504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__A2
timestamp 1698431365
transform -1 0 22176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__A2
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__B
timestamp 1698431365
transform -1 0 25872 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__I
timestamp 1698431365
transform 1 0 35504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__A2
timestamp 1698431365
transform 1 0 39536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A1
timestamp 1698431365
transform 1 0 37856 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A2
timestamp 1698431365
transform -1 0 37968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1024__A1
timestamp 1698431365
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__A1
timestamp 1698431365
transform 1 0 36064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__A2
timestamp 1698431365
transform -1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A1
timestamp 1698431365
transform 1 0 35056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1029__A2
timestamp 1698431365
transform 1 0 19824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__A2
timestamp 1698431365
transform 1 0 20832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__B
timestamp 1698431365
transform 1 0 39984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1033__A2
timestamp 1698431365
transform -1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A2
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__I
timestamp 1698431365
transform 1 0 22400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__I
timestamp 1698431365
transform -1 0 14448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__I
timestamp 1698431365
transform 1 0 24528 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__B1
timestamp 1698431365
transform 1 0 28224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A1
timestamp 1698431365
transform 1 0 28224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A2
timestamp 1698431365
transform 1 0 27776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A3
timestamp 1698431365
transform -1 0 27776 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__A1
timestamp 1698431365
transform 1 0 25424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__A1
timestamp 1698431365
transform 1 0 37296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__B
timestamp 1698431365
transform 1 0 35952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A2
timestamp 1698431365
transform 1 0 30128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__I
timestamp 1698431365
transform 1 0 34944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__I
timestamp 1698431365
transform -1 0 10640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__I
timestamp 1698431365
transform -1 0 31024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A1
timestamp 1698431365
transform -1 0 31360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A2
timestamp 1698431365
transform 1 0 32704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A1
timestamp 1698431365
transform -1 0 33824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A2
timestamp 1698431365
transform 1 0 30464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__I
timestamp 1698431365
transform -1 0 12208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__I
timestamp 1698431365
transform 1 0 13104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1110__A1
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__I
timestamp 1698431365
transform -1 0 23856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A1
timestamp 1698431365
transform 1 0 22400 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__I
timestamp 1698431365
transform -1 0 14112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__A1
timestamp 1698431365
transform -1 0 22960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1128__I
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__I
timestamp 1698431365
transform -1 0 23968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__A3
timestamp 1698431365
transform 1 0 22064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__A1
timestamp 1698431365
transform 1 0 21392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__A1
timestamp 1698431365
transform 1 0 24080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__A2
timestamp 1698431365
transform -1 0 23856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1140__A1
timestamp 1698431365
transform 1 0 18816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__I
timestamp 1698431365
transform -1 0 30128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__S
timestamp 1698431365
transform 1 0 25424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__I
timestamp 1698431365
transform 1 0 25200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__I
timestamp 1698431365
transform 1 0 31584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1167__A1
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1169__A1
timestamp 1698431365
transform 1 0 24864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A1
timestamp 1698431365
transform 1 0 23520 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__C
timestamp 1698431365
transform -1 0 25200 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__A1
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__A2
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__A1
timestamp 1698431365
transform 1 0 21280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__A1
timestamp 1698431365
transform -1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1178__A2
timestamp 1698431365
transform 1 0 19712 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1178__B
timestamp 1698431365
transform -1 0 20384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1179__A2
timestamp 1698431365
transform 1 0 18480 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1180__A1
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1184__I
timestamp 1698431365
transform -1 0 13776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__A1
timestamp 1698431365
transform -1 0 24752 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1186__I
timestamp 1698431365
transform -1 0 14784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__C
timestamp 1698431365
transform 1 0 24080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1189__A2
timestamp 1698431365
transform 1 0 26768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__A2
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__A1
timestamp 1698431365
transform 1 0 26432 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A1
timestamp 1698431365
transform 1 0 25424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1194__C
timestamp 1698431365
transform 1 0 26992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1196__I
timestamp 1698431365
transform -1 0 36064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__A1
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__B
timestamp 1698431365
transform 1 0 30912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__B
timestamp 1698431365
transform 1 0 28224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1203__B
timestamp 1698431365
transform 1 0 26992 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__A1
timestamp 1698431365
transform 1 0 32032 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__I
timestamp 1698431365
transform -1 0 34048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1209__A2
timestamp 1698431365
transform -1 0 28224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__A2
timestamp 1698431365
transform 1 0 29680 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__A1
timestamp 1698431365
transform 1 0 31584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__A1
timestamp 1698431365
transform 1 0 34496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__B
timestamp 1698431365
transform -1 0 31808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__I
timestamp 1698431365
transform 1 0 41216 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__C
timestamp 1698431365
transform 1 0 39424 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__I
timestamp 1698431365
transform 1 0 38304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__S
timestamp 1698431365
transform 1 0 45360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__B
timestamp 1698431365
transform -1 0 39984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__I
timestamp 1698431365
transform 1 0 13552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1228__C
timestamp 1698431365
transform 1 0 44016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__I
timestamp 1698431365
transform -1 0 41328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1231__I0
timestamp 1698431365
transform 1 0 43232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1234__C
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__B
timestamp 1698431365
transform -1 0 31696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__C
timestamp 1698431365
transform 1 0 31472 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1237__B
timestamp 1698431365
transform 1 0 27888 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__S
timestamp 1698431365
transform 1 0 19152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1240__I
timestamp 1698431365
transform 1 0 44128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__A1
timestamp 1698431365
transform -1 0 19376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__A1
timestamp 1698431365
transform -1 0 20720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__A1
timestamp 1698431365
transform 1 0 19936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__C
timestamp 1698431365
transform 1 0 20608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1248__A1
timestamp 1698431365
transform -1 0 18144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1250__A2
timestamp 1698431365
transform -1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1250__B
timestamp 1698431365
transform -1 0 20496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1251__A2
timestamp 1698431365
transform 1 0 18144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1252__A1
timestamp 1698431365
transform 1 0 25312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__I
timestamp 1698431365
transform 1 0 15344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1256__A1
timestamp 1698431365
transform -1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__A1
timestamp 1698431365
transform -1 0 9968 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__A2
timestamp 1698431365
transform -1 0 11424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1259__A2
timestamp 1698431365
transform -1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__A1
timestamp 1698431365
transform -1 0 14224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__A1
timestamp 1698431365
transform 1 0 14000 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A1
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__C
timestamp 1698431365
transform -1 0 11760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__S
timestamp 1698431365
transform -1 0 10192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__A1
timestamp 1698431365
transform 1 0 15008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__B
timestamp 1698431365
transform -1 0 15568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1266__B
timestamp 1698431365
transform -1 0 13776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__B
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1269__A2
timestamp 1698431365
transform -1 0 22960 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__A1
timestamp 1698431365
transform -1 0 23856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__C
timestamp 1698431365
transform 1 0 24080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A1
timestamp 1698431365
transform 1 0 16240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A2
timestamp 1698431365
transform -1 0 19824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__A2
timestamp 1698431365
transform -1 0 21056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A1
timestamp 1698431365
transform 1 0 23184 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1276__A1
timestamp 1698431365
transform 1 0 30800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__A1
timestamp 1698431365
transform 1 0 28672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__B
timestamp 1698431365
transform 1 0 31360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1281__A1
timestamp 1698431365
transform -1 0 39424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__A2
timestamp 1698431365
transform 1 0 40992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__C
timestamp 1698431365
transform 1 0 40320 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1288__B
timestamp 1698431365
transform 1 0 43008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1289__C
timestamp 1698431365
transform -1 0 39984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__C
timestamp 1698431365
transform -1 0 29456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__I3
timestamp 1698431365
transform -1 0 36736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__S0
timestamp 1698431365
transform 1 0 40544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__S1
timestamp 1698431365
transform -1 0 37296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A1
timestamp 1698431365
transform 1 0 39200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__S0
timestamp 1698431365
transform 1 0 45472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__S1
timestamp 1698431365
transform 1 0 42448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1298__A1
timestamp 1698431365
transform -1 0 34720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1301__I
timestamp 1698431365
transform -1 0 9072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1303__I
timestamp 1698431365
transform 1 0 13104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1304__A1
timestamp 1698431365
transform -1 0 9072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1306__A2
timestamp 1698431365
transform -1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1306__C
timestamp 1698431365
transform 1 0 14000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__A1
timestamp 1698431365
transform 1 0 10192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1309__A2
timestamp 1698431365
transform -1 0 10976 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1309__C
timestamp 1698431365
transform -1 0 11424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1311__C
timestamp 1698431365
transform -1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1312__A1
timestamp 1698431365
transform -1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1313__A1
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1314__A2
timestamp 1698431365
transform -1 0 13552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1314__C
timestamp 1698431365
transform -1 0 11200 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1316__A1
timestamp 1698431365
transform 1 0 11536 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__A1
timestamp 1698431365
transform 1 0 8400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__A2
timestamp 1698431365
transform -1 0 14448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__B1
timestamp 1698431365
transform 1 0 14672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__B2
timestamp 1698431365
transform -1 0 8176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__C
timestamp 1698431365
transform -1 0 14000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__C
timestamp 1698431365
transform -1 0 13104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1319__A1
timestamp 1698431365
transform 1 0 15680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__A1
timestamp 1698431365
transform 1 0 9744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1321__A1
timestamp 1698431365
transform 1 0 10640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__B
timestamp 1698431365
transform 1 0 11984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1325__A2
timestamp 1698431365
transform -1 0 10528 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1326__A2
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1326__C
timestamp 1698431365
transform 1 0 12432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1327__A1
timestamp 1698431365
transform -1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__A1
timestamp 1698431365
transform -1 0 10752 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1329__B
timestamp 1698431365
transform 1 0 11648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__A2
timestamp 1698431365
transform 1 0 10416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1332__A2
timestamp 1698431365
transform 1 0 11088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1332__C
timestamp 1698431365
transform 1 0 10864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1333__C
timestamp 1698431365
transform 1 0 12544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1336__A1
timestamp 1698431365
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1336__A2
timestamp 1698431365
transform -1 0 10304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A2
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A1
timestamp 1698431365
transform -1 0 11872 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1340__C
timestamp 1698431365
transform -1 0 10416 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1341__S
timestamp 1698431365
transform 1 0 5712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__B
timestamp 1698431365
transform -1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__B
timestamp 1698431365
transform -1 0 12208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1344__B
timestamp 1698431365
transform 1 0 14224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__B
timestamp 1698431365
transform 1 0 17584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__S
timestamp 1698431365
transform 1 0 15344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__A2
timestamp 1698431365
transform 1 0 14784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__A2
timestamp 1698431365
transform 1 0 14896 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A1
timestamp 1698431365
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1352__A1
timestamp 1698431365
transform 1 0 18592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__A2
timestamp 1698431365
transform -1 0 20832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__B
timestamp 1698431365
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1355__A2
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__A1
timestamp 1698431365
transform 1 0 19264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A1
timestamp 1698431365
transform 1 0 21616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__C
timestamp 1698431365
transform 1 0 25424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__A2
timestamp 1698431365
transform -1 0 24304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__A2
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1361__A1
timestamp 1698431365
transform -1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__A2
timestamp 1698431365
transform 1 0 27440 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A1
timestamp 1698431365
transform 1 0 29232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__C
timestamp 1698431365
transform 1 0 26096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1365__B
timestamp 1698431365
transform 1 0 29344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__B
timestamp 1698431365
transform 1 0 27552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1367__B
timestamp 1698431365
transform 1 0 25648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1369__A1
timestamp 1698431365
transform 1 0 39424 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A2
timestamp 1698431365
transform 1 0 38528 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__A1
timestamp 1698431365
transform -1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__A2
timestamp 1698431365
transform 1 0 27776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__B
timestamp 1698431365
transform -1 0 28896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__A2
timestamp 1698431365
transform 1 0 28224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1373__A1
timestamp 1698431365
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1373__A2
timestamp 1698431365
transform 1 0 34496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__B
timestamp 1698431365
transform -1 0 32480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__C
timestamp 1698431365
transform -1 0 45136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1380__S
timestamp 1698431365
transform -1 0 45248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1382__A1
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1383__C
timestamp 1698431365
transform 1 0 39648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1384__S
timestamp 1698431365
transform -1 0 42784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__B
timestamp 1698431365
transform 1 0 38864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__C
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__C
timestamp 1698431365
transform 1 0 27776 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A2
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__C
timestamp 1698431365
transform 1 0 26096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__A2
timestamp 1698431365
transform 1 0 23184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__A3
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1405__A2
timestamp 1698431365
transform 1 0 27104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1405__B
timestamp 1698431365
transform -1 0 27552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__1_I
timestamp 1698431365
transform 1 0 36400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1416__I
timestamp 1698431365
transform -1 0 14560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__I
timestamp 1698431365
transform 1 0 16016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__A1
timestamp 1698431365
transform 1 0 27776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1422__A1
timestamp 1698431365
transform 1 0 26992 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A1
timestamp 1698431365
transform -1 0 25984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1424__A1
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1424__A3
timestamp 1698431365
transform -1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__I
timestamp 1698431365
transform -1 0 20496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A1
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__I
timestamp 1698431365
transform -1 0 23744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__A2
timestamp 1698431365
transform 1 0 24192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__C
timestamp 1698431365
transform -1 0 15120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__B
timestamp 1698431365
transform 1 0 15792 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1499__A1
timestamp 1698431365
transform 1 0 13888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1499__A2
timestamp 1698431365
transform -1 0 15680 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__I1
timestamp 1698431365
transform 1 0 9632 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__I
timestamp 1698431365
transform 1 0 17584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__I
timestamp 1698431365
transform 1 0 17696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__I
timestamp 1698431365
transform 1 0 18592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__I0
timestamp 1698431365
transform 1 0 22624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__I
timestamp 1698431365
transform -1 0 27440 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1560__I1
timestamp 1698431365
transform 1 0 26880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__I0
timestamp 1698431365
transform 1 0 40320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__I1
timestamp 1698431365
transform 1 0 40208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__I
timestamp 1698431365
transform 1 0 27664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__I
timestamp 1698431365
transform 1 0 20384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__I0
timestamp 1698431365
transform 1 0 44912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__I
timestamp 1698431365
transform 1 0 47712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I1
timestamp 1698431365
transform -1 0 45136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__I
timestamp 1698431365
transform 1 0 47152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I0
timestamp 1698431365
transform 1 0 48272 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1698431365
transform -1 0 24304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A1
timestamp 1698431365
transform 1 0 27328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__I1
timestamp 1698431365
transform 1 0 45472 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__I
timestamp 1698431365
transform -1 0 45696 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__I0
timestamp 1698431365
transform 1 0 48272 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__I
timestamp 1698431365
transform -1 0 46704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__I1
timestamp 1698431365
transform 1 0 48272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__I
timestamp 1698431365
transform 1 0 38752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__I
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__I0
timestamp 1698431365
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__I
timestamp 1698431365
transform -1 0 21840 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__I1
timestamp 1698431365
transform 1 0 23072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A2
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__I
timestamp 1698431365
transform 1 0 18816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A2
timestamp 1698431365
transform 1 0 13552 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__I
timestamp 1698431365
transform 1 0 6720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__I
timestamp 1698431365
transform 1 0 6160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A2
timestamp 1698431365
transform 1 0 9968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__I
timestamp 1698431365
transform 1 0 6944 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__A2
timestamp 1698431365
transform -1 0 7840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__I
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__I
timestamp 1698431365
transform 1 0 6048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__I0
timestamp 1698431365
transform 1 0 5152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__I0
timestamp 1698431365
transform -1 0 3136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__I1
timestamp 1698431365
transform 1 0 4256 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__I
timestamp 1698431365
transform 1 0 6720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__I1
timestamp 1698431365
transform 1 0 5264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__I
timestamp 1698431365
transform 1 0 35728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__S
timestamp 1698431365
transform -1 0 9520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__S
timestamp 1698431365
transform 1 0 9632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__I0
timestamp 1698431365
transform -1 0 8288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__S
timestamp 1698431365
transform -1 0 7840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__I1
timestamp 1698431365
transform -1 0 35616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__S
timestamp 1698431365
transform 1 0 37520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__I
timestamp 1698431365
transform 1 0 38192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__S
timestamp 1698431365
transform 1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__S
timestamp 1698431365
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__A1
timestamp 1698431365
transform -1 0 33376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__A3
timestamp 1698431365
transform 1 0 35056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A1
timestamp 1698431365
transform 1 0 34048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__A1
timestamp 1698431365
transform 1 0 31248 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A3
timestamp 1698431365
transform 1 0 33152 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A1
timestamp 1698431365
transform 1 0 34832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A2
timestamp 1698431365
transform 1 0 34048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A1
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__A1
timestamp 1698431365
transform 1 0 28448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__C
timestamp 1698431365
transform 1 0 27552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__S
timestamp 1698431365
transform -1 0 11984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A1
timestamp 1698431365
transform -1 0 12432 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__A1
timestamp 1698431365
transform -1 0 11088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A1
timestamp 1698431365
transform 1 0 33600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__A1
timestamp 1698431365
transform 1 0 35056 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__A1
timestamp 1698431365
transform -1 0 15008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__I
timestamp 1698431365
transform 1 0 38192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A1
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A2
timestamp 1698431365
transform -1 0 34048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__A2
timestamp 1698431365
transform 1 0 38416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A2
timestamp 1698431365
transform 1 0 37968 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__A2
timestamp 1698431365
transform -1 0 32256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__I
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A1
timestamp 1698431365
transform 1 0 42336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__I
timestamp 1698431365
transform -1 0 37968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__CLK
timestamp 1698431365
transform 1 0 5712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__CLK
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__CLK
timestamp 1698431365
transform 1 0 23520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__CLK
timestamp 1698431365
transform 1 0 23744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__CLK
timestamp 1698431365
transform 1 0 22176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__CLK
timestamp 1698431365
transform 1 0 14336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__CLK
timestamp 1698431365
transform -1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__CLK
timestamp 1698431365
transform 1 0 14896 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__CLK
timestamp 1698431365
transform 1 0 35840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__CLK
timestamp 1698431365
transform 1 0 24528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__CLK
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__CLKN
timestamp 1698431365
transform 1 0 9632 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__CLKN
timestamp 1698431365
transform 1 0 12880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__CLKN
timestamp 1698431365
transform 1 0 9184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__CLKN
timestamp 1698431365
transform 1 0 8848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__CLKN
timestamp 1698431365
transform 1 0 10864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__CLKN
timestamp 1698431365
transform 1 0 11648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__CLKN
timestamp 1698431365
transform 1 0 13552 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__CLKN
timestamp 1698431365
transform 1 0 10752 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__CLKN
timestamp 1698431365
transform 1 0 17136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__CLKN
timestamp 1698431365
transform 1 0 18144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__CLKN
timestamp 1698431365
transform 1 0 18816 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__CLKN
timestamp 1698431365
transform 1 0 11536 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__CLKN
timestamp 1698431365
transform 1 0 12880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__CLKN
timestamp 1698431365
transform 1 0 16240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__CLKN
timestamp 1698431365
transform 1 0 19600 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__CLKN
timestamp 1698431365
transform 1 0 19600 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__CLKN
timestamp 1698431365
transform 1 0 17584 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__CLKN
timestamp 1698431365
transform -1 0 21168 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__CLKN
timestamp 1698431365
transform -1 0 21616 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__CLKN
timestamp 1698431365
transform 1 0 30128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__CLKN
timestamp 1698431365
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__CLKN
timestamp 1698431365
transform 1 0 33824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__CLKN
timestamp 1698431365
transform 1 0 33376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__CLKN
timestamp 1698431365
transform 1 0 40208 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__CLKN
timestamp 1698431365
transform 1 0 39424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__CLKN
timestamp 1698431365
transform 1 0 40432 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__CLKN
timestamp 1698431365
transform 1 0 41104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__CLKN
timestamp 1698431365
transform 1 0 38416 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__CLKN
timestamp 1698431365
transform 1 0 41664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__CLKN
timestamp 1698431365
transform 1 0 42336 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__CLKN
timestamp 1698431365
transform 1 0 41776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__CLKN
timestamp 1698431365
transform 1 0 35952 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__CLKN
timestamp 1698431365
transform 1 0 36176 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1929__CLKN
timestamp 1698431365
transform 1 0 32368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__CLKN
timestamp 1698431365
transform -1 0 29008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__CLKN
timestamp 1698431365
transform 1 0 22960 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__CLKN
timestamp 1698431365
transform 1 0 23072 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__CLKN
timestamp 1698431365
transform 1 0 23520 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__CLKN
timestamp 1698431365
transform 1 0 22960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__CLKN
timestamp 1698431365
transform -1 0 20272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1936__CLKN
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__CLKN
timestamp 1698431365
transform 1 0 22400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1939__CLKN
timestamp 1698431365
transform 1 0 23632 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__CLKN
timestamp 1698431365
transform 1 0 21056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__CLKN
timestamp 1698431365
transform 1 0 24080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__CLKN
timestamp 1698431365
transform 1 0 29568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__CLKN
timestamp 1698431365
transform 1 0 30464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__CLKN
timestamp 1698431365
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__CLKN
timestamp 1698431365
transform 1 0 34272 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__CLKN
timestamp 1698431365
transform 1 0 36288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__CLKN
timestamp 1698431365
transform 1 0 40992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__CLKN
timestamp 1698431365
transform 1 0 39984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__CLKN
timestamp 1698431365
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__CLKN
timestamp 1698431365
transform 1 0 40320 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__CLKN
timestamp 1698431365
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__CLKN
timestamp 1698431365
transform 1 0 41888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1954__CLKN
timestamp 1698431365
transform 1 0 45360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__CLKN
timestamp 1698431365
transform 1 0 44912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1956__CLKN
timestamp 1698431365
transform 1 0 44688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__CLKN
timestamp 1698431365
transform 1 0 45360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1958__CLKN
timestamp 1698431365
transform 1 0 44912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__CLKN
timestamp 1698431365
transform 1 0 44912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__CLKN
timestamp 1698431365
transform 1 0 31920 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1967__CLKN
timestamp 1698431365
transform 1 0 44912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__CLKN
timestamp 1698431365
transform 1 0 44912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__CLKN
timestamp 1698431365
transform 1 0 45472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__CLKN
timestamp 1698431365
transform 1 0 40992 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__CLKN
timestamp 1698431365
transform 1 0 44912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__CLKN
timestamp 1698431365
transform 1 0 43232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__CLKN
timestamp 1698431365
transform 1 0 45584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__CLKN
timestamp 1698431365
transform -1 0 35168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1979__CLKN
timestamp 1698431365
transform 1 0 18928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__CLKN
timestamp 1698431365
transform 1 0 18704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__CLKN
timestamp 1698431365
transform 1 0 20944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__CLKN
timestamp 1698431365
transform -1 0 23632 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__CLKN
timestamp 1698431365
transform 1 0 14672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__CLKN
timestamp 1698431365
transform 1 0 5152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__CLKN
timestamp 1698431365
transform 1 0 5712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__CLKN
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__CLKN
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__CLKN
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__CLKN
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__CLKN
timestamp 1698431365
transform 1 0 9296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__CLKN
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__CLKN
timestamp 1698431365
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__CLKN
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__CLKN
timestamp 1698431365
transform 1 0 8400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__CLKN
timestamp 1698431365
transform 1 0 5712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__CLKN
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__CLKN
timestamp 1698431365
transform 1 0 9632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__CLKN
timestamp 1698431365
transform 1 0 5040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__CLKN
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__CLKN
timestamp 1698431365
transform 1 0 5040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__CLKN
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__CLKN
timestamp 1698431365
transform 1 0 1792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__CLKN
timestamp 1698431365
transform 1 0 5712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__CLKN
timestamp 1698431365
transform 1 0 6944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__CLKN
timestamp 1698431365
transform -1 0 11648 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__CLKN
timestamp 1698431365
transform 1 0 11424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__CLKN
timestamp 1698431365
transform 1 0 8624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__CLKN
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__CLKN
timestamp 1698431365
transform 1 0 7168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__CLKN
timestamp 1698431365
transform 1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__CLKN
timestamp 1698431365
transform 1 0 39760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__CLKN
timestamp 1698431365
transform 1 0 40992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2027__CLKN
timestamp 1698431365
transform 1 0 40320 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__CLKN
timestamp 1698431365
transform 1 0 43232 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__CLKN
timestamp 1698431365
transform 1 0 44912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__CLKN
timestamp 1698431365
transform 1 0 44912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__CLK
timestamp 1698431365
transform 1 0 11312 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__CLK
timestamp 1698431365
transform 1 0 6048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2033__CLK
timestamp 1698431365
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2034__CLK
timestamp 1698431365
transform 1 0 14336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__CLK
timestamp 1698431365
transform 1 0 35504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__CLK
timestamp 1698431365
transform 1 0 35952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__CLK
timestamp 1698431365
transform 1 0 9744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__CLK
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__CLK
timestamp 1698431365
transform 1 0 35504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__CLK
timestamp 1698431365
transform -1 0 39648 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__CLK
timestamp 1698431365
transform 1 0 40320 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__CLK
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__CLK
timestamp 1698431365
transform 1 0 41664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__CLK
timestamp 1698431365
transform 1 0 41664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__CLK
timestamp 1698431365
transform 1 0 38752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__CLK
timestamp 1698431365
transform 1 0 42336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__CLK
timestamp 1698431365
transform 1 0 38528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__CLK
timestamp 1698431365
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__I
timestamp 1698431365
transform -1 0 42224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 25200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_clk_I
timestamp 1698431365
transform 1 0 15120 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_clk_I
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_clk_I
timestamp 1698431365
transform 1 0 20384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_clk_I
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_clk_I
timestamp 1698431365
transform 1 0 14224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_clk_I
timestamp 1698431365
transform 1 0 15792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_clk_I
timestamp 1698431365
transform 1 0 21280 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_clk_I
timestamp 1698431365
transform -1 0 18816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_clk_I
timestamp 1698431365
transform -1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_clk_I
timestamp 1698431365
transform 1 0 38528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_clk_I
timestamp 1698431365
transform 1 0 38976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_clk_I
timestamp 1698431365
transform 1 0 43568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_clk_I
timestamp 1698431365
transform 1 0 31136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_clk_I
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_clk_I
timestamp 1698431365
transform 1 0 39648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_clk_I
timestamp 1698431365
transform 1 0 37408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold1_I
timestamp 1698431365
transform -1 0 13552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold5_I
timestamp 1698431365
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold13_I
timestamp 1698431365
transform 1 0 21392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold14_I
timestamp 1698431365
transform -1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold15_I
timestamp 1698431365
transform -1 0 13776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 2016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 3584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 6496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 3360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 2912 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output12_I
timestamp 1698431365
transform 1 0 45360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output14_I
timestamp 1698431365
transform 1 0 38976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output17_I
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_clk asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13552 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1698431365
transform -1 0 13104 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1698431365
transform 1 0 17472 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1698431365
transform -1 0 13552 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1698431365
transform -1 0 14112 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1698431365
transform 1 0 18368 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1698431365
transform -1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1698431365
transform -1 0 39760 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1698431365
transform -1 0 40880 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1698431365
transform -1 0 43344 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1698431365
transform -1 0 43680 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1698431365
transform 1 0 31360 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1698431365
transform 1 0 38864 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1698431365
transform -1 0 40544 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_46 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_106 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13216 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_134
timestamp 1698431365
transform 1 0 16352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_163
timestamp 1698431365
transform 1 0 19600 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_338
timestamp 1698431365
transform 1 0 39200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_372
timestamp 1698431365
transform 1 0 43008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_406
timestamp 1698431365
transform 1 0 46816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_414
timestamp 1698431365
transform 1 0 47712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_416
timestamp 1698431365
transform 1 0 47936 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_33
timestamp 1698431365
transform 1 0 5040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_74
timestamp 1698431365
transform 1 0 9632 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_155
timestamp 1698431365
transform 1 0 18704 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_180
timestamp 1698431365
transform 1 0 21504 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_310
timestamp 1698431365
transform 1 0 36064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_312
timestamp 1698431365
transform 1 0 36288 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_343
timestamp 1698431365
transform 1 0 39760 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_412 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47488 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_420
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_12
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_16
timestamp 1698431365
transform 1 0 3136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_94
timestamp 1698431365
transform 1 0 11872 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_96
timestamp 1698431365
transform 1 0 12096 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_170
timestamp 1698431365
transform 1 0 20384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_172
timestamp 1698431365
transform 1 0 20608 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_299
timestamp 1698431365
transform 1 0 34832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_303
timestamp 1698431365
transform 1 0 35280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_307
timestamp 1698431365
transform 1 0 35728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_321
timestamp 1698431365
transform 1 0 37296 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_369 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42672 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_373
timestamp 1698431365
transform 1 0 43120 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_382
timestamp 1698431365
transform 1 0 44128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_384
timestamp 1698431365
transform 1 0 44352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_32
timestamp 1698431365
transform 1 0 4928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_36
timestamp 1698431365
transform 1 0 5376 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_67
timestamp 1698431365
transform 1 0 8848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_114
timestamp 1698431365
transform 1 0 14112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_200
timestamp 1698431365
transform 1 0 23744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_233
timestamp 1698431365
transform 1 0 27440 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_235
timestamp 1698431365
transform 1 0 27664 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_284
timestamp 1698431365
transform 1 0 33152 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_327
timestamp 1698431365
transform 1 0 37968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_331
timestamp 1698431365
transform 1 0 38416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_356
timestamp 1698431365
transform 1 0 41216 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_361
timestamp 1698431365
transform 1 0 41776 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_365
timestamp 1698431365
transform 1 0 42224 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_384
timestamp 1698431365
transform 1 0 44352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_388
timestamp 1698431365
transform 1 0 44800 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_391
timestamp 1698431365
transform 1 0 45136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_6
timestamp 1698431365
transform 1 0 2016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_10
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_14
timestamp 1698431365
transform 1 0 2912 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_33
timestamp 1698431365
transform 1 0 5040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_41
timestamp 1698431365
transform 1 0 5936 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_50
timestamp 1698431365
transform 1 0 6944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_52
timestamp 1698431365
transform 1 0 7168 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_68
timestamp 1698431365
transform 1 0 8960 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_130
timestamp 1698431365
transform 1 0 15904 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_147
timestamp 1698431365
transform 1 0 17808 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_192
timestamp 1698431365
transform 1 0 22848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_194
timestamp 1698431365
transform 1 0 23072 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_197
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_217
timestamp 1698431365
transform 1 0 25648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_232
timestamp 1698431365
transform 1 0 27328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_234
timestamp 1698431365
transform 1 0 27552 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_243
timestamp 1698431365
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_265
timestamp 1698431365
transform 1 0 31024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_269
timestamp 1698431365
transform 1 0 31472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_321
timestamp 1698431365
transform 1 0 37296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_325
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_334
timestamp 1698431365
transform 1 0 38752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_338
timestamp 1698431365
transform 1 0 39200 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_342
timestamp 1698431365
transform 1 0 39648 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_345
timestamp 1698431365
transform 1 0 39984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_347
timestamp 1698431365
transform 1 0 40208 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_380
timestamp 1698431365
transform 1 0 43904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_384
timestamp 1698431365
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_389
timestamp 1698431365
transform 1 0 44912 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_392
timestamp 1698431365
transform 1 0 45248 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_417
timestamp 1698431365
transform 1 0 48048 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_12
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_20
timestamp 1698431365
transform 1 0 3584 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_24
timestamp 1698431365
transform 1 0 4032 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_28
timestamp 1698431365
transform 1 0 4480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_40
timestamp 1698431365
transform 1 0 5824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_44
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_48
timestamp 1698431365
transform 1 0 6720 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_54
timestamp 1698431365
transform 1 0 7392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_58
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_62
timestamp 1698431365
transform 1 0 8288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_74
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_83
timestamp 1698431365
transform 1 0 10640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_85
timestamp 1698431365
transform 1 0 10864 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_106
timestamp 1698431365
transform 1 0 13216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_114
timestamp 1698431365
transform 1 0 14112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_116
timestamp 1698431365
transform 1 0 14336 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_166
timestamp 1698431365
transform 1 0 19936 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_196
timestamp 1698431365
transform 1 0 23296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_200
timestamp 1698431365
transform 1 0 23744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_202
timestamp 1698431365
transform 1 0 23968 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_205
timestamp 1698431365
transform 1 0 24304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_230
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_234
timestamp 1698431365
transform 1 0 27552 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_243
timestamp 1698431365
transform 1 0 28560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_272
timestamp 1698431365
transform 1 0 31808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_286
timestamp 1698431365
transform 1 0 33376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_290
timestamp 1698431365
transform 1 0 33824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_294
timestamp 1698431365
transform 1 0 34272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_298
timestamp 1698431365
transform 1 0 34720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_302
timestamp 1698431365
transform 1 0 35168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_306
timestamp 1698431365
transform 1 0 35616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_310
timestamp 1698431365
transform 1 0 36064 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_316
timestamp 1698431365
transform 1 0 36736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_420
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_96
timestamp 1698431365
transform 1 0 12096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_98
timestamp 1698431365
transform 1 0 12320 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_120
timestamp 1698431365
transform 1 0 14784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_122
timestamp 1698431365
transform 1 0 15008 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_129
timestamp 1698431365
transform 1 0 15792 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_137
timestamp 1698431365
transform 1 0 16688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_158
timestamp 1698431365
transform 1 0 19040 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_165
timestamp 1698431365
transform 1 0 19824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_173
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_206
timestamp 1698431365
transform 1 0 24416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_208
timestamp 1698431365
transform 1 0 24640 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_240
timestamp 1698431365
transform 1 0 28224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_290
timestamp 1698431365
transform 1 0 33824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_294
timestamp 1698431365
transform 1 0 34272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_296
timestamp 1698431365
transform 1 0 34496 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_305
timestamp 1698431365
transform 1 0 35504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_309
timestamp 1698431365
transform 1 0 35952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_313
timestamp 1698431365
transform 1 0 36400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_323
timestamp 1698431365
transform 1 0 37520 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_327
timestamp 1698431365
transform 1 0 37968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_331
timestamp 1698431365
transform 1 0 38416 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_334 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38752 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_352
timestamp 1698431365
transform 1 0 40768 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_362
timestamp 1698431365
transform 1 0 41888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_366
timestamp 1698431365
transform 1 0 42336 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_369
timestamp 1698431365
transform 1 0 42672 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_10
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_14
timestamp 1698431365
transform 1 0 2912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_31
timestamp 1698431365
transform 1 0 4816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_35
timestamp 1698431365
transform 1 0 5264 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_49
timestamp 1698431365
transform 1 0 6832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_51
timestamp 1698431365
transform 1 0 7056 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_76
timestamp 1698431365
transform 1 0 9856 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_84
timestamp 1698431365
transform 1 0 10752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_87
timestamp 1698431365
transform 1 0 11088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_91
timestamp 1698431365
transform 1 0 11536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_107
timestamp 1698431365
transform 1 0 13328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_111
timestamp 1698431365
transform 1 0 13776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_115
timestamp 1698431365
transform 1 0 14224 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_184
timestamp 1698431365
transform 1 0 21952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_188
timestamp 1698431365
transform 1 0 22400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_198
timestamp 1698431365
transform 1 0 23520 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_219
timestamp 1698431365
transform 1 0 25872 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_227
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_229
timestamp 1698431365
transform 1 0 26992 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_232
timestamp 1698431365
transform 1 0 27328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_290
timestamp 1698431365
transform 1 0 33824 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_297
timestamp 1698431365
transform 1 0 34608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_301
timestamp 1698431365
transform 1 0 35056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_332
timestamp 1698431365
transform 1 0 38528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_342
timestamp 1698431365
transform 1 0 39648 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_352 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_384
timestamp 1698431365
transform 1 0 44352 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_392
timestamp 1698431365
transform 1 0 45248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_396
timestamp 1698431365
transform 1 0 45696 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_403
timestamp 1698431365
transform 1 0 46480 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_12
timestamp 1698431365
transform 1 0 2688 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_16
timestamp 1698431365
transform 1 0 3136 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_47
timestamp 1698431365
transform 1 0 6608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_51
timestamp 1698431365
transform 1 0 7056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_73
timestamp 1698431365
transform 1 0 9520 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_87
timestamp 1698431365
transform 1 0 11088 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_91
timestamp 1698431365
transform 1 0 11536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_95
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_99
timestamp 1698431365
transform 1 0 12432 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_103
timestamp 1698431365
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_111
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_118
timestamp 1698431365
transform 1 0 14560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_128
timestamp 1698431365
transform 1 0 15680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_130
timestamp 1698431365
transform 1 0 15904 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_133
timestamp 1698431365
transform 1 0 16240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_146
timestamp 1698431365
transform 1 0 17696 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_148
timestamp 1698431365
transform 1 0 17920 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_154
timestamp 1698431365
transform 1 0 18592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_158
timestamp 1698431365
transform 1 0 19040 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_163
timestamp 1698431365
transform 1 0 19600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_167
timestamp 1698431365
transform 1 0 20048 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_186
timestamp 1698431365
transform 1 0 22176 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_193
timestamp 1698431365
transform 1 0 22960 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_197
timestamp 1698431365
transform 1 0 23408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_199
timestamp 1698431365
transform 1 0 23632 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_231
timestamp 1698431365
transform 1 0 27216 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_255
timestamp 1698431365
transform 1 0 29904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_257
timestamp 1698431365
transform 1 0 30128 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_299
timestamp 1698431365
transform 1 0 34832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_312
timestamp 1698431365
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_333
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_335
timestamp 1698431365
transform 1 0 38864 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_365
timestamp 1698431365
transform 1 0 42224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_369
timestamp 1698431365
transform 1 0 42672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_371
timestamp 1698431365
transform 1 0 42896 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_378
timestamp 1698431365
transform 1 0 43680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_32
timestamp 1698431365
transform 1 0 4928 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_63
timestamp 1698431365
transform 1 0 8400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_67
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_116
timestamp 1698431365
transform 1 0 14336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_118
timestamp 1698431365
transform 1 0 14560 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_127
timestamp 1698431365
transform 1 0 15568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_131
timestamp 1698431365
transform 1 0 16016 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_144
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_151
timestamp 1698431365
transform 1 0 18256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_155
timestamp 1698431365
transform 1 0 18704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_180
timestamp 1698431365
transform 1 0 21504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_182
timestamp 1698431365
transform 1 0 21728 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_197
timestamp 1698431365
transform 1 0 23408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_205
timestamp 1698431365
transform 1 0 24304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_252
timestamp 1698431365
transform 1 0 29568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_319
timestamp 1698431365
transform 1 0 37072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_345
timestamp 1698431365
transform 1 0 39984 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_360
timestamp 1698431365
transform 1 0 41664 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_415
timestamp 1698431365
transform 1 0 47824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_419
timestamp 1698431365
transform 1 0 48272 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_18
timestamp 1698431365
transform 1 0 3360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_26
timestamp 1698431365
transform 1 0 4256 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_30
timestamp 1698431365
transform 1 0 4704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_57
timestamp 1698431365
transform 1 0 7728 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_88
timestamp 1698431365
transform 1 0 11200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_92
timestamp 1698431365
transform 1 0 11648 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_96
timestamp 1698431365
transform 1 0 12096 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_134
timestamp 1698431365
transform 1 0 16352 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_154
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_164
timestamp 1698431365
transform 1 0 19712 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_187
timestamp 1698431365
transform 1 0 22288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_226
timestamp 1698431365
transform 1 0 26656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_228
timestamp 1698431365
transform 1 0 26880 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_313
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_332
timestamp 1698431365
transform 1 0 38528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_334
timestamp 1698431365
transform 1 0 38752 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_364
timestamp 1698431365
transform 1 0 42112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_368
timestamp 1698431365
transform 1 0 42560 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_391
timestamp 1698431365
transform 1 0 45136 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_393
timestamp 1698431365
transform 1 0 45360 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_396
timestamp 1698431365
transform 1 0 45696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_400
timestamp 1698431365
transform 1 0 46144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_417
timestamp 1698431365
transform 1 0 48048 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_32
timestamp 1698431365
transform 1 0 4928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_34
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_37
timestamp 1698431365
transform 1 0 5488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_41
timestamp 1698431365
transform 1 0 5936 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_63
timestamp 1698431365
transform 1 0 8400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_67
timestamp 1698431365
transform 1 0 8848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_104
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_107
timestamp 1698431365
transform 1 0 13328 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_123
timestamp 1698431365
transform 1 0 15120 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_125
timestamp 1698431365
transform 1 0 15344 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_128
timestamp 1698431365
transform 1 0 15680 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_135
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1698431365
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_157
timestamp 1698431365
transform 1 0 18928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_165
timestamp 1698431365
transform 1 0 19824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_169
timestamp 1698431365
transform 1 0 20272 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_171
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_196
timestamp 1698431365
transform 1 0 23296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_200
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_216
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_237
timestamp 1698431365
transform 1 0 27888 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_290
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_292
timestamp 1698431365
transform 1 0 34048 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_315
timestamp 1698431365
transform 1 0 36624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_317
timestamp 1698431365
transform 1 0 36848 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_336
timestamp 1698431365
transform 1 0 38976 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_340
timestamp 1698431365
transform 1 0 39424 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_356
timestamp 1698431365
transform 1 0 41216 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_370
timestamp 1698431365
transform 1 0 42784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_387
timestamp 1698431365
transform 1 0 44688 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_395
timestamp 1698431365
transform 1 0 45584 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_399
timestamp 1698431365
transform 1 0 46032 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_406
timestamp 1698431365
transform 1 0 46816 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_414
timestamp 1698431365
transform 1 0 47712 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_418
timestamp 1698431365
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_420
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_6
timestamp 1698431365
transform 1 0 2016 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_13
timestamp 1698431365
transform 1 0 2800 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_17
timestamp 1698431365
transform 1 0 3248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_19
timestamp 1698431365
transform 1 0 3472 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_46
timestamp 1698431365
transform 1 0 6496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_50
timestamp 1698431365
transform 1 0 6944 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_85
timestamp 1698431365
transform 1 0 10864 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_93
timestamp 1698431365
transform 1 0 11760 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_141
timestamp 1698431365
transform 1 0 17136 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_150
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_166
timestamp 1698431365
transform 1 0 19936 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_183
timestamp 1698431365
transform 1 0 21840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_195
timestamp 1698431365
transform 1 0 23184 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_199
timestamp 1698431365
transform 1 0 23632 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_202
timestamp 1698431365
transform 1 0 23968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_255
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_282
timestamp 1698431365
transform 1 0 32928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_286
timestamp 1698431365
transform 1 0 33376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_297
timestamp 1698431365
transform 1 0 34608 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_310
timestamp 1698431365
transform 1 0 36064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_319
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_48
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_84
timestamp 1698431365
transform 1 0 10752 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_86
timestamp 1698431365
transform 1 0 10976 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_116
timestamp 1698431365
transform 1 0 14336 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_120
timestamp 1698431365
transform 1 0 14784 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_134
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_149
timestamp 1698431365
transform 1 0 18032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_153
timestamp 1698431365
transform 1 0 18480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_155
timestamp 1698431365
transform 1 0 18704 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_174
timestamp 1698431365
transform 1 0 20832 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_218
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_294
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_323
timestamp 1698431365
transform 1 0 37520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_327
timestamp 1698431365
transform 1 0 37968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_331
timestamp 1698431365
transform 1 0 38416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_335
timestamp 1698431365
transform 1 0 38864 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_343
timestamp 1698431365
transform 1 0 39760 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_354
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_357
timestamp 1698431365
transform 1 0 41328 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_389
timestamp 1698431365
transform 1 0 44912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_407
timestamp 1698431365
transform 1 0 46928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_415
timestamp 1698431365
transform 1 0 47824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_32
timestamp 1698431365
transform 1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_88
timestamp 1698431365
transform 1 0 11200 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_92
timestamp 1698431365
transform 1 0 11648 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_96
timestamp 1698431365
transform 1 0 12096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_98
timestamp 1698431365
transform 1 0 12320 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_118
timestamp 1698431365
transform 1 0 14560 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_134
timestamp 1698431365
transform 1 0 16352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_151
timestamp 1698431365
transform 1 0 18256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_153
timestamp 1698431365
transform 1 0 18480 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_196
timestamp 1698431365
transform 1 0 23296 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_207
timestamp 1698431365
transform 1 0 24528 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_209
timestamp 1698431365
transform 1 0 24752 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_228
timestamp 1698431365
transform 1 0 26880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_230
timestamp 1698431365
transform 1 0 27104 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_308
timestamp 1698431365
transform 1 0 35840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_324
timestamp 1698431365
transform 1 0 37632 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_328
timestamp 1698431365
transform 1 0 38080 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_358
timestamp 1698431365
transform 1 0 41440 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_362
timestamp 1698431365
transform 1 0 41888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_372
timestamp 1698431365
transform 1 0 43008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_380
timestamp 1698431365
transform 1 0 43904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_391
timestamp 1698431365
transform 1 0 45136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_395
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_403
timestamp 1698431365
transform 1 0 46480 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_419
timestamp 1698431365
transform 1 0 48272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_12
timestamp 1698431365
transform 1 0 2688 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_20
timestamp 1698431365
transform 1 0 3584 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_24
timestamp 1698431365
transform 1 0 4032 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_31
timestamp 1698431365
transform 1 0 4816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_35
timestamp 1698431365
transform 1 0 5264 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_67
timestamp 1698431365
transform 1 0 8848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_81
timestamp 1698431365
transform 1 0 10416 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_89
timestamp 1698431365
transform 1 0 11312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_119
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_158
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_175
timestamp 1698431365
transform 1 0 20944 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698431365
transform 1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_223
timestamp 1698431365
transform 1 0 26320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_225
timestamp 1698431365
transform 1 0 26544 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_339
timestamp 1698431365
transform 1 0 39312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_343
timestamp 1698431365
transform 1 0 39760 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_347
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_390
timestamp 1698431365
transform 1 0 45024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_392
timestamp 1698431365
transform 1 0 45248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_399
timestamp 1698431365
transform 1 0 46032 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_413
timestamp 1698431365
transform 1 0 47600 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_18
timestamp 1698431365
transform 1 0 3360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_53
timestamp 1698431365
transform 1 0 7280 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_89
timestamp 1698431365
transform 1 0 11312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_93
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_141
timestamp 1698431365
transform 1 0 17136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_143
timestamp 1698431365
transform 1 0 17360 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_150
timestamp 1698431365
transform 1 0 18144 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_164
timestamp 1698431365
transform 1 0 19712 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_168
timestamp 1698431365
transform 1 0 20160 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_179
timestamp 1698431365
transform 1 0 21392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_226
timestamp 1698431365
transform 1 0 26656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_233
timestamp 1698431365
transform 1 0 27440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_235
timestamp 1698431365
transform 1 0 27664 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_263
timestamp 1698431365
transform 1 0 30800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_265
timestamp 1698431365
transform 1 0 31024 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_268
timestamp 1698431365
transform 1 0 31360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_358
timestamp 1698431365
transform 1 0 41440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_362
timestamp 1698431365
transform 1 0 41888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_366
timestamp 1698431365
transform 1 0 42336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_368
timestamp 1698431365
transform 1 0 42560 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_32
timestamp 1698431365
transform 1 0 4928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_36
timestamp 1698431365
transform 1 0 5376 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_76
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_78
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_81
timestamp 1698431365
transform 1 0 10416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_83
timestamp 1698431365
transform 1 0 10640 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_86
timestamp 1698431365
transform 1 0 10976 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_90
timestamp 1698431365
transform 1 0 11424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_92
timestamp 1698431365
transform 1 0 11648 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_101
timestamp 1698431365
transform 1 0 12656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_105
timestamp 1698431365
transform 1 0 13104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_109
timestamp 1698431365
transform 1 0 13552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_111
timestamp 1698431365
transform 1 0 13776 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_120
timestamp 1698431365
transform 1 0 14784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_122
timestamp 1698431365
transform 1 0 15008 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_163
timestamp 1698431365
transform 1 0 19600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_186
timestamp 1698431365
transform 1 0 22176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_198
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698431365
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_218
timestamp 1698431365
transform 1 0 25760 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_226
timestamp 1698431365
transform 1 0 26656 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_245
timestamp 1698431365
transform 1 0 28784 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_360
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_364
timestamp 1698431365
transform 1 0 42112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_383
timestamp 1698431365
transform 1 0 44240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_412
timestamp 1698431365
transform 1 0 47488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_420
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_12
timestamp 1698431365
transform 1 0 2688 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_56
timestamp 1698431365
transform 1 0 7616 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_60
timestamp 1698431365
transform 1 0 8064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_62
timestamp 1698431365
transform 1 0 8288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_82
timestamp 1698431365
transform 1 0 10528 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_99
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_117
timestamp 1698431365
transform 1 0 14448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_121
timestamp 1698431365
transform 1 0 14896 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_125
timestamp 1698431365
transform 1 0 15344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_135
timestamp 1698431365
transform 1 0 16464 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_150
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_163
timestamp 1698431365
transform 1 0 19600 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_165
timestamp 1698431365
transform 1 0 19824 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_189
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_193
timestamp 1698431365
transform 1 0 22960 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_278
timestamp 1698431365
transform 1 0 32480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_308
timestamp 1698431365
transform 1 0 35840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698431365
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_391
timestamp 1698431365
transform 1 0 45136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_393
timestamp 1698431365
transform 1 0 45360 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_409
timestamp 1698431365
transform 1 0 47152 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_417
timestamp 1698431365
transform 1 0 48048 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_6
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_13
timestamp 1698431365
transform 1 0 2800 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_21
timestamp 1698431365
transform 1 0 3696 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_37
timestamp 1698431365
transform 1 0 5488 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_41
timestamp 1698431365
transform 1 0 5936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_43
timestamp 1698431365
transform 1 0 6160 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_50
timestamp 1698431365
transform 1 0 6944 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_87
timestamp 1698431365
transform 1 0 11088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_89
timestamp 1698431365
transform 1 0 11312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_101
timestamp 1698431365
transform 1 0 12656 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_107
timestamp 1698431365
transform 1 0 13328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_109
timestamp 1698431365
transform 1 0 13552 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_126
timestamp 1698431365
transform 1 0 15456 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_130
timestamp 1698431365
transform 1 0 15904 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_165
timestamp 1698431365
transform 1 0 19824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_169
timestamp 1698431365
transform 1 0 20272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_172
timestamp 1698431365
transform 1 0 20608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_176
timestamp 1698431365
transform 1 0 21056 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_184
timestamp 1698431365
transform 1 0 21952 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_187
timestamp 1698431365
transform 1 0 22288 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_195
timestamp 1698431365
transform 1 0 23184 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_236
timestamp 1698431365
transform 1 0 27776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_240
timestamp 1698431365
transform 1 0 28224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_254
timestamp 1698431365
transform 1 0 29792 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_258
timestamp 1698431365
transform 1 0 30240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_270
timestamp 1698431365
transform 1 0 31584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_299
timestamp 1698431365
transform 1 0 34832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_303
timestamp 1698431365
transform 1 0 35280 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_307
timestamp 1698431365
transform 1 0 35728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_343
timestamp 1698431365
transform 1 0 39760 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_347
timestamp 1698431365
transform 1 0 40208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_375
timestamp 1698431365
transform 1 0 43344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_379
timestamp 1698431365
transform 1 0 43792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_383
timestamp 1698431365
transform 1 0 44240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_41
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_51
timestamp 1698431365
transform 1 0 7056 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_55
timestamp 1698431365
transform 1 0 7504 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_65
timestamp 1698431365
transform 1 0 8624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_113
timestamp 1698431365
transform 1 0 14000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_170
timestamp 1698431365
transform 1 0 20384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_186
timestamp 1698431365
transform 1 0 22176 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_256
timestamp 1698431365
transform 1 0 30016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_260
timestamp 1698431365
transform 1 0 30464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_305
timestamp 1698431365
transform 1 0 35504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_420
timestamp 1698431365
transform 1 0 48384 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_74
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_109
timestamp 1698431365
transform 1 0 13552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_113
timestamp 1698431365
transform 1 0 14000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_117
timestamp 1698431365
transform 1 0 14448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_121
timestamp 1698431365
transform 1 0 14896 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_125
timestamp 1698431365
transform 1 0 15344 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_129
timestamp 1698431365
transform 1 0 15792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_131
timestamp 1698431365
transform 1 0 16016 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_234
timestamp 1698431365
transform 1 0 27552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_238
timestamp 1698431365
transform 1 0 28000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_242
timestamp 1698431365
transform 1 0 28448 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_261
timestamp 1698431365
transform 1 0 30576 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_269
timestamp 1698431365
transform 1 0 31472 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_273
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_296
timestamp 1698431365
transform 1 0 34496 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_330
timestamp 1698431365
transform 1 0 38304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_334
timestamp 1698431365
transform 1 0 38752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_378
timestamp 1698431365
transform 1 0 43680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_380
timestamp 1698431365
transform 1 0 43904 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_414
timestamp 1698431365
transform 1 0 47712 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_418
timestamp 1698431365
transform 1 0 48160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_420
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_16
timestamp 1698431365
transform 1 0 3136 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_39
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_55
timestamp 1698431365
transform 1 0 7504 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_61
timestamp 1698431365
transform 1 0 8176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_65
timestamp 1698431365
transform 1 0 8624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_69
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_102
timestamp 1698431365
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_118
timestamp 1698431365
transform 1 0 14560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_126
timestamp 1698431365
transform 1 0 15456 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_134
timestamp 1698431365
transform 1 0 16352 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_138
timestamp 1698431365
transform 1 0 16800 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_142
timestamp 1698431365
transform 1 0 17248 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_170
timestamp 1698431365
transform 1 0 20384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698431365
transform 1 0 21392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_182
timestamp 1698431365
transform 1 0 21728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_199
timestamp 1698431365
transform 1 0 23632 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_238
timestamp 1698431365
transform 1 0 28000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_251
timestamp 1698431365
transform 1 0 29456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_271
timestamp 1698431365
transform 1 0 31696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_290
timestamp 1698431365
transform 1 0 33824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_303
timestamp 1698431365
transform 1 0 35280 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_48
timestamp 1698431365
transform 1 0 6720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_52
timestamp 1698431365
transform 1 0 7168 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_133
timestamp 1698431365
transform 1 0 16240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_160
timestamp 1698431365
transform 1 0 19264 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_178
timestamp 1698431365
transform 1 0 21280 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_182
timestamp 1698431365
transform 1 0 21728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_184
timestamp 1698431365
transform 1 0 21952 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698431365
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698431365
transform 1 0 25312 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_242
timestamp 1698431365
transform 1 0 28448 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_256
timestamp 1698431365
transform 1 0 30016 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_264
timestamp 1698431365
transform 1 0 30912 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_268
timestamp 1698431365
transform 1 0 31360 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_299
timestamp 1698431365
transform 1 0 34832 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_303
timestamp 1698431365
transform 1 0 35280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_305
timestamp 1698431365
transform 1 0 35504 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_314
timestamp 1698431365
transform 1 0 36512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_6
timestamp 1698431365
transform 1 0 2016 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_13
timestamp 1698431365
transform 1 0 2800 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_29
timestamp 1698431365
transform 1 0 4592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_31
timestamp 1698431365
transform 1 0 4816 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_80
timestamp 1698431365
transform 1 0 10304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_84
timestamp 1698431365
transform 1 0 10752 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_131
timestamp 1698431365
transform 1 0 16016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_135
timestamp 1698431365
transform 1 0 16464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_181
timestamp 1698431365
transform 1 0 21616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_199
timestamp 1698431365
transform 1 0 23632 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_211
timestamp 1698431365
transform 1 0 24976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_215
timestamp 1698431365
transform 1 0 25424 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_219
timestamp 1698431365
transform 1 0 25872 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_227
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_255
timestamp 1698431365
transform 1 0 29904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_259
timestamp 1698431365
transform 1 0 30352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_276
timestamp 1698431365
transform 1 0 32256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_278
timestamp 1698431365
transform 1 0 32480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_285
timestamp 1698431365
transform 1 0 33264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_287
timestamp 1698431365
transform 1 0 33488 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_333
timestamp 1698431365
transform 1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_335
timestamp 1698431365
transform 1 0 38864 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_338
timestamp 1698431365
transform 1 0 39200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_372
timestamp 1698431365
transform 1 0 43008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_376
timestamp 1698431365
transform 1 0 43456 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_383
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_391
timestamp 1698431365
transform 1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_395
timestamp 1698431365
transform 1 0 45584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_403
timestamp 1698431365
transform 1 0 46480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_419
timestamp 1698431365
transform 1 0 48272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_32
timestamp 1698431365
transform 1 0 4928 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_48
timestamp 1698431365
transform 1 0 6720 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_56
timestamp 1698431365
transform 1 0 7616 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_74
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_90
timestamp 1698431365
transform 1 0 11424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_94
timestamp 1698431365
transform 1 0 11872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_98
timestamp 1698431365
transform 1 0 12320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_196
timestamp 1698431365
transform 1 0 23296 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_204
timestamp 1698431365
transform 1 0 24192 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698431365
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_234
timestamp 1698431365
transform 1 0 27552 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_250
timestamp 1698431365
transform 1 0 29344 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_254
timestamp 1698431365
transform 1 0 29792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_319
timestamp 1698431365
transform 1 0 37072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_323
timestamp 1698431365
transform 1 0 37520 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_329
timestamp 1698431365
transform 1 0 38192 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_333
timestamp 1698431365
transform 1 0 38640 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_336
timestamp 1698431365
transform 1 0 38976 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_340
timestamp 1698431365
transform 1 0 39424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_367
timestamp 1698431365
transform 1 0 42448 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_390
timestamp 1698431365
transform 1 0 45024 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_16
timestamp 1698431365
transform 1 0 3136 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_49
timestamp 1698431365
transform 1 0 6832 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_53
timestamp 1698431365
transform 1 0 7280 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_55
timestamp 1698431365
transform 1 0 7504 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_129
timestamp 1698431365
transform 1 0 15792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_143
timestamp 1698431365
transform 1 0 17360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_147
timestamp 1698431365
transform 1 0 17808 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_163
timestamp 1698431365
transform 1 0 19600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_183
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_188
timestamp 1698431365
transform 1 0 22400 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_234
timestamp 1698431365
transform 1 0 27552 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_238
timestamp 1698431365
transform 1 0 28000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_261
timestamp 1698431365
transform 1 0 30576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_265
timestamp 1698431365
transform 1 0 31024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_269
timestamp 1698431365
transform 1 0 31472 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_273
timestamp 1698431365
transform 1 0 31920 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_335
timestamp 1698431365
transform 1 0 38864 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_362
timestamp 1698431365
transform 1 0 41888 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_378
timestamp 1698431365
transform 1 0 43680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_382
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_395
timestamp 1698431365
transform 1 0 45584 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_399
timestamp 1698431365
transform 1 0 46032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_407
timestamp 1698431365
transform 1 0 46928 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_415
timestamp 1698431365
transform 1 0 47824 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_419
timestamp 1698431365
transform 1 0 48272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_34
timestamp 1698431365
transform 1 0 5152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_79
timestamp 1698431365
transform 1 0 10192 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_83
timestamp 1698431365
transform 1 0 10640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_117
timestamp 1698431365
transform 1 0 14448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_121
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_125
timestamp 1698431365
transform 1 0 15344 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_133
timestamp 1698431365
transform 1 0 16240 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698431365
transform 1 0 16688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_176
timestamp 1698431365
transform 1 0 21056 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_192
timestamp 1698431365
transform 1 0 22848 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_200
timestamp 1698431365
transform 1 0 23744 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_234
timestamp 1698431365
transform 1 0 27552 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_238
timestamp 1698431365
transform 1 0 28000 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_242
timestamp 1698431365
transform 1 0 28448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_246
timestamp 1698431365
transform 1 0 28896 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_263
timestamp 1698431365
transform 1 0 30800 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_298
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_337
timestamp 1698431365
transform 1 0 39088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_345
timestamp 1698431365
transform 1 0 39984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_362
timestamp 1698431365
transform 1 0 41888 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_393
timestamp 1698431365
transform 1 0 45360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_397
timestamp 1698431365
transform 1 0 45808 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_413
timestamp 1698431365
transform 1 0 47600 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_53
timestamp 1698431365
transform 1 0 7280 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_93
timestamp 1698431365
transform 1 0 11760 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_113
timestamp 1698431365
transform 1 0 14000 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_145
timestamp 1698431365
transform 1 0 17584 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_168
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_190
timestamp 1698431365
transform 1 0 22624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_200
timestamp 1698431365
transform 1 0 23744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_202
timestamp 1698431365
transform 1 0 23968 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_210
timestamp 1698431365
transform 1 0 24864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_212
timestamp 1698431365
transform 1 0 25088 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_223
timestamp 1698431365
transform 1 0 26320 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_282
timestamp 1698431365
transform 1 0 32928 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_346
timestamp 1698431365
transform 1 0 40096 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_350
timestamp 1698431365
transform 1 0 40544 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_358
timestamp 1698431365
transform 1 0 41440 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_360
timestamp 1698431365
transform 1 0 41664 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_382
timestamp 1698431365
transform 1 0 44128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_391
timestamp 1698431365
transform 1 0 45136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_410
timestamp 1698431365
transform 1 0 47264 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_418
timestamp 1698431365
transform 1 0 48160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_420
timestamp 1698431365
transform 1 0 48384 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_32
timestamp 1698431365
transform 1 0 4928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_36
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_52
timestamp 1698431365
transform 1 0 7168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_60
timestamp 1698431365
transform 1 0 8064 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_81
timestamp 1698431365
transform 1 0 10416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_85
timestamp 1698431365
transform 1 0 10864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_89
timestamp 1698431365
transform 1 0 11312 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_97
timestamp 1698431365
transform 1 0 12208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_101
timestamp 1698431365
transform 1 0 12656 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_109
timestamp 1698431365
transform 1 0 13552 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_125
timestamp 1698431365
transform 1 0 15344 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_133
timestamp 1698431365
transform 1 0 16240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_135
timestamp 1698431365
transform 1 0 16464 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_158
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_170
timestamp 1698431365
transform 1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_174
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_178
timestamp 1698431365
transform 1 0 21280 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_274
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_310
timestamp 1698431365
transform 1 0 36064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_318
timestamp 1698431365
transform 1 0 36960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_324
timestamp 1698431365
transform 1 0 37632 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_340
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_342
timestamp 1698431365
transform 1 0 39648 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_345
timestamp 1698431365
transform 1 0 39984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_347
timestamp 1698431365
transform 1 0 40208 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_375
timestamp 1698431365
transform 1 0 43344 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_383
timestamp 1698431365
transform 1 0 44240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_387
timestamp 1698431365
transform 1 0 44688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_6
timestamp 1698431365
transform 1 0 2016 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_13
timestamp 1698431365
transform 1 0 2800 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_17
timestamp 1698431365
transform 1 0 3248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_19
timestamp 1698431365
transform 1 0 3472 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_75
timestamp 1698431365
transform 1 0 9744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_79
timestamp 1698431365
transform 1 0 10192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_99
timestamp 1698431365
transform 1 0 12432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_148
timestamp 1698431365
transform 1 0 17920 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_156
timestamp 1698431365
transform 1 0 18816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_160
timestamp 1698431365
transform 1 0 19264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_170
timestamp 1698431365
transform 1 0 20384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_183
timestamp 1698431365
transform 1 0 21840 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_191
timestamp 1698431365
transform 1 0 22736 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_195
timestamp 1698431365
transform 1 0 23184 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_202
timestamp 1698431365
transform 1 0 23968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_204
timestamp 1698431365
transform 1 0 24192 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_209
timestamp 1698431365
transform 1 0 24752 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_213
timestamp 1698431365
transform 1 0 25200 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_221
timestamp 1698431365
transform 1 0 26096 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_223
timestamp 1698431365
transform 1 0 26320 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_230
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_234
timestamp 1698431365
transform 1 0 27552 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_253
timestamp 1698431365
transform 1 0 29680 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_257
timestamp 1698431365
transform 1 0 30128 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_293
timestamp 1698431365
transform 1 0 34160 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_297
timestamp 1698431365
transform 1 0 34608 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_308
timestamp 1698431365
transform 1 0 35840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_329
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_333
timestamp 1698431365
transform 1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_366
timestamp 1698431365
transform 1 0 42336 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_395
timestamp 1698431365
transform 1 0 45584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_397
timestamp 1698431365
transform 1 0 45808 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_419
timestamp 1698431365
transform 1 0 48272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_6
timestamp 1698431365
transform 1 0 2016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_8
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_15
timestamp 1698431365
transform 1 0 3024 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_19
timestamp 1698431365
transform 1 0 3472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_21
timestamp 1698431365
transform 1 0 3696 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_37
timestamp 1698431365
transform 1 0 5488 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_39
timestamp 1698431365
transform 1 0 5712 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_125
timestamp 1698431365
transform 1 0 15344 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_133
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_152
timestamp 1698431365
transform 1 0 18368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_186
timestamp 1698431365
transform 1 0 22176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_190
timestamp 1698431365
transform 1 0 22624 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_198
timestamp 1698431365
transform 1 0 23520 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_202
timestamp 1698431365
transform 1 0 23968 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_205
timestamp 1698431365
transform 1 0 24304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_218
timestamp 1698431365
transform 1 0 25760 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_271
timestamp 1698431365
transform 1 0 31696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_275
timestamp 1698431365
transform 1 0 32144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_299
timestamp 1698431365
transform 1 0 34832 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_338
timestamp 1698431365
transform 1 0 39200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_342
timestamp 1698431365
transform 1 0 39648 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_407
timestamp 1698431365
transform 1 0 46928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_411
timestamp 1698431365
transform 1 0 47376 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_33
timestamp 1698431365
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_53
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_57
timestamp 1698431365
transform 1 0 7728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_67
timestamp 1698431365
transform 1 0 8848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_71
timestamp 1698431365
transform 1 0 9296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_73
timestamp 1698431365
transform 1 0 9520 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_78
timestamp 1698431365
transform 1 0 10080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_87
timestamp 1698431365
transform 1 0 11088 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_89
timestamp 1698431365
transform 1 0 11312 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_96
timestamp 1698431365
transform 1 0 12096 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_119
timestamp 1698431365
transform 1 0 14672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_123
timestamp 1698431365
transform 1 0 15120 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_131
timestamp 1698431365
transform 1 0 16016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_141
timestamp 1698431365
transform 1 0 17136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_145
timestamp 1698431365
transform 1 0 17584 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_155
timestamp 1698431365
transform 1 0 18704 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_159
timestamp 1698431365
transform 1 0 19152 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_192
timestamp 1698431365
transform 1 0 22848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_196
timestamp 1698431365
transform 1 0 23296 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_235
timestamp 1698431365
transform 1 0 27664 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698431365
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_249
timestamp 1698431365
transform 1 0 29232 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_264
timestamp 1698431365
transform 1 0 30912 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_281
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_289
timestamp 1698431365
transform 1 0 33712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_291
timestamp 1698431365
transform 1 0 33936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_331
timestamp 1698431365
transform 1 0 38416 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_365
timestamp 1698431365
transform 1 0 42224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_367
timestamp 1698431365
transform 1 0 42448 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_374
timestamp 1698431365
transform 1 0 43232 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_382
timestamp 1698431365
transform 1 0 44128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_391
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_393
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_419
timestamp 1698431365
transform 1 0 48272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_104
timestamp 1698431365
transform 1 0 12992 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_120
timestamp 1698431365
transform 1 0 14784 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_124
timestamp 1698431365
transform 1 0 15232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_134
timestamp 1698431365
transform 1 0 16352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_138
timestamp 1698431365
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_144
timestamp 1698431365
transform 1 0 17472 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_161
timestamp 1698431365
transform 1 0 19376 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_177
timestamp 1698431365
transform 1 0 21168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_179
timestamp 1698431365
transform 1 0 21392 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_218
timestamp 1698431365
transform 1 0 25760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_222
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_252
timestamp 1698431365
transform 1 0 29568 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_256
timestamp 1698431365
transform 1 0 30016 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_263
timestamp 1698431365
transform 1 0 30800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_265
timestamp 1698431365
transform 1 0 31024 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_274
timestamp 1698431365
transform 1 0 32032 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_288
timestamp 1698431365
transform 1 0 33600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_298
timestamp 1698431365
transform 1 0 34720 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_321
timestamp 1698431365
transform 1 0 37296 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_329
timestamp 1698431365
transform 1 0 38192 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_348
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_358
timestamp 1698431365
transform 1 0 41440 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_360
timestamp 1698431365
transform 1 0 41664 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_41
timestamp 1698431365
transform 1 0 5936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_45
timestamp 1698431365
transform 1 0 6384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_47
timestamp 1698431365
transform 1 0 6608 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_54
timestamp 1698431365
transform 1 0 7392 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_73
timestamp 1698431365
transform 1 0 9520 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_77
timestamp 1698431365
transform 1 0 9968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_85
timestamp 1698431365
transform 1 0 10864 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_89
timestamp 1698431365
transform 1 0 11312 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_123
timestamp 1698431365
transform 1 0 15120 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_127
timestamp 1698431365
transform 1 0 15568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_129
timestamp 1698431365
transform 1 0 15792 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_136
timestamp 1698431365
transform 1 0 16576 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_144
timestamp 1698431365
transform 1 0 17472 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_151
timestamp 1698431365
transform 1 0 18256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_155
timestamp 1698431365
transform 1 0 18704 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_159
timestamp 1698431365
transform 1 0 19152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_187
timestamp 1698431365
transform 1 0 22288 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_190
timestamp 1698431365
transform 1 0 22624 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_197
timestamp 1698431365
transform 1 0 23408 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_201
timestamp 1698431365
transform 1 0 23856 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_209
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_212
timestamp 1698431365
transform 1 0 25088 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_220
timestamp 1698431365
transform 1 0 25984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_236
timestamp 1698431365
transform 1 0 27776 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_251
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_261
timestamp 1698431365
transform 1 0 30576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_265
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_273
timestamp 1698431365
transform 1 0 31920 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_303
timestamp 1698431365
transform 1 0 35280 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_307
timestamp 1698431365
transform 1 0 35728 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_321
timestamp 1698431365
transform 1 0 37296 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_338
timestamp 1698431365
transform 1 0 39200 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_342
timestamp 1698431365
transform 1 0 39648 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_364
timestamp 1698431365
transform 1 0 42112 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_368
timestamp 1698431365
transform 1 0 42560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_391
timestamp 1698431365
transform 1 0 45136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_393
timestamp 1698431365
transform 1 0 45360 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_402
timestamp 1698431365
transform 1 0 46368 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_412
timestamp 1698431365
transform 1 0 47488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_420
timestamp 1698431365
transform 1 0 48384 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_12
timestamp 1698431365
transform 1 0 2688 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_20
timestamp 1698431365
transform 1 0 3584 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_102
timestamp 1698431365
transform 1 0 12768 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_106
timestamp 1698431365
transform 1 0 13216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_123
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_127
timestamp 1698431365
transform 1 0 15568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_135
timestamp 1698431365
transform 1 0 16464 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_152
timestamp 1698431365
transform 1 0 18368 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_193
timestamp 1698431365
transform 1 0 22960 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_197
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_222
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_226
timestamp 1698431365
transform 1 0 26656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_243
timestamp 1698431365
transform 1 0 28560 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_251
timestamp 1698431365
transform 1 0 29456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_261
timestamp 1698431365
transform 1 0 30576 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_286
timestamp 1698431365
transform 1 0 33376 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_294
timestamp 1698431365
transform 1 0 34272 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_298
timestamp 1698431365
transform 1 0 34720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_308
timestamp 1698431365
transform 1 0 35840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_310
timestamp 1698431365
transform 1 0 36064 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_341
timestamp 1698431365
transform 1 0 39536 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_345
timestamp 1698431365
transform 1 0 39984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_347
timestamp 1698431365
transform 1 0 40208 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_362
timestamp 1698431365
transform 1 0 41888 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_364
timestamp 1698431365
transform 1 0 42112 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_395
timestamp 1698431365
transform 1 0 45584 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_399
timestamp 1698431365
transform 1 0 46032 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_401
timestamp 1698431365
transform 1 0 46256 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_417
timestamp 1698431365
transform 1 0 48048 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_12
timestamp 1698431365
transform 1 0 2688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_16
timestamp 1698431365
transform 1 0 3136 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_33
timestamp 1698431365
transform 1 0 5040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_69
timestamp 1698431365
transform 1 0 9072 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_85
timestamp 1698431365
transform 1 0 10864 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_89
timestamp 1698431365
transform 1 0 11312 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_98
timestamp 1698431365
transform 1 0 12320 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_115
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_119
timestamp 1698431365
transform 1 0 14672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_121
timestamp 1698431365
transform 1 0 14896 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_158
timestamp 1698431365
transform 1 0 19040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_209
timestamp 1698431365
transform 1 0 24752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_213
timestamp 1698431365
transform 1 0 25200 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_217
timestamp 1698431365
transform 1 0 25648 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_235
timestamp 1698431365
transform 1 0 27664 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_239
timestamp 1698431365
transform 1 0 28112 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_253
timestamp 1698431365
transform 1 0 29680 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_276
timestamp 1698431365
transform 1 0 32256 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_294
timestamp 1698431365
transform 1 0 34272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_298
timestamp 1698431365
transform 1 0 34720 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_306
timestamp 1698431365
transform 1 0 35616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_310
timestamp 1698431365
transform 1 0 36064 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_324
timestamp 1698431365
transform 1 0 37632 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_340
timestamp 1698431365
transform 1 0 39424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_342
timestamp 1698431365
transform 1 0 39648 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_382
timestamp 1698431365
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_32
timestamp 1698431365
transform 1 0 4928 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_41
timestamp 1698431365
transform 1 0 5936 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_45
timestamp 1698431365
transform 1 0 6384 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_81
timestamp 1698431365
transform 1 0 10416 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_92
timestamp 1698431365
transform 1 0 11648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_94
timestamp 1698431365
transform 1 0 11872 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_113
timestamp 1698431365
transform 1 0 14000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_117
timestamp 1698431365
transform 1 0 14448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_121
timestamp 1698431365
transform 1 0 14896 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_128
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_150
timestamp 1698431365
transform 1 0 18144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_154
timestamp 1698431365
transform 1 0 18592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_158
timestamp 1698431365
transform 1 0 19040 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_162
timestamp 1698431365
transform 1 0 19488 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_166
timestamp 1698431365
transform 1 0 19936 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_176
timestamp 1698431365
transform 1 0 21056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_180
timestamp 1698431365
transform 1 0 21504 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_196
timestamp 1698431365
transform 1 0 23296 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_204
timestamp 1698431365
transform 1 0 24192 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_208
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_250
timestamp 1698431365
transform 1 0 29344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_266
timestamp 1698431365
transform 1 0 31136 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_293
timestamp 1698431365
transform 1 0 34160 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_301
timestamp 1698431365
transform 1 0 35056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_333
timestamp 1698431365
transform 1 0 38640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_337
timestamp 1698431365
transform 1 0 39088 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_348
timestamp 1698431365
transform 1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_370
timestamp 1698431365
transform 1 0 42784 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_374
timestamp 1698431365
transform 1 0 43232 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_390
timestamp 1698431365
transform 1 0 45024 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_398
timestamp 1698431365
transform 1 0 45920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_406
timestamp 1698431365
transform 1 0 46816 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_414
timestamp 1698431365
transform 1 0 47712 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_418
timestamp 1698431365
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_420
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_10
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_14
timestamp 1698431365
transform 1 0 2912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_16
timestamp 1698431365
transform 1 0 3136 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_39
timestamp 1698431365
transform 1 0 5712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_70
timestamp 1698431365
transform 1 0 9184 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_87
timestamp 1698431365
transform 1 0 11088 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_91
timestamp 1698431365
transform 1 0 11536 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_94
timestamp 1698431365
transform 1 0 11872 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_113
timestamp 1698431365
transform 1 0 14000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_117
timestamp 1698431365
transform 1 0 14448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_139
timestamp 1698431365
transform 1 0 16912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_143
timestamp 1698431365
transform 1 0 17360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_145
timestamp 1698431365
transform 1 0 17584 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_148
timestamp 1698431365
transform 1 0 17920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_152
timestamp 1698431365
transform 1 0 18368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_156
timestamp 1698431365
transform 1 0 18816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_158
timestamp 1698431365
transform 1 0 19040 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_167
timestamp 1698431365
transform 1 0 20048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_212
timestamp 1698431365
transform 1 0 25088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_216
timestamp 1698431365
transform 1 0 25536 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_224
timestamp 1698431365
transform 1 0 26432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_232
timestamp 1698431365
transform 1 0 27328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_236
timestamp 1698431365
transform 1 0 27776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_249
timestamp 1698431365
transform 1 0 29232 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_258
timestamp 1698431365
transform 1 0 30240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_260
timestamp 1698431365
transform 1 0 30464 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_267
timestamp 1698431365
transform 1 0 31248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_271
timestamp 1698431365
transform 1 0 31696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_275
timestamp 1698431365
transform 1 0 32144 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_286
timestamp 1698431365
transform 1 0 33376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_292
timestamp 1698431365
transform 1 0 34048 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_323
timestamp 1698431365
transform 1 0 37520 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_369
timestamp 1698431365
transform 1 0 42672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_6
timestamp 1698431365
transform 1 0 2016 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_14
timestamp 1698431365
transform 1 0 2912 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_22
timestamp 1698431365
transform 1 0 3808 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_46
timestamp 1698431365
transform 1 0 6496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_50
timestamp 1698431365
transform 1 0 6944 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_74
timestamp 1698431365
transform 1 0 9632 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_109
timestamp 1698431365
transform 1 0 13552 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_164
timestamp 1698431365
transform 1 0 19712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_168
timestamp 1698431365
transform 1 0 20160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_174
timestamp 1698431365
transform 1 0 20832 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_239
timestamp 1698431365
transform 1 0 28112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_241
timestamp 1698431365
transform 1 0 28336 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_267
timestamp 1698431365
transform 1 0 31248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_271
timestamp 1698431365
transform 1 0 31696 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_298
timestamp 1698431365
transform 1 0 34720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_302
timestamp 1698431365
transform 1 0 35168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_319
timestamp 1698431365
transform 1 0 37072 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_323
timestamp 1698431365
transform 1 0 37520 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_340
timestamp 1698431365
transform 1 0 39424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_344
timestamp 1698431365
transform 1 0 39872 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_348
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_356
timestamp 1698431365
transform 1 0 41216 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_417
timestamp 1698431365
transform 1 0 48048 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_41
timestamp 1698431365
transform 1 0 5936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_43
timestamp 1698431365
transform 1 0 6160 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_50
timestamp 1698431365
transform 1 0 6944 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_54
timestamp 1698431365
transform 1 0 7392 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_56
timestamp 1698431365
transform 1 0 7616 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_72
timestamp 1698431365
transform 1 0 9408 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_76
timestamp 1698431365
transform 1 0 9856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_78
timestamp 1698431365
transform 1 0 10080 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_113
timestamp 1698431365
transform 1 0 14000 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_123
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_127
timestamp 1698431365
transform 1 0 15568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_135
timestamp 1698431365
transform 1 0 16464 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_141
timestamp 1698431365
transform 1 0 17136 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_145
timestamp 1698431365
transform 1 0 17584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_147
timestamp 1698431365
transform 1 0 17808 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_160
timestamp 1698431365
transform 1 0 19264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_162
timestamp 1698431365
transform 1 0 19488 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_189
timestamp 1698431365
transform 1 0 22512 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_193
timestamp 1698431365
transform 1 0 22960 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_197
timestamp 1698431365
transform 1 0 23408 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_205
timestamp 1698431365
transform 1 0 24304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_294
timestamp 1698431365
transform 1 0 34272 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_298
timestamp 1698431365
transform 1 0 34720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_321
timestamp 1698431365
transform 1 0 37296 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_380
timestamp 1698431365
transform 1 0 43904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_395
timestamp 1698431365
transform 1 0 45584 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_405
timestamp 1698431365
transform 1 0 46704 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_34
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_87
timestamp 1698431365
transform 1 0 11088 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_120
timestamp 1698431365
transform 1 0 14784 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_124
timestamp 1698431365
transform 1 0 15232 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_127
timestamp 1698431365
transform 1 0 15568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_178
timestamp 1698431365
transform 1 0 21280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_201
timestamp 1698431365
transform 1 0 23856 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_205
timestamp 1698431365
transform 1 0 24304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_219
timestamp 1698431365
transform 1 0 25872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_231
timestamp 1698431365
transform 1 0 27216 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_243
timestamp 1698431365
transform 1 0 28560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_245
timestamp 1698431365
transform 1 0 28784 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_262
timestamp 1698431365
transform 1 0 30688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_266
timestamp 1698431365
transform 1 0 31136 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_270
timestamp 1698431365
transform 1 0 31584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_292
timestamp 1698431365
transform 1 0 34048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_354
timestamp 1698431365
transform 1 0 40992 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_372
timestamp 1698431365
transform 1 0 43008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_376
timestamp 1698431365
transform 1 0 43456 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_408
timestamp 1698431365
transform 1 0 47040 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698431365
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_420
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_6
timestamp 1698431365
transform 1 0 2016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_8
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_15
timestamp 1698431365
transform 1 0 3024 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_31
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_52
timestamp 1698431365
transform 1 0 7168 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_56
timestamp 1698431365
transform 1 0 7616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_58
timestamp 1698431365
transform 1 0 7840 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_74
timestamp 1698431365
transform 1 0 9632 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_76
timestamp 1698431365
transform 1 0 9856 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_79
timestamp 1698431365
transform 1 0 10192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_96
timestamp 1698431365
transform 1 0 12096 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_111
timestamp 1698431365
transform 1 0 13776 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_159
timestamp 1698431365
transform 1 0 19152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_170
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_202
timestamp 1698431365
transform 1 0 23968 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_213
timestamp 1698431365
transform 1 0 25200 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_217
timestamp 1698431365
transform 1 0 25648 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_227
timestamp 1698431365
transform 1 0 26768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_231
timestamp 1698431365
transform 1 0 27216 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_242
timestamp 1698431365
transform 1 0 28448 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_251
timestamp 1698431365
transform 1 0 29456 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_262
timestamp 1698431365
transform 1 0 30688 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_268
timestamp 1698431365
transform 1 0 31360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_272
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_306
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_321
timestamp 1698431365
transform 1 0 37296 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_324
timestamp 1698431365
transform 1 0 37632 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_340
timestamp 1698431365
transform 1 0 39424 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_348
timestamp 1698431365
transform 1 0 40320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_352
timestamp 1698431365
transform 1 0 40768 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_368
timestamp 1698431365
transform 1 0 42560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_391
timestamp 1698431365
transform 1 0 45136 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_407
timestamp 1698431365
transform 1 0 46928 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_415
timestamp 1698431365
transform 1 0 47824 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_419
timestamp 1698431365
transform 1 0 48272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_32
timestamp 1698431365
transform 1 0 4928 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_36
timestamp 1698431365
transform 1 0 5376 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_74
timestamp 1698431365
transform 1 0 9632 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_116
timestamp 1698431365
transform 1 0 14336 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_120
timestamp 1698431365
transform 1 0 14784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_138
timestamp 1698431365
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_169
timestamp 1698431365
transform 1 0 20272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_173
timestamp 1698431365
transform 1 0 20720 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_177
timestamp 1698431365
transform 1 0 21168 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_180
timestamp 1698431365
transform 1 0 21504 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_222
timestamp 1698431365
transform 1 0 26208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_226
timestamp 1698431365
transform 1 0 26656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_228
timestamp 1698431365
transform 1 0 26880 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_231
timestamp 1698431365
transform 1 0 27216 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_239
timestamp 1698431365
transform 1 0 28112 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_242
timestamp 1698431365
transform 1 0 28448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_261
timestamp 1698431365
transform 1 0 30576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_265
timestamp 1698431365
transform 1 0 31024 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_269
timestamp 1698431365
transform 1 0 31472 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_272
timestamp 1698431365
transform 1 0 31808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_308
timestamp 1698431365
transform 1 0 35840 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_316
timestamp 1698431365
transform 1 0 36736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_368
timestamp 1698431365
transform 1 0 42560 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_405
timestamp 1698431365
transform 1 0 46704 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_6
timestamp 1698431365
transform 1 0 2016 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_13
timestamp 1698431365
transform 1 0 2800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_17
timestamp 1698431365
transform 1 0 3248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_19
timestamp 1698431365
transform 1 0 3472 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_52
timestamp 1698431365
transform 1 0 7168 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_59
timestamp 1698431365
transform 1 0 7952 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_67
timestamp 1698431365
transform 1 0 8848 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_111
timestamp 1698431365
transform 1 0 13776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_123
timestamp 1698431365
transform 1 0 15120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_127
timestamp 1698431365
transform 1 0 15568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_131
timestamp 1698431365
transform 1 0 16016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_149
timestamp 1698431365
transform 1 0 18032 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_153
timestamp 1698431365
transform 1 0 18480 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698431365
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_191
timestamp 1698431365
transform 1 0 22736 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_200
timestamp 1698431365
transform 1 0 23744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_202
timestamp 1698431365
transform 1 0 23968 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_210
timestamp 1698431365
transform 1 0 24864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_212
timestamp 1698431365
transform 1 0 25088 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_228
timestamp 1698431365
transform 1 0 26880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_230
timestamp 1698431365
transform 1 0 27104 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_251
timestamp 1698431365
transform 1 0 29456 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_255
timestamp 1698431365
transform 1 0 29904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_259
timestamp 1698431365
transform 1 0 30352 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_261
timestamp 1698431365
transform 1 0 30576 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_292
timestamp 1698431365
transform 1 0 34048 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_296
timestamp 1698431365
transform 1 0 34496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_300
timestamp 1698431365
transform 1 0 34944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_310
timestamp 1698431365
transform 1 0 36064 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698431365
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_347
timestamp 1698431365
transform 1 0 40208 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_349
timestamp 1698431365
transform 1 0 40432 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_380
timestamp 1698431365
transform 1 0 43904 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_419
timestamp 1698431365
transform 1 0 48272 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_32
timestamp 1698431365
transform 1 0 4928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_36
timestamp 1698431365
transform 1 0 5376 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_76
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_86
timestamp 1698431365
transform 1 0 10976 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_134
timestamp 1698431365
transform 1 0 16352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_138
timestamp 1698431365
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_150
timestamp 1698431365
transform 1 0 18144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_157
timestamp 1698431365
transform 1 0 18928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_165
timestamp 1698431365
transform 1 0 19824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_197
timestamp 1698431365
transform 1 0 23408 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_201
timestamp 1698431365
transform 1 0 23856 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_214
timestamp 1698431365
transform 1 0 25312 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_225
timestamp 1698431365
transform 1 0 26544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_252
timestamp 1698431365
transform 1 0 29568 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_256
timestamp 1698431365
transform 1 0 30016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_258
timestamp 1698431365
transform 1 0 30240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_290
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_306
timestamp 1698431365
transform 1 0 35616 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_343
timestamp 1698431365
transform 1 0 39760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_347
timestamp 1698431365
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_349
timestamp 1698431365
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_358
timestamp 1698431365
transform 1 0 41440 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_390
timestamp 1698431365
transform 1 0 45024 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_406
timestamp 1698431365
transform 1 0 46816 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_414
timestamp 1698431365
transform 1 0 47712 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_420
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_10
timestamp 1698431365
transform 1 0 2464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_14
timestamp 1698431365
transform 1 0 2912 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_22
timestamp 1698431365
transform 1 0 3808 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_30
timestamp 1698431365
transform 1 0 4704 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_41
timestamp 1698431365
transform 1 0 5936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_45
timestamp 1698431365
transform 1 0 6384 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_61
timestamp 1698431365
transform 1 0 8176 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_69
timestamp 1698431365
transform 1 0 9072 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_72
timestamp 1698431365
transform 1 0 9408 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_88
timestamp 1698431365
transform 1 0 11200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_90
timestamp 1698431365
transform 1 0 11424 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_121
timestamp 1698431365
transform 1 0 14896 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_167
timestamp 1698431365
transform 1 0 20048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_179
timestamp 1698431365
transform 1 0 21392 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_195
timestamp 1698431365
transform 1 0 23184 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_226
timestamp 1698431365
transform 1 0 26656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_228
timestamp 1698431365
transform 1 0 26880 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_235
timestamp 1698431365
transform 1 0 27664 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_255
timestamp 1698431365
transform 1 0 29904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_259
timestamp 1698431365
transform 1 0 30352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_262
timestamp 1698431365
transform 1 0 30688 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_294
timestamp 1698431365
transform 1 0 34272 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_303
timestamp 1698431365
transform 1 0 35280 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_323
timestamp 1698431365
transform 1 0 37520 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_339
timestamp 1698431365
transform 1 0 39312 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_347
timestamp 1698431365
transform 1 0 40208 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_350
timestamp 1698431365
transform 1 0 40544 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_358
timestamp 1698431365
transform 1 0 41440 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_362
timestamp 1698431365
transform 1 0 41888 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_370
timestamp 1698431365
transform 1 0 42784 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_378
timestamp 1698431365
transform 1 0 43680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_419
timestamp 1698431365
transform 1 0 48272 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_6
timestamp 1698431365
transform 1 0 2016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_8
timestamp 1698431365
transform 1 0 2240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_39
timestamp 1698431365
transform 1 0 5712 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_87
timestamp 1698431365
transform 1 0 11088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_95
timestamp 1698431365
transform 1 0 11984 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_131
timestamp 1698431365
transform 1 0 16016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_135
timestamp 1698431365
transform 1 0 16464 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698431365
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_157
timestamp 1698431365
transform 1 0 18928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_161
timestamp 1698431365
transform 1 0 19376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_165
timestamp 1698431365
transform 1 0 19824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_169
timestamp 1698431365
transform 1 0 20272 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_173
timestamp 1698431365
transform 1 0 20720 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_176
timestamp 1698431365
transform 1 0 21056 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_180
timestamp 1698431365
transform 1 0 21504 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_183
timestamp 1698431365
transform 1 0 21840 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_191
timestamp 1698431365
transform 1 0 22736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_195
timestamp 1698431365
transform 1 0 23184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_199
timestamp 1698431365
transform 1 0 23632 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_205
timestamp 1698431365
transform 1 0 24304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_227
timestamp 1698431365
transform 1 0 26768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_229
timestamp 1698431365
transform 1 0 26992 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_275
timestamp 1698431365
transform 1 0 32144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_277
timestamp 1698431365
transform 1 0 32368 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_288
timestamp 1698431365
transform 1 0 33600 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_320
timestamp 1698431365
transform 1 0 37184 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_328
timestamp 1698431365
transform 1 0 38080 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_332
timestamp 1698431365
transform 1 0 38528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_334
timestamp 1698431365
transform 1 0 38752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_392
timestamp 1698431365
transform 1 0 45248 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_408
timestamp 1698431365
transform 1 0 47040 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_420
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_41
timestamp 1698431365
transform 1 0 5936 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_43
timestamp 1698431365
transform 1 0 6160 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_50
timestamp 1698431365
transform 1 0 6944 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_66
timestamp 1698431365
transform 1 0 8736 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_70
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_127
timestamp 1698431365
transform 1 0 15568 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_161
timestamp 1698431365
transform 1 0 19376 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_165
timestamp 1698431365
transform 1 0 19824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_173
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_192
timestamp 1698431365
transform 1 0 22848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_196
timestamp 1698431365
transform 1 0 23296 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_200
timestamp 1698431365
transform 1 0 23744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_208
timestamp 1698431365
transform 1 0 24640 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_224
timestamp 1698431365
transform 1 0 26432 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_233
timestamp 1698431365
transform 1 0 27440 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_237
timestamp 1698431365
transform 1 0 27888 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_249
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_280
timestamp 1698431365
transform 1 0 32704 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_296
timestamp 1698431365
transform 1 0 34496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_313
timestamp 1698431365
transform 1 0 36400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_329
timestamp 1698431365
transform 1 0 38192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_378
timestamp 1698431365
transform 1 0 43680 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_382
timestamp 1698431365
transform 1 0 44128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_419
timestamp 1698431365
transform 1 0 48272 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_34
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_42
timestamp 1698431365
transform 1 0 6048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_59
timestamp 1698431365
transform 1 0 7952 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_67
timestamp 1698431365
transform 1 0 8848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_69
timestamp 1698431365
transform 1 0 9072 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_79
timestamp 1698431365
transform 1 0 10192 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_111
timestamp 1698431365
transform 1 0 13776 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_127
timestamp 1698431365
transform 1 0 15568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_135
timestamp 1698431365
transform 1 0 16464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_150
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_154
timestamp 1698431365
transform 1 0 18592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_156
timestamp 1698431365
transform 1 0 18816 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_189
timestamp 1698431365
transform 1 0 22512 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_205
timestamp 1698431365
transform 1 0 24304 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_227
timestamp 1698431365
transform 1 0 26768 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_231
timestamp 1698431365
transform 1 0 27216 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_233
timestamp 1698431365
transform 1 0 27440 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_270
timestamp 1698431365
transform 1 0 31584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_274
timestamp 1698431365
transform 1 0 32032 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_278
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_356
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_364
timestamp 1698431365
transform 1 0 42112 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_398
timestamp 1698431365
transform 1 0 45920 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_414
timestamp 1698431365
transform 1 0 47712 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_418
timestamp 1698431365
transform 1 0 48160 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_420
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_43
timestamp 1698431365
transform 1 0 6160 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_59
timestamp 1698431365
transform 1 0 7952 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_78
timestamp 1698431365
transform 1 0 10080 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_80
timestamp 1698431365
transform 1 0 10304 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_97
timestamp 1698431365
transform 1 0 12208 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_122
timestamp 1698431365
transform 1 0 15008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_154
timestamp 1698431365
transform 1 0 18592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_158
timestamp 1698431365
transform 1 0 19040 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_192
timestamp 1698431365
transform 1 0 22848 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_196
timestamp 1698431365
transform 1 0 23296 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_230
timestamp 1698431365
transform 1 0 27104 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_238
timestamp 1698431365
transform 1 0 28000 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_242
timestamp 1698431365
transform 1 0 28448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_279
timestamp 1698431365
transform 1 0 32592 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_295
timestamp 1698431365
transform 1 0 34384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_299
timestamp 1698431365
transform 1 0 34832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_301
timestamp 1698431365
transform 1 0 35056 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_308
timestamp 1698431365
transform 1 0 35840 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_314
timestamp 1698431365
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_321
timestamp 1698431365
transform 1 0 37296 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_353
timestamp 1698431365
transform 1 0 40880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_357
timestamp 1698431365
transform 1 0 41328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_365
timestamp 1698431365
transform 1 0 42224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_382
timestamp 1698431365
transform 1 0 44128 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_384
timestamp 1698431365
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_419
timestamp 1698431365
transform 1 0 48272 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_18
timestamp 1698431365
transform 1 0 3360 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_26
timestamp 1698431365
transform 1 0 4256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_58
timestamp 1698431365
transform 1 0 7840 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_65
timestamp 1698431365
transform 1 0 8624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_88
timestamp 1698431365
transform 1 0 11200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_90
timestamp 1698431365
transform 1 0 11424 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_129
timestamp 1698431365
transform 1 0 15792 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_137
timestamp 1698431365
transform 1 0 16688 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698431365
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_144
timestamp 1698431365
transform 1 0 17472 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_153
timestamp 1698431365
transform 1 0 18480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_187
timestamp 1698431365
transform 1 0 22288 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_191
timestamp 1698431365
transform 1 0 22736 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_193
timestamp 1698431365
transform 1 0 22960 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_196
timestamp 1698431365
transform 1 0 23296 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_204
timestamp 1698431365
transform 1 0 24192 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_208
timestamp 1698431365
transform 1 0 24640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_218
timestamp 1698431365
transform 1 0 25760 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_234
timestamp 1698431365
transform 1 0 27552 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_257
timestamp 1698431365
transform 1 0 30128 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_261
timestamp 1698431365
transform 1 0 30576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_263
timestamp 1698431365
transform 1 0 30800 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_305
timestamp 1698431365
transform 1 0 35504 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_321
timestamp 1698431365
transform 1 0 37296 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_325
timestamp 1698431365
transform 1 0 37744 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_347
timestamp 1698431365
transform 1 0 40208 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_349
timestamp 1698431365
transform 1 0 40432 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_375
timestamp 1698431365
transform 1 0 43344 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_407
timestamp 1698431365
transform 1 0 46928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_415
timestamp 1698431365
transform 1 0 47824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_419
timestamp 1698431365
transform 1 0 48272 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_83
timestamp 1698431365
transform 1 0 10640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_87
timestamp 1698431365
transform 1 0 11088 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_89
timestamp 1698431365
transform 1 0 11312 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_98
timestamp 1698431365
transform 1 0 12320 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_102
timestamp 1698431365
transform 1 0 12768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_139
timestamp 1698431365
transform 1 0 16912 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_155
timestamp 1698431365
transform 1 0 18704 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_163
timestamp 1698431365
transform 1 0 19600 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_170
timestamp 1698431365
transform 1 0 20384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_194
timestamp 1698431365
transform 1 0 23072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_226
timestamp 1698431365
transform 1 0 26656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_230
timestamp 1698431365
transform 1 0 27104 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_239
timestamp 1698431365
transform 1 0 28112 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_243
timestamp 1698431365
transform 1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_255
timestamp 1698431365
transform 1 0 29904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_259
timestamp 1698431365
transform 1 0 30352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_311
timestamp 1698431365
transform 1 0 36176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_333
timestamp 1698431365
transform 1 0 38640 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_341
timestamp 1698431365
transform 1 0 39536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_345
timestamp 1698431365
transform 1 0 39984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_349
timestamp 1698431365
transform 1 0 40432 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_357
timestamp 1698431365
transform 1 0 41328 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_363
timestamp 1698431365
transform 1 0 42000 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_380
timestamp 1698431365
transform 1 0 43904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698431365
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_419
timestamp 1698431365
transform 1 0 48272 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_92
timestamp 1698431365
transform 1 0 11648 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_114
timestamp 1698431365
transform 1 0 14112 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_130
timestamp 1698431365
transform 1 0 15904 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_138
timestamp 1698431365
transform 1 0 16800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_157
timestamp 1698431365
transform 1 0 18928 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_173
timestamp 1698431365
transform 1 0 20720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_177
timestamp 1698431365
transform 1 0 21168 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_271
timestamp 1698431365
transform 1 0 31696 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_279
timestamp 1698431365
transform 1 0 32592 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_288
timestamp 1698431365
transform 1 0 33600 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_292
timestamp 1698431365
transform 1 0 34048 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_330
timestamp 1698431365
transform 1 0 38304 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_346
timestamp 1698431365
transform 1 0 40096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_360
timestamp 1698431365
transform 1 0 41664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_362
timestamp 1698431365
transform 1 0 41888 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_393
timestamp 1698431365
transform 1 0 45360 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_409
timestamp 1698431365
transform 1 0 47152 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_417
timestamp 1698431365
transform 1 0 48048 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_53
timestamp 1698431365
transform 1 0 7280 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_57
timestamp 1698431365
transform 1 0 7728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_59
timestamp 1698431365
transform 1 0 7952 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_123
timestamp 1698431365
transform 1 0 15120 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_161
timestamp 1698431365
transform 1 0 19376 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_165
timestamp 1698431365
transform 1 0 19824 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_213
timestamp 1698431365
transform 1 0 25200 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_221
timestamp 1698431365
transform 1 0 26096 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_225
timestamp 1698431365
transform 1 0 26544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_227
timestamp 1698431365
transform 1 0 26768 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_311
timestamp 1698431365
transform 1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_347
timestamp 1698431365
transform 1 0 40208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_349
timestamp 1698431365
transform 1 0 40432 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_365
timestamp 1698431365
transform 1 0 42224 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_375
timestamp 1698431365
transform 1 0 43344 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_383
timestamp 1698431365
transform 1 0 44240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_419
timestamp 1698431365
transform 1 0 48272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1698431365
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_78
timestamp 1698431365
transform 1 0 10080 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_82
timestamp 1698431365
transform 1 0 10528 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_90
timestamp 1698431365
transform 1 0 11424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_94
timestamp 1698431365
transform 1 0 11872 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_102
timestamp 1698431365
transform 1 0 12768 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_135
timestamp 1698431365
transform 1 0 16464 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_139
timestamp 1698431365
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_148
timestamp 1698431365
transform 1 0 17920 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_180
timestamp 1698431365
transform 1 0 21504 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_196
timestamp 1698431365
transform 1 0 23296 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_204
timestamp 1698431365
transform 1 0 24192 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_208
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_227
timestamp 1698431365
transform 1 0 26768 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_231
timestamp 1698431365
transform 1 0 27216 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_238
timestamp 1698431365
transform 1 0 28000 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_254
timestamp 1698431365
transform 1 0 29792 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_263
timestamp 1698431365
transform 1 0 30800 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_290
timestamp 1698431365
transform 1 0 33824 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_294
timestamp 1698431365
transform 1 0 34272 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_310
timestamp 1698431365
transform 1 0 36064 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_318
timestamp 1698431365
transform 1 0 36960 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_322
timestamp 1698431365
transform 1 0 37408 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_338
timestamp 1698431365
transform 1 0 39200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_342
timestamp 1698431365
transform 1 0 39648 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_346
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_349
timestamp 1698431365
transform 1 0 40432 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_416
timestamp 1698431365
transform 1 0 47936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_420
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_69
timestamp 1698431365
transform 1 0 9072 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_73
timestamp 1698431365
transform 1 0 9520 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_111
timestamp 1698431365
transform 1 0 13776 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_127
timestamp 1698431365
transform 1 0 15568 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_135
timestamp 1698431365
transform 1 0 16464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_139
timestamp 1698431365
transform 1 0 16912 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_155
timestamp 1698431365
transform 1 0 18704 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_183
timestamp 1698431365
transform 1 0 21840 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_191
timestamp 1698431365
transform 1 0 22736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_225
timestamp 1698431365
transform 1 0 26544 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_241
timestamp 1698431365
transform 1 0 28336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_263
timestamp 1698431365
transform 1 0 30800 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_307
timestamp 1698431365
transform 1 0 35728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_311
timestamp 1698431365
transform 1 0 36176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_321
timestamp 1698431365
transform 1 0 37296 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_368
timestamp 1698431365
transform 1 0 42560 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_384
timestamp 1698431365
transform 1 0 44352 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_419
timestamp 1698431365
transform 1 0 48272 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_104
timestamp 1698431365
transform 1 0 12992 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_120
timestamp 1698431365
transform 1 0 14784 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_128
timestamp 1698431365
transform 1 0 15680 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_138
timestamp 1698431365
transform 1 0 16800 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_144
timestamp 1698431365
transform 1 0 17472 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_147
timestamp 1698431365
transform 1 0 17808 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_170
timestamp 1698431365
transform 1 0 20384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_172
timestamp 1698431365
transform 1 0 20608 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_188
timestamp 1698431365
transform 1 0 22400 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_192
timestamp 1698431365
transform 1 0 22848 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_200
timestamp 1698431365
transform 1 0 23744 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_208
timestamp 1698431365
transform 1 0 24640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_228
timestamp 1698431365
transform 1 0 26880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_245
timestamp 1698431365
transform 1 0 28784 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_268
timestamp 1698431365
transform 1 0 31360 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_276
timestamp 1698431365
transform 1 0 32256 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698431365
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_297
timestamp 1698431365
transform 1 0 34608 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_313
timestamp 1698431365
transform 1 0 36400 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_317
timestamp 1698431365
transform 1 0 36848 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_346
timestamp 1698431365
transform 1 0 40096 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_416
timestamp 1698431365
transform 1 0 47936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_420
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_207
timestamp 1698431365
transform 1 0 24528 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_277
timestamp 1698431365
transform 1 0 32368 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_309
timestamp 1698431365
transform 1 0 35952 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_313
timestamp 1698431365
transform 1 0 36400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_347
timestamp 1698431365
transform 1 0 40208 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_351
timestamp 1698431365
transform 1 0 40656 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_383
timestamp 1698431365
transform 1 0 44240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_419
timestamp 1698431365
transform 1 0 48272 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_36
timestamp 1698431365
transform 1 0 5376 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_70
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_104
timestamp 1698431365
transform 1 0 12992 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_138
timestamp 1698431365
transform 1 0 16800 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_172
timestamp 1698431365
transform 1 0 20608 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_174
timestamp 1698431365
transform 1 0 20832 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_177
timestamp 1698431365
transform 1 0 21168 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_181
timestamp 1698431365
transform 1 0 21616 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_197
timestamp 1698431365
transform 1 0 23408 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_201
timestamp 1698431365
transform 1 0 23856 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_203
timestamp 1698431365
transform 1 0 24080 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_222
timestamp 1698431365
transform 1 0 26208 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_224
timestamp 1698431365
transform 1 0 26432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_231
timestamp 1698431365
transform 1 0 27216 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_235
timestamp 1698431365
transform 1 0 27664 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_237
timestamp 1698431365
transform 1 0 27888 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_240
timestamp 1698431365
transform 1 0 28224 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_244
timestamp 1698431365
transform 1 0 28672 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_247
timestamp 1698431365
transform 1 0 29008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_249
timestamp 1698431365
transform 1 0 29232 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_256
timestamp 1698431365
transform 1 0 30016 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_274
timestamp 1698431365
transform 1 0 32032 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_276
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_283
timestamp 1698431365
transform 1 0 33040 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_299
timestamp 1698431365
transform 1 0 34832 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_303
timestamp 1698431365
transform 1 0 35280 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_305
timestamp 1698431365
transform 1 0 35504 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_308
timestamp 1698431365
transform 1 0 35840 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_342
timestamp 1698431365
transform 1 0 39648 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_376
timestamp 1698431365
transform 1 0 43456 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_410
timestamp 1698431365
transform 1 0 47264 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_418
timestamp 1698431365
transform 1 0 48160 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_420
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold2 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14224 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 17808 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 16240 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 20384 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform 1 0 18816 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform 1 0 21504 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 25648 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform -1 0 20608 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 10976 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform 1 0 13552 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold13
timestamp 1698431365
transform -1 0 19600 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold14
timestamp 1698431365
transform -1 0 14224 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold15
timestamp 1698431365
transform -1 0 16352 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 2240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698431365
transform 1 0 7952 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 7280 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform -1 0 9744 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 6608 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 3584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 2912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 14560 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input9
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 6720 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 5264 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45584 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698431365
transform 1 0 39088 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output16
timestamp 1698431365
transform 1 0 34944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform -1 0 32592 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform 1 0 26768 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform 1 0 25088 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform -1 0 27440 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 21280 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_60 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 48720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 48720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 48720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 48720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 48720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 48720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 48720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 48720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 48720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 48720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 48720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 48720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 48720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 48720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 48720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 48720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 48720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 48720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 48720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 48720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 48720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 48720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 48720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 48720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 48720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 48720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 48720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 48720 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 48720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 48720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 48720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 48720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 48720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 48720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 48720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 48720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 48720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 48720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 48720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 48720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 48720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 48720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 48720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 48720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 48720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 48720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 48720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 48720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 48720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 48720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 48720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 48720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 48720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 48720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 48720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 48720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 48720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 48720 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 48720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 48720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_122
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_123
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_124
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_125
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_126
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_127
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_128
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_129
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_130
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_131
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_132
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_133
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_134
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_135
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_136
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_137
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_138
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_139
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_140
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_141
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_142
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_143
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_144
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_145
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_146
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_147
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_148
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_149
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_150
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_151
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_152
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_153
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_154
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_155
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_156
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_157
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_158
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_159
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_160
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_161
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_162
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_163
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_164
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_165
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_166
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_167
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_168
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_169
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_170
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_171
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_173
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_174
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_175
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_176
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_177
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_178
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_179
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_180
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_181
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_182
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_183
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_184
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_185
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_186
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_187
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_188
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_189
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_190
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_191
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_192
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_193
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_194
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_195
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_196
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_197
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_198
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_199
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_200
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_201
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_202
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_203
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_204
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_205
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_206
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_207
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_208
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_209
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_210
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_211
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_212
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_213
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_214
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_215
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_216
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_217
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_218
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_219
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_220
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_221
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_222
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_223
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_224
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_225
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_226
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_227
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_228
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_229
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_230
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_231
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_232
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_233
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_234
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_235
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_236
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_237
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_238
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_239
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_240
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_241
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_242
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_243
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_244
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_245
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_246
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_247
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_248
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_249
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_250
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_251
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_252
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_253
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_254
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_255
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_256
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_257
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_258
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_259
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_260
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_261
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_262
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_263
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_264
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_265
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_266
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_267
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_268
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_269
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_270
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_271
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_272
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_273
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_274
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_275
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_276
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_277
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_278
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_279
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_280
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_281
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_282
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_283
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_284
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_285
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_286
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_287
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_288
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_289
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_290
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_291
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_292
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_293
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_294
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_295
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_296
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_297
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_298
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_299
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_300
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_301
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_302
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_303
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_304
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_305
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_306
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_307
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_308
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_309
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_310
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_311
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_312
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_313
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_314
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_315
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_316
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_317
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_318
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_319
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_320
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_321
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_322
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_323
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_324
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_325
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_326
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_327
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_328
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_329
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_330
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_331
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_332
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_333
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_334
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_335
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_336
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_337
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_338
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_339
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_340
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_341
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_342
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_343
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_344
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_345
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_346
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_347
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_348
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_349
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_350
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_351
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_352
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_353
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_354
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_355
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_356
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_357
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_358
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_359
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_360
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_361
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_362
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_363
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_364
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_365
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_366
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_367
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_368
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_369
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_370
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_371
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_372
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_373
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_374
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_375
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_376
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_377
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_378
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_379
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_380
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_381
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_382
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_383
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_384
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_385
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_386
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_387
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_388
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_389
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_390
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_391
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_392
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_393
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_394
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_395
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_396
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_397
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_398
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_399
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_400
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_401
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_402
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_403
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_404
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_405
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_406
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_407
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_408
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_409
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_410
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_411
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_412
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_413
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_414
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_415
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_416
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_417
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_418
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_419
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_420
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_421
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_422
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_423
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_424
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_425
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_426
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_427
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_428
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_429
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_430
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_431
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_432
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_433
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_434
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_435
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_436
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_437
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_438
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_439
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_440
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_441
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_442
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_443
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_444
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_445
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_446
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_447
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_448
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_449
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_450
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_451
timestamp 1698431365
transform 1 0 5152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_452
timestamp 1698431365
transform 1 0 8960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_453
timestamp 1698431365
transform 1 0 12768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_454
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_455
timestamp 1698431365
transform 1 0 20384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_456
timestamp 1698431365
transform 1 0 24192 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_457
timestamp 1698431365
transform 1 0 28000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_458
timestamp 1698431365
transform 1 0 31808 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_459
timestamp 1698431365
transform 1 0 35616 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_460
timestamp 1698431365
transform 1 0 39424 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_461
timestamp 1698431365
transform 1 0 43232 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_462
timestamp 1698431365
transform 1 0 47040 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_vga_spi_rom_26 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 47712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_vga_spi_rom_27
timestamp 1698431365
transform -1 0 41776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_vga_spi_rom_28
timestamp 1698431365
transform -1 0 43008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_vga_spi_rom_29
timestamp 1698431365
transform -1 0 39200 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_vga_spi_rom_30
timestamp 1698431365
transform -1 0 35168 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_vga_spi_rom_31
timestamp 1698431365
transform -1 0 34720 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  top_vga_spi_rom_32 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  top_vga_spi_rom_33
timestamp 1698431365
transform -1 0 45136 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  top_vga_spi_rom_34
timestamp 1698431365
transform -1 0 46816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  top_vga_spi_rom_35
timestamp 1698431365
transform -1 0 35616 0 -1 4704
box -86 -86 534 870
<< labels >>
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 3136 0 3248 800 0 FreeSans 448 90 0 0 rst
port 1 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 ui_in[0]
port 2 nsew signal input
flabel metal2 s 10976 0 11088 800 0 FreeSans 448 90 0 0 ui_in[1]
port 3 nsew signal input
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 ui_in[2]
port 4 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 ui_in[3]
port 5 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 ui_in[4]
port 6 nsew signal input
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 ui_in[5]
port 7 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 ui_in[6]
port 8 nsew signal input
flabel metal2 s 4256 0 4368 800 0 FreeSans 448 90 0 0 ui_in[7]
port 9 nsew signal input
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 uio_in[0]
port 10 nsew signal input
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 uio_in[1]
port 11 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 uio_in[2]
port 12 nsew signal input
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 uio_in[3]
port 13 nsew signal input
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 uio_in[4]
port 14 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 uio_in[5]
port 15 nsew signal input
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 uio_in[6]
port 16 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 uio_in[7]
port 17 nsew signal input
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 uio_oe[0]
port 18 nsew signal tristate
flabel metal2 s 46816 0 46928 800 0 FreeSans 448 90 0 0 uio_oe[1]
port 19 nsew signal tristate
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 uio_oe[2]
port 20 nsew signal tristate
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 uio_oe[3]
port 21 nsew signal tristate
flabel metal2 s 43456 0 43568 800 0 FreeSans 448 90 0 0 uio_oe[4]
port 22 nsew signal tristate
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 uio_oe[5]
port 23 nsew signal tristate
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 uio_oe[6]
port 24 nsew signal tristate
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 uio_oe[7]
port 25 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 uio_out[0]
port 26 nsew signal tristate
flabel metal2 s 37856 0 37968 800 0 FreeSans 448 90 0 0 uio_out[1]
port 27 nsew signal tristate
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 uio_out[2]
port 28 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 uio_out[3]
port 29 nsew signal tristate
flabel metal2 s 34496 0 34608 800 0 FreeSans 448 90 0 0 uio_out[4]
port 30 nsew signal tristate
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 uio_out[5]
port 31 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 uio_out[6]
port 32 nsew signal tristate
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 uio_out[7]
port 33 nsew signal tristate
flabel metal2 s 30016 0 30128 800 0 FreeSans 448 90 0 0 uo_out[0]
port 34 nsew signal tristate
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 uo_out[1]
port 35 nsew signal tristate
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 uo_out[2]
port 36 nsew signal tristate
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 uo_out[3]
port 37 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 uo_out[4]
port 38 nsew signal tristate
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 uo_out[5]
port 39 nsew signal tristate
flabel metal2 s 23296 0 23408 800 0 FreeSans 448 90 0 0 uo_out[6]
port 40 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 uo_out[7]
port 41 nsew signal tristate
flabel metal4 s 4448 3076 4768 50236 0 FreeSans 1280 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 35168 3076 35488 50236 0 FreeSans 1280 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 19808 3076 20128 50236 0 FreeSans 1280 90 0 0 vss
port 43 nsew ground bidirectional
rlabel metal1 25032 49392 25032 49392 0 vdd
rlabel metal1 25032 50176 25032 50176 0 vss
rlabel metal2 9576 5320 9576 5320 0 _0000_
rlabel metal2 22568 12992 22568 12992 0 _0001_
rlabel metal3 23800 11256 23800 11256 0 _0002_
rlabel metal3 23800 9912 23800 9912 0 _0003_
rlabel metal3 21280 7336 21280 7336 0 _0004_
rlabel metal2 12040 13888 12040 13888 0 _0005_
rlabel metal2 14952 18872 14952 18872 0 _0006_
rlabel metal2 12376 15148 12376 15148 0 _0007_
rlabel metal2 23352 7784 23352 7784 0 _0008_
rlabel metal3 22232 8344 22232 8344 0 _0009_
rlabel metal2 18816 16184 18816 16184 0 _0010_
rlabel metal2 10584 10080 10584 10080 0 _0011_
rlabel metal2 6440 35224 6440 35224 0 _0012_
rlabel metal2 7448 38080 7448 38080 0 _0013_
rlabel metal2 10024 41608 10024 41608 0 _0014_
rlabel metal2 6496 40936 6496 40936 0 _0015_
rlabel metal2 5656 43064 5656 43064 0 _0016_
rlabel metal2 8120 44016 8120 44016 0 _0017_
rlabel metal2 8904 46312 8904 46312 0 _0018_
rlabel metal2 10920 47152 10920 47152 0 _0019_
rlabel metal3 14112 38136 14112 38136 0 _0020_
rlabel metal2 14504 33768 14504 33768 0 _0021_
rlabel metal2 16296 36176 16296 36176 0 _0022_
rlabel metal2 16240 42728 16240 42728 0 _0023_
rlabel metal3 12712 43624 12712 43624 0 _0024_
rlabel metal2 13944 45976 13944 45976 0 _0025_
rlabel metal2 12824 40488 12824 40488 0 _0026_
rlabel metal2 16856 39900 16856 39900 0 _0027_
rlabel metal2 16800 45864 16800 45864 0 _0028_
rlabel metal2 15064 48888 15064 48888 0 _0029_
rlabel metal2 18200 48720 18200 48720 0 _0030_
rlabel metal2 21672 48160 21672 48160 0 _0031_
rlabel metal2 27608 45920 27608 45920 0 _0032_
rlabel metal2 28280 42784 28280 42784 0 _0033_
rlabel metal2 31192 44800 31192 44800 0 _0034_
rlabel metal3 35392 44072 35392 44072 0 _0035_
rlabel metal2 37800 45584 37800 45584 0 _0036_
rlabel metal2 39928 47880 39928 47880 0 _0037_
rlabel metal2 37576 48720 37576 48720 0 _0038_
rlabel metal2 38024 43176 38024 43176 0 _0039_
rlabel metal2 39648 41160 39648 41160 0 _0040_
rlabel metal2 42616 39928 42616 39928 0 _0041_
rlabel metal2 43176 42784 43176 42784 0 _0042_
rlabel metal2 42840 45360 42840 45360 0 _0043_
rlabel metal2 32200 47376 32200 47376 0 _0044_
rlabel metal2 32872 49448 32872 49448 0 _0045_
rlabel metal2 29512 49448 29512 49448 0 _0046_
rlabel metal2 27048 50176 27048 50176 0 _0047_
rlabel metal2 24024 47880 24024 47880 0 _0048_
rlabel metal2 24304 44296 24304 44296 0 _0049_
rlabel metal3 24920 42728 24920 42728 0 _0050_
rlabel metal2 24136 40264 24136 40264 0 _0051_
rlabel metal2 17528 39312 17528 39312 0 _0052_
rlabel metal3 16688 31192 16688 31192 0 _0053_
rlabel metal2 18088 24864 18088 24864 0 _0054_
rlabel metal2 19656 28112 19656 28112 0 _0055_
rlabel metal2 20328 31416 20328 31416 0 _0056_
rlabel metal2 22008 34384 22008 34384 0 _0057_
rlabel metal3 22680 25592 22680 25592 0 _0058_
rlabel metal3 24360 28616 24360 28616 0 _0059_
rlabel metal2 26824 32816 26824 32816 0 _0060_
rlabel metal2 27944 39928 27944 39928 0 _0061_
rlabel metal2 30184 41384 30184 41384 0 _0062_
rlabel metal2 31136 38920 31136 38920 0 _0063_
rlabel metal2 33488 40600 33488 40600 0 _0064_
rlabel metal2 35672 42168 35672 42168 0 _0065_
rlabel metal2 37352 39088 37352 39088 0 _0066_
rlabel metal2 39648 37240 39648 37240 0 _0067_
rlabel metal2 41272 38472 41272 38472 0 _0068_
rlabel metal3 43624 37352 43624 37352 0 _0069_
rlabel metal2 41832 17864 41832 17864 0 _0070_
rlabel metal2 42504 14840 42504 14840 0 _0071_
rlabel metal2 45864 15792 45864 15792 0 _0072_
rlabel metal2 44968 18480 44968 18480 0 _0073_
rlabel metal2 45976 21224 45976 21224 0 _0074_
rlabel metal2 45976 23408 45976 23408 0 _0075_
rlabel metal2 45976 26544 45976 26544 0 _0076_
rlabel metal2 24136 24248 24136 24248 0 _0077_
rlabel metal3 26516 27720 26516 27720 0 _0078_
rlabel metal2 45864 29680 45864 29680 0 _0079_
rlabel metal2 43960 31248 43960 31248 0 _0080_
rlabel metal2 43736 34384 43736 34384 0 _0081_
rlabel metal2 45976 33992 45976 33992 0 _0082_
rlabel metal2 45976 32200 45976 32200 0 _0083_
rlabel metal2 46312 12656 46312 12656 0 _0084_
rlabel metal2 45976 10248 45976 10248 0 _0085_
rlabel metal2 43176 10136 43176 10136 0 _0086_
rlabel metal2 42280 12656 42280 12656 0 _0087_
rlabel metal3 44632 22232 44632 22232 0 _0088_
rlabel metal2 40376 22792 40376 22792 0 _0089_
rlabel metal2 42280 24976 42280 24976 0 _0090_
rlabel metal2 42728 28952 42728 28952 0 _0091_
rlabel metal2 37464 31248 37464 31248 0 _0092_
rlabel metal2 37352 32816 37352 32816 0 _0093_
rlabel metal3 40600 34776 40600 34776 0 _0094_
rlabel metal2 35112 35952 35112 35952 0 _0095_
rlabel metal2 20216 41496 20216 41496 0 _0096_
rlabel metal2 19656 43792 19656 43792 0 _0097_
rlabel metal2 20776 45808 20776 45808 0 _0098_
rlabel metal2 20776 39088 20776 39088 0 _0099_
rlabel metal2 20776 23632 20776 23632 0 _0100_
rlabel metal2 20216 22344 20216 22344 0 _0101_
rlabel metal2 14560 23128 14560 23128 0 _0102_
rlabel metal2 14168 26544 14168 26544 0 _0103_
rlabel metal2 11536 27832 11536 27832 0 _0104_
rlabel metal2 13608 21672 13608 21672 0 _0105_
rlabel metal2 11928 24808 11928 24808 0 _0106_
rlabel metal2 10360 30520 10360 30520 0 _0107_
rlabel metal2 6888 30520 6888 30520 0 _0108_
rlabel metal2 7000 33040 7000 33040 0 _0109_
rlabel metal2 2520 36792 2520 36792 0 _0110_
rlabel metal2 3304 39928 3304 39928 0 _0111_
rlabel metal2 2296 38360 2296 38360 0 _0112_
rlabel metal2 2408 34608 2408 34608 0 _0113_
rlabel metal2 2184 31780 2184 31780 0 _0114_
rlabel metal2 2184 30632 2184 30632 0 _0115_
rlabel metal2 2520 28336 2520 28336 0 _0116_
rlabel metal2 6664 28224 6664 28224 0 _0117_
rlabel metal3 8792 27048 8792 27048 0 _0118_
rlabel metal2 2296 26544 2296 26544 0 _0119_
rlabel metal2 2632 24248 2632 24248 0 _0120_
rlabel metal2 7336 22512 7336 22512 0 _0121_
rlabel metal2 8008 24360 8008 24360 0 _0122_
rlabel metal2 2296 22680 2296 22680 0 _0123_
rlabel metal2 2576 20664 2576 20664 0 _0124_
rlabel metal2 5656 20048 5656 20048 0 _0125_
rlabel metal2 2296 18928 2296 18928 0 _0126_
rlabel metal2 2184 17136 2184 17136 0 _0127_
rlabel metal2 6664 17304 6664 17304 0 _0128_
rlabel metal2 2184 14952 2184 14952 0 _0129_
rlabel metal2 2184 10136 2184 10136 0 _0130_
rlabel metal2 2184 7952 2184 7952 0 _0131_
rlabel metal2 2184 5432 2184 5432 0 _0132_
rlabel metal2 2072 3360 2072 3360 0 _0133_
rlabel metal2 2296 12432 2296 12432 0 _0134_
rlabel metal2 4312 15260 4312 15260 0 _0135_
rlabel metal2 7672 14448 7672 14448 0 _0136_
rlabel metal2 8232 11816 8232 11816 0 _0137_
rlabel metal2 6104 10136 6104 10136 0 _0138_
rlabel metal2 6328 8680 6328 8680 0 _0139_
rlabel metal2 6384 5880 6384 5880 0 _0140_
rlabel metal2 33992 6104 33992 6104 0 _0141_
rlabel metal2 37240 5152 37240 5152 0 _0142_
rlabel metal3 41832 4424 41832 4424 0 _0143_
rlabel metal2 41384 7336 41384 7336 0 _0144_
rlabel metal2 43960 4480 43960 4480 0 _0145_
rlabel metal2 45976 8680 45976 8680 0 _0146_
rlabel metal2 45864 5768 45864 5768 0 _0147_
rlabel metal2 10136 7896 10136 7896 0 _0148_
rlabel metal2 6832 4424 6832 4424 0 _0149_
rlabel metal2 23576 6272 23576 6272 0 _0150_
rlabel metal2 16296 5320 16296 5320 0 _0151_
rlabel metal2 31752 6048 31752 6048 0 _0152_
rlabel metal2 34104 4760 34104 4760 0 _0153_
rlabel metal2 15232 6888 15232 6888 0 _0154_
rlabel metal2 20552 7000 20552 7000 0 _0155_
rlabel metal2 33040 29288 33040 29288 0 _0156_
rlabel metal2 37352 27496 37352 27496 0 _0157_
rlabel metal2 38696 24752 38696 24752 0 _0158_
rlabel metal3 33264 24024 33264 24024 0 _0159_
rlabel metal2 38696 15148 38696 15148 0 _0160_
rlabel metal2 39144 16352 39144 16352 0 _0161_
rlabel metal3 40376 9240 40376 9240 0 _0162_
rlabel metal2 41160 11032 41160 11032 0 _0163_
rlabel metal2 37520 9128 37520 9128 0 _0164_
rlabel metal3 39480 12040 39480 12040 0 _0165_
rlabel metal2 39144 40768 39144 40768 0 _0166_
rlabel metal2 42280 40264 42280 40264 0 _0167_
rlabel metal2 42784 42952 42784 42952 0 _0168_
rlabel metal2 42504 45192 42504 45192 0 _0169_
rlabel metal2 30744 47600 30744 47600 0 _0170_
rlabel metal2 31304 47096 31304 47096 0 _0171_
rlabel metal2 33208 48664 33208 48664 0 _0172_
rlabel metal2 29904 48440 29904 48440 0 _0173_
rlabel metal2 27384 49112 27384 49112 0 _0174_
rlabel metal2 27272 39088 27272 39088 0 _0175_
rlabel metal2 26152 45864 26152 45864 0 _0176_
rlabel metal3 24920 46872 24920 46872 0 _0177_
rlabel metal2 25256 45304 25256 45304 0 _0178_
rlabel metal2 25424 42168 25424 42168 0 _0179_
rlabel metal2 25368 40824 25368 40824 0 _0180_
rlabel metal3 18480 38808 18480 38808 0 _0181_
rlabel metal2 17976 31304 17976 31304 0 _0182_
rlabel metal3 19096 25368 19096 25368 0 _0183_
rlabel metal2 19992 25424 19992 25424 0 _0184_
rlabel metal2 18648 25592 18648 25592 0 _0185_
rlabel metal2 23576 28728 23576 28728 0 _0186_
rlabel metal2 25592 27440 25592 27440 0 _0187_
rlabel metal2 20440 28672 20440 28672 0 _0188_
rlabel metal2 27776 38696 27776 38696 0 _0189_
rlabel metal2 21336 31976 21336 31976 0 _0190_
rlabel metal2 22568 34160 22568 34160 0 _0191_
rlabel metal2 23520 26824 23520 26824 0 _0192_
rlabel metal2 25480 28280 25480 28280 0 _0193_
rlabel metal2 27160 32200 27160 32200 0 _0194_
rlabel metal2 28168 39312 28168 39312 0 _0195_
rlabel metal2 31752 40320 31752 40320 0 _0196_
rlabel metal2 30744 40824 30744 40824 0 _0197_
rlabel metal2 30632 38752 30632 38752 0 _0198_
rlabel metal2 33096 40712 33096 40712 0 _0199_
rlabel metal2 35000 42000 35000 42000 0 _0200_
rlabel metal2 41944 37184 41944 37184 0 _0201_
rlabel metal2 37128 38920 37128 38920 0 _0202_
rlabel metal2 39256 38724 39256 38724 0 _0203_
rlabel metal2 41104 37464 41104 37464 0 _0204_
rlabel metal2 43064 36960 43064 36960 0 _0205_
rlabel metal3 23016 21672 23016 21672 0 _0206_
rlabel metal2 24360 22568 24360 22568 0 _0207_
rlabel metal2 43624 16800 43624 16800 0 _0208_
rlabel metal2 42896 17080 42896 17080 0 _0209_
rlabel metal2 42952 15484 42952 15484 0 _0210_
rlabel metal2 45472 15400 45472 15400 0 _0211_
rlabel metal3 45248 17864 45248 17864 0 _0212_
rlabel metal2 47432 20664 47432 20664 0 _0213_
rlabel metal2 48104 20496 48104 20496 0 _0214_
rlabel metal2 46872 23184 46872 23184 0 _0215_
rlabel metal2 46648 26936 46648 26936 0 _0216_
rlabel metal2 24696 24976 24696 24976 0 _0217_
rlabel metal2 26712 27496 26712 27496 0 _0218_
rlabel metal2 46032 28840 46032 28840 0 _0219_
rlabel metal2 47208 32648 47208 32648 0 _0220_
rlabel metal2 43064 30296 43064 30296 0 _0221_
rlabel metal2 43120 33544 43120 33544 0 _0222_
rlabel metal2 46592 34328 46592 34328 0 _0223_
rlabel metal2 46648 31864 46648 31864 0 _0224_
rlabel metal2 47208 14392 47208 14392 0 _0225_
rlabel metal2 46648 13272 46648 13272 0 _0226_
rlabel metal2 47656 10920 47656 10920 0 _0227_
rlabel metal2 43512 10080 43512 10080 0 _0228_
rlabel metal2 42952 12152 42952 12152 0 _0229_
rlabel metal2 19656 22344 19656 22344 0 _0230_
rlabel metal2 44184 23352 44184 23352 0 _0231_
rlabel metal2 43736 22624 43736 22624 0 _0232_
rlabel metal3 40600 23128 40600 23128 0 _0233_
rlabel metal2 41944 25592 41944 25592 0 _0234_
rlabel metal3 44296 28056 44296 28056 0 _0235_
rlabel metal2 38528 33432 38528 33432 0 _0236_
rlabel metal2 37800 31080 37800 31080 0 _0237_
rlabel metal2 36960 33320 36960 33320 0 _0238_
rlabel metal2 38024 34608 38024 34608 0 _0239_
rlabel metal2 35168 35112 35168 35112 0 _0240_
rlabel metal2 22344 42728 22344 42728 0 _0241_
rlabel metal2 21000 41048 21000 41048 0 _0242_
rlabel metal3 20832 42952 20832 42952 0 _0243_
rlabel metal2 21672 44688 21672 44688 0 _0244_
rlabel metal2 20552 39536 20552 39536 0 _0245_
rlabel metal2 21952 25256 21952 25256 0 _0246_
rlabel metal3 20888 26824 20888 26824 0 _0247_
rlabel metal2 8008 23520 8008 23520 0 _0248_
rlabel metal3 10696 42280 10696 42280 0 _0249_
rlabel metal2 15344 24136 15344 24136 0 _0250_
rlabel metal3 13104 26264 13104 26264 0 _0251_
rlabel metal2 8680 25872 8680 25872 0 _0252_
rlabel metal3 14728 26264 14728 26264 0 _0253_
rlabel metal2 17304 30968 17304 30968 0 _0254_
rlabel metal2 11928 28896 11928 28896 0 _0255_
rlabel metal2 13664 23128 13664 23128 0 _0256_
rlabel metal2 13608 25536 13608 25536 0 _0257_
rlabel metal3 11200 30184 11200 30184 0 _0258_
rlabel metal2 7672 30072 7672 30072 0 _0259_
rlabel metal2 7560 32536 7560 32536 0 _0260_
rlabel metal3 6384 22120 6384 22120 0 _0261_
rlabel metal3 5600 38024 5600 38024 0 _0262_
rlabel metal3 4312 36344 4312 36344 0 _0263_
rlabel metal2 3752 39480 3752 39480 0 _0264_
rlabel metal3 4200 37912 4200 37912 0 _0265_
rlabel metal3 3472 34104 3472 34104 0 _0266_
rlabel metal2 4872 27440 4872 27440 0 _0267_
rlabel metal2 2520 32424 2520 32424 0 _0268_
rlabel metal2 2520 31304 2520 31304 0 _0269_
rlabel metal3 3472 27832 3472 27832 0 _0270_
rlabel metal2 9184 27832 9184 27832 0 _0271_
rlabel metal2 9016 26544 9016 26544 0 _0272_
rlabel metal3 3248 26936 3248 26936 0 _0273_
rlabel metal3 5432 23240 5432 23240 0 _0274_
rlabel metal3 3416 23800 3416 23800 0 _0275_
rlabel metal2 8680 23408 8680 23408 0 _0276_
rlabel metal2 8456 24416 8456 24416 0 _0277_
rlabel metal2 2632 22624 2632 22624 0 _0278_
rlabel metal2 2968 21056 2968 21056 0 _0279_
rlabel metal2 5432 20160 5432 20160 0 _0280_
rlabel metal2 4648 17248 4648 17248 0 _0281_
rlabel metal3 3360 18424 3360 18424 0 _0282_
rlabel metal3 3192 17528 3192 17528 0 _0283_
rlabel metal2 6216 18144 6216 18144 0 _0284_
rlabel metal2 2520 15624 2520 15624 0 _0285_
rlabel metal2 23800 12096 23800 12096 0 _0286_
rlabel metal2 4816 6664 4816 6664 0 _0287_
rlabel metal3 3024 9688 3024 9688 0 _0288_
rlabel metal2 2520 8176 2520 8176 0 _0289_
rlabel metal2 2520 5768 2520 5768 0 _0290_
rlabel metal2 1848 3808 1848 3808 0 _0291_
rlabel metal2 6216 12992 6216 12992 0 _0292_
rlabel metal3 3248 12824 3248 12824 0 _0293_
rlabel metal2 5768 14896 5768 14896 0 _0294_
rlabel metal2 7448 14224 7448 14224 0 _0295_
rlabel metal2 7896 12488 7896 12488 0 _0296_
rlabel metal2 25256 8400 25256 8400 0 _0297_
rlabel metal3 7056 9688 7056 9688 0 _0298_
rlabel metal3 7056 9016 7056 9016 0 _0299_
rlabel metal3 7168 6552 7168 6552 0 _0300_
rlabel metal2 33544 6160 33544 6160 0 _0301_
rlabel metal2 42952 5936 42952 5936 0 _0302_
rlabel metal2 37688 5600 37688 5600 0 _0303_
rlabel metal3 39592 4424 39592 4424 0 _0304_
rlabel metal2 41272 7952 41272 7952 0 _0305_
rlabel metal2 43792 5096 43792 5096 0 _0306_
rlabel metal2 46536 8344 46536 8344 0 _0307_
rlabel metal2 46424 6552 46424 6552 0 _0308_
rlabel metal3 33432 12152 33432 12152 0 _0309_
rlabel metal2 33208 11032 33208 11032 0 _0310_
rlabel metal2 33432 9296 33432 9296 0 _0311_
rlabel metal2 33880 10584 33880 10584 0 _0312_
rlabel metal2 29848 8288 29848 8288 0 _0313_
rlabel metal2 31528 8512 31528 8512 0 _0314_
rlabel metal2 12824 7392 12824 7392 0 _0315_
rlabel metal2 33656 10640 33656 10640 0 _0316_
rlabel metal2 39704 10080 39704 10080 0 _0317_
rlabel metal2 33320 9800 33320 9800 0 _0318_
rlabel metal2 33656 9184 33656 9184 0 _0319_
rlabel metal2 32312 8960 32312 8960 0 _0320_
rlabel metal2 30408 11984 30408 11984 0 _0321_
rlabel metal2 29960 10360 29960 10360 0 _0322_
rlabel metal2 28840 8512 28840 8512 0 _0323_
rlabel metal2 12936 8008 12936 8008 0 _0324_
rlabel metal3 11144 7448 11144 7448 0 _0325_
rlabel metal3 13384 5096 13384 5096 0 _0326_
rlabel metal2 7112 5768 7112 5768 0 _0327_
rlabel metal3 11424 5320 11424 5320 0 _0328_
rlabel metal2 30352 6552 30352 6552 0 _0329_
rlabel metal2 33768 4648 33768 4648 0 _0330_
rlabel metal3 19432 6664 19432 6664 0 _0331_
rlabel metal2 21672 8624 21672 8624 0 _0332_
rlabel metal2 38024 22848 38024 22848 0 _0333_
rlabel metal3 37912 15176 37912 15176 0 _0334_
rlabel metal2 38696 12600 38696 12600 0 _0335_
rlabel metal3 37744 15288 37744 15288 0 _0336_
rlabel metal2 38304 9576 38304 9576 0 _0337_
rlabel metal2 38696 10920 38696 10920 0 _0338_
rlabel metal2 37240 10696 37240 10696 0 _0339_
rlabel metal2 39256 9688 39256 9688 0 _0340_
rlabel metal2 37800 10920 37800 10920 0 _0341_
rlabel metal2 37128 9912 37128 9912 0 _0342_
rlabel metal2 39480 10976 39480 10976 0 _0343_
rlabel metal2 38304 12040 38304 12040 0 _0344_
rlabel metal2 5264 3416 5264 3416 0 _0345_
rlabel metal2 32536 24528 32536 24528 0 _0346_
rlabel metal2 34552 23968 34552 23968 0 _0347_
rlabel metal2 35784 23968 35784 23968 0 _0348_
rlabel metal2 39704 20328 39704 20328 0 _0349_
rlabel metal2 30408 21952 30408 21952 0 _0350_
rlabel metal3 29680 19992 29680 19992 0 _0351_
rlabel metal2 28280 22008 28280 22008 0 _0352_
rlabel metal2 40376 26600 40376 26600 0 _0353_
rlabel metal3 32424 25256 32424 25256 0 _0354_
rlabel metal2 33824 26376 33824 26376 0 _0355_
rlabel metal2 33656 28168 33656 28168 0 _0356_
rlabel metal2 26152 23016 26152 23016 0 _0357_
rlabel metal2 32424 21392 32424 21392 0 _0358_
rlabel metal2 34776 20776 34776 20776 0 _0359_
rlabel metal2 34328 19544 34328 19544 0 _0360_
rlabel metal2 36960 24808 36960 24808 0 _0361_
rlabel metal2 20888 18200 20888 18200 0 _0362_
rlabel metal2 16968 22736 16968 22736 0 _0363_
rlabel metal2 21336 21224 21336 21224 0 _0364_
rlabel metal2 38920 17752 38920 17752 0 _0365_
rlabel metal3 40936 19768 40936 19768 0 _0366_
rlabel metal2 35224 22512 35224 22512 0 _0367_
rlabel metal3 39256 18312 39256 18312 0 _0368_
rlabel metal3 41048 18648 41048 18648 0 _0369_
rlabel metal2 37688 17920 37688 17920 0 _0370_
rlabel metal2 38808 15456 38808 15456 0 _0371_
rlabel metal2 41384 17136 41384 17136 0 _0372_
rlabel metal2 38024 18368 38024 18368 0 _0373_
rlabel metal3 40320 18424 40320 18424 0 _0374_
rlabel metal2 23912 18256 23912 18256 0 _0375_
rlabel metal3 25032 18648 25032 18648 0 _0376_
rlabel metal2 27272 20496 27272 20496 0 _0377_
rlabel metal2 26152 20104 26152 20104 0 _0378_
rlabel metal2 30856 31472 30856 31472 0 _0379_
rlabel metal2 22120 21336 22120 21336 0 _0380_
rlabel metal2 22680 20272 22680 20272 0 _0381_
rlabel metal2 33152 21672 33152 21672 0 _0382_
rlabel metal2 31192 16408 31192 16408 0 _0383_
rlabel metal2 30744 11368 30744 11368 0 _0384_
rlabel metal3 30296 10584 30296 10584 0 _0385_
rlabel metal2 35896 9968 35896 9968 0 _0386_
rlabel metal2 31752 12936 31752 12936 0 _0387_
rlabel metal2 24360 14056 24360 14056 0 _0388_
rlabel metal3 29344 17864 29344 17864 0 _0389_
rlabel metal2 28560 11368 28560 11368 0 _0390_
rlabel metal3 28560 15624 28560 15624 0 _0391_
rlabel metal2 31640 11704 31640 11704 0 _0392_
rlabel metal2 33768 15680 33768 15680 0 _0393_
rlabel metal3 30744 11368 30744 11368 0 _0394_
rlabel metal2 28616 13328 28616 13328 0 _0395_
rlabel metal2 28728 14168 28728 14168 0 _0396_
rlabel metal3 27944 15176 27944 15176 0 _0397_
rlabel metal3 28168 16184 28168 16184 0 _0398_
rlabel metal2 33432 15680 33432 15680 0 _0399_
rlabel metal2 31920 15960 31920 15960 0 _0400_
rlabel metal2 33096 15848 33096 15848 0 _0401_
rlabel metal2 26712 20384 26712 20384 0 _0402_
rlabel metal2 37464 24976 37464 24976 0 _0403_
rlabel metal2 31752 23128 31752 23128 0 _0404_
rlabel metal2 17752 21672 17752 21672 0 _0405_
rlabel metal2 30856 21056 30856 21056 0 _0406_
rlabel metal2 31024 20888 31024 20888 0 _0407_
rlabel metal2 31976 24304 31976 24304 0 _0408_
rlabel metal2 23464 21896 23464 21896 0 _0409_
rlabel metal2 38696 16352 38696 16352 0 _0410_
rlabel metal2 30632 22064 30632 22064 0 _0411_
rlabel metal2 29848 21112 29848 21112 0 _0412_
rlabel metal2 23464 29232 23464 29232 0 _0413_
rlabel metal2 31304 26124 31304 26124 0 _0414_
rlabel metal2 31528 26040 31528 26040 0 _0415_
rlabel metal2 29736 20328 29736 20328 0 _0416_
rlabel metal3 32984 20104 32984 20104 0 _0417_
rlabel metal3 31080 20104 31080 20104 0 _0418_
rlabel metal2 29848 20216 29848 20216 0 _0419_
rlabel metal2 26824 16408 26824 16408 0 _0420_
rlabel metal2 30520 20216 30520 20216 0 _0421_
rlabel metal2 32872 20608 32872 20608 0 _0422_
rlabel metal2 33208 19488 33208 19488 0 _0423_
rlabel metal2 39928 18256 39928 18256 0 _0424_
rlabel metal3 39816 21672 39816 21672 0 _0425_
rlabel metal2 41048 19096 41048 19096 0 _0426_
rlabel metal2 41608 29792 41608 29792 0 _0427_
rlabel metal2 36120 16968 36120 16968 0 _0428_
rlabel metal2 38808 18928 38808 18928 0 _0429_
rlabel metal2 40152 21112 40152 21112 0 _0430_
rlabel metal2 17640 17416 17640 17416 0 _0431_
rlabel metal2 36568 16128 36568 16128 0 _0432_
rlabel metal2 39032 18256 39032 18256 0 _0433_
rlabel metal2 39480 18984 39480 18984 0 _0434_
rlabel metal2 35224 17248 35224 17248 0 _0435_
rlabel metal3 36456 21336 36456 21336 0 _0436_
rlabel metal2 37016 21168 37016 21168 0 _0437_
rlabel metal2 17976 18144 17976 18144 0 _0438_
rlabel metal2 17752 17248 17752 17248 0 _0439_
rlabel metal2 38248 19600 38248 19600 0 _0440_
rlabel metal2 32480 26488 32480 26488 0 _0441_
rlabel metal2 37240 20776 37240 20776 0 _0442_
rlabel metal2 32536 22736 32536 22736 0 _0443_
rlabel metal2 31920 9688 31920 9688 0 _0444_
rlabel metal3 35560 20664 35560 20664 0 _0445_
rlabel metal3 36288 20552 36288 20552 0 _0446_
rlabel metal2 33376 18424 33376 18424 0 _0447_
rlabel via1 33768 19991 33768 19991 0 _0448_
rlabel metal2 26712 19040 26712 19040 0 _0449_
rlabel metal3 34664 17752 34664 17752 0 _0450_
rlabel metal2 20776 27160 20776 27160 0 _0451_
rlabel metal3 25088 21672 25088 21672 0 _0452_
rlabel metal2 29232 18648 29232 18648 0 _0453_
rlabel metal3 26096 21000 26096 21000 0 _0454_
rlabel metal2 38696 29344 38696 29344 0 _0455_
rlabel metal2 15400 34552 15400 34552 0 _0456_
rlabel metal2 26600 20944 26600 20944 0 _0457_
rlabel metal2 26712 21224 26712 21224 0 _0458_
rlabel metal2 15848 18760 15848 18760 0 _0459_
rlabel metal2 25928 19936 25928 19936 0 _0460_
rlabel metal2 26040 20944 26040 20944 0 _0461_
rlabel metal2 25256 18480 25256 18480 0 _0462_
rlabel metal2 26376 20272 26376 20272 0 _0463_
rlabel metal3 29232 14952 29232 14952 0 _0464_
rlabel metal3 32424 21672 32424 21672 0 _0465_
rlabel metal2 33096 22904 33096 22904 0 _0466_
rlabel metal2 32200 21448 32200 21448 0 _0467_
rlabel metal3 32144 19096 32144 19096 0 _0468_
rlabel metal2 33432 19656 33432 19656 0 _0469_
rlabel metal2 34440 22008 34440 22008 0 _0470_
rlabel metal3 33376 23352 33376 23352 0 _0471_
rlabel metal3 38304 23800 38304 23800 0 _0472_
rlabel metal2 37744 22344 37744 22344 0 _0473_
rlabel metal3 37352 21672 37352 21672 0 _0474_
rlabel metal2 38360 22008 38360 22008 0 _0475_
rlabel metal2 37352 21560 37352 21560 0 _0476_
rlabel metal2 37128 21952 37128 21952 0 _0477_
rlabel metal2 36120 21728 36120 21728 0 _0478_
rlabel metal3 35168 21560 35168 21560 0 _0479_
rlabel metal2 29624 24080 29624 24080 0 _0480_
rlabel metal2 24472 30856 24472 30856 0 _0481_
rlabel metal2 24472 17864 24472 17864 0 _0482_
rlabel metal3 30184 22232 30184 22232 0 _0483_
rlabel metal2 30296 24080 30296 24080 0 _0484_
rlabel metal3 40320 22120 40320 22120 0 _0485_
rlabel metal2 30184 23912 30184 23912 0 _0486_
rlabel metal2 31080 23016 31080 23016 0 _0487_
rlabel metal2 34104 21672 34104 21672 0 _0488_
rlabel metal2 33656 20664 33656 20664 0 _0489_
rlabel metal2 35000 9632 35000 9632 0 _0490_
rlabel metal3 26264 5880 26264 5880 0 _0491_
rlabel metal3 18760 36064 18760 36064 0 _0492_
rlabel metal3 9912 37912 9912 37912 0 _0493_
rlabel metal3 10416 26376 10416 26376 0 _0494_
rlabel metal2 18200 29680 18200 29680 0 _0495_
rlabel metal2 11648 23352 11648 23352 0 _0496_
rlabel metal2 23240 34552 23240 34552 0 _0497_
rlabel metal3 32480 9688 32480 9688 0 _0498_
rlabel metal2 26712 17864 26712 17864 0 _0499_
rlabel metal2 33544 16688 33544 16688 0 _0500_
rlabel metal2 32648 16128 32648 16128 0 _0501_
rlabel metal2 34664 15232 34664 15232 0 _0502_
rlabel metal2 27720 12768 27720 12768 0 _0503_
rlabel metal3 35392 15176 35392 15176 0 _0504_
rlabel metal2 35784 15456 35784 15456 0 _0505_
rlabel metal3 31304 12264 31304 12264 0 _0506_
rlabel metal2 30072 17192 30072 17192 0 _0507_
rlabel metal2 30520 16408 30520 16408 0 _0508_
rlabel metal2 30632 15568 30632 15568 0 _0509_
rlabel metal2 31864 12208 31864 12208 0 _0510_
rlabel metal3 9240 4312 9240 4312 0 _0511_
rlabel metal3 10304 6664 10304 6664 0 _0512_
rlabel metal2 22232 16464 22232 16464 0 _0513_
rlabel metal2 15848 10416 15848 10416 0 _0514_
rlabel metal3 11704 8120 11704 8120 0 _0515_
rlabel metal2 11144 5880 11144 5880 0 _0516_
rlabel metal2 28504 17864 28504 17864 0 _0517_
rlabel metal2 27720 16464 27720 16464 0 _0518_
rlabel metal2 27160 16520 27160 16520 0 _0519_
rlabel metal2 26488 16744 26488 16744 0 _0520_
rlabel metal2 24136 18760 24136 18760 0 _0521_
rlabel via2 23800 16968 23800 16968 0 _0522_
rlabel metal2 20776 16800 20776 16800 0 _0523_
rlabel metal2 15848 17304 15848 17304 0 _0524_
rlabel metal3 21000 17864 21000 17864 0 _0525_
rlabel metal3 18144 17416 18144 17416 0 _0526_
rlabel metal2 20832 17640 20832 17640 0 _0527_
rlabel metal3 22008 17528 22008 17528 0 _0528_
rlabel metal2 22400 17416 22400 17416 0 _0529_
rlabel metal2 22456 16240 22456 16240 0 _0530_
rlabel metal2 20888 15624 20888 15624 0 _0531_
rlabel metal2 20160 15512 20160 15512 0 _0532_
rlabel metal3 21112 13720 21112 13720 0 _0533_
rlabel metal3 21112 16072 21112 16072 0 _0534_
rlabel metal2 18760 17472 18760 17472 0 _0535_
rlabel metal2 25928 12544 25928 12544 0 _0536_
rlabel metal2 22960 14840 22960 14840 0 _0537_
rlabel metal3 23520 16632 23520 16632 0 _0538_
rlabel metal2 23296 16856 23296 16856 0 _0539_
rlabel metal2 24024 15596 24024 15596 0 _0540_
rlabel metal3 25760 7448 25760 7448 0 _0541_
rlabel metal2 25592 6384 25592 6384 0 _0542_
rlabel metal3 19824 7448 19824 7448 0 _0543_
rlabel metal2 17360 7224 17360 7224 0 _0544_
rlabel metal2 15176 8344 15176 8344 0 _0545_
rlabel metal2 9688 6160 9688 6160 0 _0546_
rlabel metal2 7672 4200 7672 4200 0 _0547_
rlabel metal2 18256 16856 18256 16856 0 _0548_
rlabel metal2 18536 7504 18536 7504 0 _0549_
rlabel metal3 24976 6104 24976 6104 0 _0550_
rlabel metal2 18144 7448 18144 7448 0 _0551_
rlabel metal2 18312 7000 18312 7000 0 _0552_
rlabel metal2 21448 4424 21448 4424 0 _0553_
rlabel metal2 22456 5768 22456 5768 0 _0554_
rlabel metal2 25312 15960 25312 15960 0 _0555_
rlabel metal2 30632 17360 30632 17360 0 _0556_
rlabel metal2 28896 17528 28896 17528 0 _0557_
rlabel metal2 28280 17192 28280 17192 0 _0558_
rlabel metal2 27888 29848 27888 29848 0 _0559_
rlabel metal2 25928 7840 25928 7840 0 _0560_
rlabel metal2 17752 30464 17752 30464 0 _0561_
rlabel metal2 30632 31360 30632 31360 0 _0562_
rlabel metal2 15400 30744 15400 30744 0 _0563_
rlabel metal2 23856 31080 23856 31080 0 _0564_
rlabel metal2 25256 22624 25256 22624 0 _0565_
rlabel metal2 24248 22512 24248 22512 0 _0566_
rlabel metal2 23912 28448 23912 28448 0 _0567_
rlabel metal2 17528 40096 17528 40096 0 _0568_
rlabel metal3 24752 29176 24752 29176 0 _0569_
rlabel metal3 19096 36120 19096 36120 0 _0570_
rlabel metal2 24360 30184 24360 30184 0 _0571_
rlabel metal2 25480 31080 25480 31080 0 _0572_
rlabel metal2 10808 21896 10808 21896 0 _0573_
rlabel metal2 16632 24920 16632 24920 0 _0574_
rlabel metal2 19096 25088 19096 25088 0 _0575_
rlabel metal2 30632 32816 30632 32816 0 _0576_
rlabel metal2 20104 30576 20104 30576 0 _0577_
rlabel metal2 19376 30744 19376 30744 0 _0578_
rlabel metal2 19656 32312 19656 32312 0 _0579_
rlabel metal2 19432 31080 19432 31080 0 _0580_
rlabel metal2 25704 30688 25704 30688 0 _0581_
rlabel metal2 26152 31416 26152 31416 0 _0582_
rlabel metal2 40936 28280 40936 28280 0 _0583_
rlabel metal2 26488 13608 26488 13608 0 _0584_
rlabel metal2 29848 35112 29848 35112 0 _0585_
rlabel via2 13272 39480 13272 39480 0 _0586_
rlabel metal2 24696 38416 24696 38416 0 _0587_
rlabel metal2 12264 38752 12264 38752 0 _0588_
rlabel metal2 25928 37464 25928 37464 0 _0589_
rlabel metal2 26656 22456 26656 22456 0 _0590_
rlabel metal2 25592 37576 25592 37576 0 _0591_
rlabel metal2 23016 35728 23016 35728 0 _0592_
rlabel metal3 25144 36680 25144 36680 0 _0593_
rlabel metal2 26208 36456 26208 36456 0 _0594_
rlabel metal2 26376 38304 26376 38304 0 _0595_
rlabel metal2 27832 37296 27832 37296 0 _0596_
rlabel metal3 11200 35000 11200 35000 0 _0597_
rlabel metal2 34888 45528 34888 45528 0 _0598_
rlabel metal2 30576 39032 30576 39032 0 _0599_
rlabel metal2 26824 24864 26824 24864 0 _0600_
rlabel metal2 28168 36176 28168 36176 0 _0601_
rlabel metal3 21224 37800 21224 37800 0 _0602_
rlabel metal3 27272 36344 27272 36344 0 _0603_
rlabel metal2 26264 23744 26264 23744 0 _0604_
rlabel metal2 26040 33992 26040 33992 0 _0605_
rlabel metal4 26824 20944 26824 20944 0 _0606_
rlabel metal2 32760 36288 32760 36288 0 _0607_
rlabel metal2 42168 33656 42168 33656 0 _0608_
rlabel metal2 30520 35168 30520 35168 0 _0609_
rlabel metal2 22904 21392 22904 21392 0 _0610_
rlabel metal2 28728 34048 28728 34048 0 _0611_
rlabel metal2 29176 36512 29176 36512 0 _0612_
rlabel metal2 30968 34440 30968 34440 0 _0613_
rlabel metal2 33432 34776 33432 34776 0 _0614_
rlabel metal2 32312 34048 32312 34048 0 _0615_
rlabel metal3 31808 33208 31808 33208 0 _0616_
rlabel metal3 33320 38584 33320 38584 0 _0617_
rlabel metal2 32032 34216 32032 34216 0 _0618_
rlabel metal2 31080 34048 31080 34048 0 _0619_
rlabel metal2 42840 21616 42840 21616 0 _0620_
rlabel via2 43624 20888 43624 20888 0 _0621_
rlabel metal2 43512 21280 43512 21280 0 _0622_
rlabel metal2 43568 22680 43568 22680 0 _0623_
rlabel metal2 40264 28560 40264 28560 0 _0624_
rlabel metal2 40712 27160 40712 27160 0 _0625_
rlabel metal2 39872 26488 39872 26488 0 _0626_
rlabel metal2 41160 27328 41160 27328 0 _0627_
rlabel metal2 43176 19712 43176 19712 0 _0628_
rlabel metal2 46312 19600 46312 19600 0 _0629_
rlabel metal2 44632 23324 44632 23324 0 _0630_
rlabel metal2 40936 29960 40936 29960 0 _0631_
rlabel metal3 41888 40376 41888 40376 0 _0632_
rlabel metal2 41664 35448 41664 35448 0 _0633_
rlabel metal2 41048 28112 41048 28112 0 _0634_
rlabel metal2 17416 25704 17416 25704 0 _0635_
rlabel metal2 39032 32144 39032 32144 0 _0636_
rlabel metal3 16408 18424 16408 18424 0 _0637_
rlabel metal2 27048 32592 27048 32592 0 _0638_
rlabel metal2 26712 30912 26712 30912 0 _0639_
rlabel metal2 18704 40152 18704 40152 0 _0640_
rlabel metal2 40432 24920 40432 24920 0 _0641_
rlabel metal2 42616 21000 42616 21000 0 _0642_
rlabel metal2 14616 40824 14616 40824 0 _0643_
rlabel metal2 19880 36904 19880 36904 0 _0644_
rlabel metal3 19880 35112 19880 35112 0 _0645_
rlabel metal3 22456 33432 22456 33432 0 _0646_
rlabel metal2 16408 36568 16408 36568 0 _0647_
rlabel metal2 26488 36120 26488 36120 0 _0648_
rlabel metal2 18872 35168 18872 35168 0 _0649_
rlabel metal2 19152 34104 19152 34104 0 _0650_
rlabel metal3 17696 33320 17696 33320 0 _0651_
rlabel metal2 19432 33768 19432 33768 0 _0652_
rlabel metal3 22064 33544 22064 33544 0 _0653_
rlabel metal2 25032 33656 25032 33656 0 _0654_
rlabel metal2 12992 39368 12992 39368 0 _0655_
rlabel metal2 11088 37800 11088 37800 0 _0656_
rlabel metal3 12768 31640 12768 31640 0 _0657_
rlabel metal2 12488 37576 12488 37576 0 _0658_
rlabel metal2 12152 22568 12152 22568 0 _0659_
rlabel metal2 11256 36960 11256 36960 0 _0660_
rlabel metal3 11144 37240 11144 37240 0 _0661_
rlabel metal3 13832 36344 13832 36344 0 _0662_
rlabel metal2 11928 39144 11928 39144 0 _0663_
rlabel metal2 12488 38696 12488 38696 0 _0664_
rlabel metal3 21672 26712 21672 26712 0 _0665_
rlabel metal2 10808 36456 10808 36456 0 _0666_
rlabel metal2 12936 36792 12936 36792 0 _0667_
rlabel metal3 13440 36456 13440 36456 0 _0668_
rlabel metal2 15288 34776 15288 34776 0 _0669_
rlabel metal2 25928 23520 25928 23520 0 _0670_
rlabel metal3 22232 35896 22232 35896 0 _0671_
rlabel metal2 22120 36736 22120 36736 0 _0672_
rlabel metal2 19544 37128 19544 37128 0 _0673_
rlabel metal3 20160 22344 20160 22344 0 _0674_
rlabel metal3 21672 36456 21672 36456 0 _0675_
rlabel metal2 22680 35672 22680 35672 0 _0676_
rlabel metal2 30072 36680 30072 36680 0 _0677_
rlabel metal2 30184 35840 30184 35840 0 _0678_
rlabel metal2 29512 35672 29512 35672 0 _0679_
rlabel metal2 29960 35840 29960 35840 0 _0680_
rlabel metal2 28616 35056 28616 35056 0 _0681_
rlabel metal3 41664 31192 41664 31192 0 _0682_
rlabel metal2 40152 32480 40152 32480 0 _0683_
rlabel metal3 40880 31752 40880 31752 0 _0684_
rlabel metal2 40712 31024 40712 31024 0 _0685_
rlabel metal2 40488 30968 40488 30968 0 _0686_
rlabel metal2 41384 31248 41384 31248 0 _0687_
rlabel metal2 41048 31472 41048 31472 0 _0688_
rlabel metal2 42392 41160 42392 41160 0 _0689_
rlabel metal2 42280 32424 42280 32424 0 _0690_
rlabel metal2 40040 32648 40040 32648 0 _0691_
rlabel metal2 26712 34160 26712 34160 0 _0692_
rlabel metal2 26600 32256 26600 32256 0 _0693_
rlabel metal3 26096 29960 26096 29960 0 _0694_
rlabel metal3 30352 13720 30352 13720 0 _0695_
rlabel metal3 36680 12824 36680 12824 0 _0696_
rlabel metal2 38136 8176 38136 8176 0 _0697_
rlabel metal2 35112 11648 35112 11648 0 _0698_
rlabel metal2 43848 8008 43848 8008 0 _0699_
rlabel metal2 34384 9240 34384 9240 0 _0700_
rlabel metal2 30296 11816 30296 11816 0 _0701_
rlabel metal2 25704 15288 25704 15288 0 _0702_
rlabel metal3 11928 20664 11928 20664 0 _0703_
rlabel metal2 9128 17976 9128 17976 0 _0704_
rlabel metal2 13944 18256 13944 18256 0 _0705_
rlabel metal3 10136 18424 10136 18424 0 _0706_
rlabel metal2 18200 22456 18200 22456 0 _0707_
rlabel metal2 10696 20104 10696 20104 0 _0708_
rlabel metal2 9576 16072 9576 16072 0 _0709_
rlabel metal2 10024 16520 10024 16520 0 _0710_
rlabel metal2 10024 17920 10024 17920 0 _0711_
rlabel metal4 25256 23352 25256 23352 0 _0712_
rlabel metal3 12432 18200 12432 18200 0 _0713_
rlabel metal2 12488 17304 12488 17304 0 _0714_
rlabel metal2 12488 18088 12488 18088 0 _0715_
rlabel metal2 12208 17752 12208 17752 0 _0716_
rlabel metal2 10248 15792 10248 15792 0 _0717_
rlabel metal2 11144 16856 11144 16856 0 _0718_
rlabel metal2 11480 19488 11480 19488 0 _0719_
rlabel metal3 13328 18424 13328 18424 0 _0720_
rlabel metal2 25032 19600 25032 19600 0 _0721_
rlabel metal2 10360 24192 10360 24192 0 _0722_
rlabel metal2 10920 25760 10920 25760 0 _0723_
rlabel metal2 11256 24584 11256 24584 0 _0724_
rlabel metal2 9352 27216 9352 27216 0 _0725_
rlabel metal2 26600 25648 26600 25648 0 _0726_
rlabel metal2 11200 28616 11200 28616 0 _0727_
rlabel metal2 12040 24472 12040 24472 0 _0728_
rlabel metal2 10920 23184 10920 23184 0 _0729_
rlabel metal2 10528 23240 10528 23240 0 _0730_
rlabel metal2 10808 23632 10808 23632 0 _0731_
rlabel metal2 8232 22848 8232 22848 0 _0732_
rlabel metal2 9968 24472 9968 24472 0 _0733_
rlabel metal2 10584 24360 10584 24360 0 _0734_
rlabel metal2 16408 24024 16408 24024 0 _0735_
rlabel metal3 10528 37352 10528 37352 0 _0736_
rlabel metal2 11256 33880 11256 33880 0 _0737_
rlabel metal2 11032 32928 11032 32928 0 _0738_
rlabel metal2 10584 32536 10584 32536 0 _0739_
rlabel metal3 12544 32536 12544 32536 0 _0740_
rlabel metal2 11816 34832 11816 34832 0 _0741_
rlabel metal4 12264 33824 12264 33824 0 _0742_
rlabel metal2 5432 31416 5432 31416 0 _0743_
rlabel metal2 11704 32200 11704 32200 0 _0744_
rlabel metal2 13160 32592 13160 32592 0 _0745_
rlabel metal2 16072 25396 16072 25396 0 _0746_
rlabel metal3 21616 20776 21616 20776 0 _0747_
rlabel metal2 13832 29680 13832 29680 0 _0748_
rlabel metal2 15176 21056 15176 21056 0 _0749_
rlabel metal2 14392 24248 14392 24248 0 _0750_
rlabel metal2 17640 26712 17640 26712 0 _0751_
rlabel metal3 17304 23688 17304 23688 0 _0752_
rlabel metal2 17864 27664 17864 27664 0 _0753_
rlabel metal2 17528 27496 17528 27496 0 _0754_
rlabel metal3 21896 25256 21896 25256 0 _0755_
rlabel metal3 18760 27048 18760 27048 0 _0756_
rlabel metal2 17808 26824 17808 26824 0 _0757_
rlabel metal2 25592 25704 25592 25704 0 _0758_
rlabel metal2 24080 37240 24080 37240 0 _0759_
rlabel metal2 23576 36792 23576 36792 0 _0760_
rlabel metal3 23856 36456 23856 36456 0 _0761_
rlabel metal2 23128 36120 23128 36120 0 _0762_
rlabel metal3 24528 34888 24528 34888 0 _0763_
rlabel metal2 27048 35168 27048 35168 0 _0764_
rlabel metal2 27608 34272 27608 34272 0 _0765_
rlabel metal2 34776 33824 34776 33824 0 _0766_
rlabel metal3 28560 34104 28560 34104 0 _0767_
rlabel metal4 27832 34384 27832 34384 0 _0768_
rlabel metal2 25368 26180 25368 26180 0 _0769_
rlabel metal3 25312 24808 25312 24808 0 _0770_
rlabel metal2 40096 29176 40096 29176 0 _0771_
rlabel metal2 39256 28280 39256 28280 0 _0772_
rlabel metal2 27160 25144 27160 25144 0 _0773_
rlabel metal3 27384 25592 27384 25592 0 _0774_
rlabel metal2 33544 32256 33544 32256 0 _0775_
rlabel metal2 32984 32088 32984 32088 0 _0776_
rlabel metal3 40124 33880 40124 33880 0 _0777_
rlabel metal2 32648 32200 32648 32200 0 _0778_
rlabel metal2 28504 26096 28504 26096 0 _0779_
rlabel metal2 44072 19040 44072 19040 0 _0780_
rlabel metal3 43680 26264 43680 26264 0 _0781_
rlabel metal2 45696 21000 45696 21000 0 _0782_
rlabel metal2 42336 26824 42336 26824 0 _0783_
rlabel metal2 40712 24080 40712 24080 0 _0784_
rlabel metal2 41496 24136 41496 24136 0 _0785_
rlabel metal2 39928 27216 39928 27216 0 _0786_
rlabel metal2 40936 26544 40936 26544 0 _0787_
rlabel metal3 40824 25760 40824 25760 0 _0788_
rlabel metal2 26152 25368 26152 25368 0 _0789_
rlabel metal2 25368 23128 25368 23128 0 _0790_
rlabel metal2 25592 20720 25592 20720 0 _0791_
rlabel metal2 25368 15568 25368 15568 0 _0792_
rlabel metal2 26040 14784 26040 14784 0 _0793_
rlabel metal2 26712 11424 26712 11424 0 _0794_
rlabel metal2 19656 9016 19656 9016 0 _0795_
rlabel metal3 25312 5768 25312 5768 0 _0796_
rlabel metal2 26376 6328 26376 6328 0 _0797_
rlabel metal2 28392 7056 28392 7056 0 _0798_
rlabel metal2 29848 6384 29848 6384 0 _0799_
rlabel metal3 28952 5096 28952 5096 0 _0800_
rlabel metal2 25816 7896 25816 7896 0 _0801_
rlabel metal2 27272 6328 27272 6328 0 _0802_
rlabel metal3 29680 5992 29680 5992 0 _0803_
rlabel metal3 30240 3528 30240 3528 0 _0804_
rlabel metal2 23184 5880 23184 5880 0 _0805_
rlabel metal3 22848 3752 22848 3752 0 _0806_
rlabel metal2 24920 4088 24920 4088 0 _0807_
rlabel metal2 19992 3808 19992 3808 0 _0808_
rlabel metal2 17752 4368 17752 4368 0 _0809_
rlabel metal2 18424 6272 18424 6272 0 _0810_
rlabel metal2 25256 5208 25256 5208 0 _0811_
rlabel metal2 21000 7840 21000 7840 0 _0812_
rlabel metal3 23688 7728 23688 7728 0 _0813_
rlabel metal2 20440 7840 20440 7840 0 _0814_
rlabel metal2 22680 12040 22680 12040 0 _0815_
rlabel metal2 27608 12880 27608 12880 0 _0816_
rlabel metal2 37576 11424 37576 11424 0 _0817_
rlabel metal2 27944 13048 27944 13048 0 _0818_
rlabel metal2 27776 12152 27776 12152 0 _0819_
rlabel metal2 26600 12432 26600 12432 0 _0820_
rlabel metal3 18424 9688 18424 9688 0 _0821_
rlabel metal2 16744 12600 16744 12600 0 _0822_
rlabel metal3 22176 12264 22176 12264 0 _0823_
rlabel metal2 18088 11704 18088 11704 0 _0824_
rlabel metal3 18480 15960 18480 15960 0 _0825_
rlabel metal2 15848 16352 15848 16352 0 _0826_
rlabel metal2 18536 16296 18536 16296 0 _0827_
rlabel metal2 16744 17192 16744 17192 0 _0828_
rlabel metal2 16576 16968 16576 16968 0 _0829_
rlabel metal3 18704 17080 18704 17080 0 _0830_
rlabel metal2 19320 16800 19320 16800 0 _0831_
rlabel metal2 18816 16744 18816 16744 0 _0832_
rlabel metal2 20440 15260 20440 15260 0 _0833_
rlabel metal3 20272 13944 20272 13944 0 _0834_
rlabel metal2 18648 16520 18648 16520 0 _0835_
rlabel metal2 19208 16408 19208 16408 0 _0836_
rlabel metal2 19264 11592 19264 11592 0 _0837_
rlabel metal2 19096 9912 19096 9912 0 _0838_
rlabel metal2 23016 11368 23016 11368 0 _0839_
rlabel metal2 23408 9016 23408 9016 0 _0840_
rlabel metal2 20160 13720 20160 13720 0 _0841_
rlabel metal3 22400 11592 22400 11592 0 _0842_
rlabel metal2 22400 11368 22400 11368 0 _0843_
rlabel metal2 20552 10696 20552 10696 0 _0844_
rlabel metal3 20440 10584 20440 10584 0 _0845_
rlabel metal2 21672 10584 21672 10584 0 _0846_
rlabel metal2 22456 10248 22456 10248 0 _0847_
rlabel metal2 19096 13664 19096 13664 0 _0848_
rlabel metal2 21784 9744 21784 9744 0 _0849_
rlabel metal2 20664 8456 20664 8456 0 _0850_
rlabel metal2 16408 14448 16408 14448 0 _0851_
rlabel metal3 19320 14392 19320 14392 0 _0852_
rlabel metal3 16520 13608 16520 13608 0 _0853_
rlabel metal2 15960 14056 15960 14056 0 _0854_
rlabel metal3 14616 13048 14616 13048 0 _0855_
rlabel metal2 19432 9408 19432 9408 0 _0856_
rlabel metal3 14280 8344 14280 8344 0 _0857_
rlabel metal2 21224 9072 21224 9072 0 _0858_
rlabel metal2 18928 8232 18928 8232 0 _0859_
rlabel metal2 17640 12488 17640 12488 0 _0860_
rlabel metal2 15064 12656 15064 12656 0 _0861_
rlabel metal2 15400 16408 15400 16408 0 _0862_
rlabel metal2 13440 13048 13440 13048 0 _0863_
rlabel metal2 16408 8232 16408 8232 0 _0864_
rlabel metal2 16520 9072 16520 9072 0 _0865_
rlabel metal3 17864 8904 17864 8904 0 _0866_
rlabel metal3 21112 9016 21112 9016 0 _0867_
rlabel metal2 17304 8736 17304 8736 0 _0868_
rlabel metal2 18088 9464 18088 9464 0 _0869_
rlabel metal2 18368 8120 18368 8120 0 _0870_
rlabel metal2 17528 9184 17528 9184 0 _0871_
rlabel metal2 18424 11704 18424 11704 0 _0872_
rlabel metal2 19712 14728 19712 14728 0 _0873_
rlabel metal3 16912 12600 16912 12600 0 _0874_
rlabel metal2 15680 15736 15680 15736 0 _0875_
rlabel metal2 14168 10248 14168 10248 0 _0876_
rlabel metal2 16296 15484 16296 15484 0 _0877_
rlabel metal2 14056 10360 14056 10360 0 _0878_
rlabel metal3 20272 14728 20272 14728 0 _0879_
rlabel metal2 19656 12096 19656 12096 0 _0880_
rlabel metal2 16184 10976 16184 10976 0 _0881_
rlabel metal2 16072 11592 16072 11592 0 _0882_
rlabel metal2 16072 15232 16072 15232 0 _0883_
rlabel metal2 15232 15064 15232 15064 0 _0884_
rlabel metal2 15064 11872 15064 11872 0 _0885_
rlabel metal2 13944 10752 13944 10752 0 _0886_
rlabel metal2 10920 10080 10920 10080 0 _0887_
rlabel metal2 26936 16520 26936 16520 0 _0888_
rlabel metal2 23016 20664 23016 20664 0 _0889_
rlabel metal2 22512 29512 22512 29512 0 _0890_
rlabel metal2 16184 28672 16184 28672 0 _0891_
rlabel metal3 7392 34776 7392 34776 0 _0892_
rlabel metal2 8232 37296 8232 37296 0 _0893_
rlabel metal2 27496 44072 27496 44072 0 _0894_
rlabel metal2 12096 42728 12096 42728 0 _0895_
rlabel metal2 7560 40768 7560 40768 0 _0896_
rlabel metal2 9688 41272 9688 41272 0 _0897_
rlabel metal2 6720 39816 6720 39816 0 _0898_
rlabel metal2 6552 42392 6552 42392 0 _0899_
rlabel metal2 8680 43232 8680 43232 0 _0900_
rlabel metal2 12712 45808 12712 45808 0 _0901_
rlabel metal2 10136 45304 10136 45304 0 _0902_
rlabel metal2 11704 46368 11704 46368 0 _0903_
rlabel metal2 15176 33544 15176 33544 0 _0904_
rlabel metal2 14672 39704 14672 39704 0 _0905_
rlabel metal2 23464 20552 23464 20552 0 _0906_
rlabel metal2 14728 39256 14728 39256 0 _0907_
rlabel metal2 14392 38696 14392 38696 0 _0908_
rlabel metal2 15512 31864 15512 31864 0 _0909_
rlabel metal3 16632 37016 16632 37016 0 _0910_
rlabel metal3 16296 33208 16296 33208 0 _0911_
rlabel metal2 16632 35336 16632 35336 0 _0912_
rlabel metal2 15848 37240 15848 37240 0 _0913_
rlabel metal2 13608 43232 13608 43232 0 _0914_
rlabel metal2 13720 45360 13720 45360 0 _0915_
rlabel metal2 15064 40880 15064 40880 0 _0916_
rlabel metal2 17192 38080 17192 38080 0 _0917_
rlabel metal2 20104 48272 20104 48272 0 _0918_
rlabel metal2 17584 45304 17584 45304 0 _0919_
rlabel metal2 17304 47936 17304 47936 0 _0920_
rlabel metal2 18760 48216 18760 48216 0 _0921_
rlabel metal2 21224 47432 21224 47432 0 _0922_
rlabel metal2 30296 45024 30296 45024 0 _0923_
rlabel metal2 30744 44912 30744 44912 0 _0924_
rlabel metal2 27384 46368 27384 46368 0 _0925_
rlabel metal3 28392 43512 28392 43512 0 _0926_
rlabel metal2 31248 43736 31248 43736 0 _0927_
rlabel metal2 35560 44296 35560 44296 0 _0928_
rlabel metal2 38920 45808 38920 45808 0 _0929_
rlabel metal2 38024 45752 38024 45752 0 _0930_
rlabel metal2 38976 47656 38976 47656 0 _0931_
rlabel metal2 37688 48216 37688 48216 0 _0932_
rlabel metal2 38584 43512 38584 43512 0 _0933_
rlabel metal2 43064 44576 43064 44576 0 _0934_
rlabel metal2 2072 1918 2072 1918 0 clk
rlabel metal2 20664 21504 20664 21504 0 clknet_0_clk
rlabel metal2 1736 5992 1736 5992 0 clknet_4_0_0_clk
rlabel metal2 41664 15512 41664 15512 0 clknet_4_10_0_clk
rlabel metal2 39648 22344 39648 22344 0 clknet_4_11_0_clk
rlabel metal2 28728 48216 28728 48216 0 clknet_4_12_0_clk
rlabel metal2 30184 44744 30184 44744 0 clknet_4_13_0_clk
rlabel metal2 45304 30184 45304 30184 0 clknet_4_14_0_clk
rlabel metal2 37128 47432 37128 47432 0 clknet_4_15_0_clk
rlabel metal2 1960 23576 1960 23576 0 clknet_4_1_0_clk
rlabel metal2 19992 19208 19992 19208 0 clknet_4_2_0_clk
rlabel metal3 22512 23912 22512 23912 0 clknet_4_3_0_clk
rlabel metal2 1848 29400 1848 29400 0 clknet_4_4_0_clk
rlabel metal2 1848 38024 1848 38024 0 clknet_4_5_0_clk
rlabel metal3 21896 40376 21896 40376 0 clknet_4_6_0_clk
rlabel metal2 17640 48720 17640 48720 0 clknet_4_7_0_clk
rlabel metal2 38696 6272 38696 6272 0 clknet_4_8_0_clk
rlabel metal3 40264 17640 40264 17640 0 clknet_4_9_0_clk
rlabel metal2 2744 4200 2744 4200 0 net1
rlabel metal2 7224 3696 7224 3696 0 net10
rlabel metal2 17416 5768 17416 5768 0 net11
rlabel metal2 41496 15372 41496 15372 0 net12
rlabel metal2 42504 4200 42504 4200 0 net13
rlabel metal2 25256 6216 25256 6216 0 net14
rlabel metal2 37128 4200 37128 4200 0 net15
rlabel metal2 15400 4816 15400 4816 0 net16
rlabel metal3 19208 3304 19208 3304 0 net17
rlabel metal2 32648 3976 32648 3976 0 net18
rlabel metal2 31640 3864 31640 3864 0 net19
rlabel metal2 23912 12432 23912 12432 0 net2
rlabel metal2 28000 4872 28000 4872 0 net20
rlabel metal3 15120 4480 15120 4480 0 net21
rlabel metal3 22736 3416 22736 3416 0 net22
rlabel metal2 28280 5152 28280 5152 0 net23
rlabel metal3 7896 3472 7896 3472 0 net24
rlabel metal3 17416 6552 17416 6552 0 net25
rlabel metal2 45752 2030 45752 2030 0 net26
rlabel metal2 41384 5992 41384 5992 0 net27
rlabel metal2 40152 2030 40152 2030 0 net28
rlabel metal2 36792 2030 36792 2030 0 net29
rlabel metal2 42168 5432 42168 5432 0 net3
rlabel metal3 33600 4424 33600 4424 0 net30
rlabel metal3 32816 3864 32816 3864 0 net31
rlabel metal2 47992 2058 47992 2058 0 net32
rlabel metal2 44632 854 44632 854 0 net33
rlabel metal3 45024 3416 45024 3416 0 net34
rlabel metal3 34384 4088 34384 4088 0 net35
rlabel metal2 35224 3640 35224 3640 0 net36
rlabel metal2 16632 6944 16632 6944 0 net37
rlabel metal2 15904 6776 15904 6776 0 net38
rlabel metal2 11816 6384 11816 6384 0 net39
rlabel metal2 18760 5936 18760 5936 0 net4
rlabel metal2 14840 5544 14840 5544 0 net40
rlabel metal2 20216 4312 20216 4312 0 net41
rlabel metal2 23016 6608 23016 6608 0 net42
rlabel metal2 22568 5264 22568 5264 0 net43
rlabel metal2 5544 4088 5544 4088 0 net44
rlabel metal3 18984 6888 18984 6888 0 net45
rlabel metal2 8288 5096 8288 5096 0 net46
rlabel metal2 15176 5768 15176 5768 0 net47
rlabel metal2 14168 4368 14168 4368 0 net48
rlabel metal2 10808 3416 10808 3416 0 net49
rlabel metal2 6104 3808 6104 3808 0 net5
rlabel metal3 13048 3416 13048 3416 0 net50
rlabel metal3 5152 3416 5152 3416 0 net6
rlabel metal2 3416 3472 3416 3472 0 net7
rlabel metal2 19096 5208 19096 5208 0 net8
rlabel metal3 25088 15176 25088 15176 0 net9
rlabel metal2 2520 2128 2520 2128 0 rst
rlabel metal2 12152 7896 12152 7896 0 tt_um_algofoogle_vga_spi_rom.hsync
rlabel metal2 9016 5152 9016 5152 0 tt_um_algofoogle_vga_spi_rom.r_hsync
rlabel metal3 25200 4200 25200 4200 0 tt_um_algofoogle_vga_spi_rom.r_rgb\[0\]
rlabel metal2 18424 5432 18424 5432 0 tt_um_algofoogle_vga_spi_rom.r_rgb\[1\]
rlabel metal2 29624 5544 29624 5544 0 tt_um_algofoogle_vga_spi_rom.r_rgb\[2\]
rlabel metal2 31752 5432 31752 5432 0 tt_um_algofoogle_vga_spi_rom.r_rgb\[3\]
rlabel metal2 13944 6216 13944 6216 0 tt_um_algofoogle_vga_spi_rom.r_rgb\[4\]
rlabel metal2 22680 6216 22680 6216 0 tt_um_algofoogle_vga_spi_rom.r_rgb\[5\]
rlabel metal2 11704 6384 11704 6384 0 tt_um_algofoogle_vga_spi_rom.r_vsync
rlabel metal2 8568 36176 8568 36176 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[0\]
rlabel metal2 4760 38668 4760 38668 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[100\]
rlabel metal3 7784 34888 7784 34888 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[101\]
rlabel metal2 3976 31472 3976 31472 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[102\]
rlabel metal2 4760 29904 4760 29904 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[103\]
rlabel metal3 10248 28056 10248 28056 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[104\]
rlabel metal2 9016 28336 9016 28336 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[105\]
rlabel metal3 4928 27048 4928 27048 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[106\]
rlabel metal3 7112 23912 7112 23912 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[107\]
rlabel metal2 9016 24024 9016 24024 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[108\]
rlabel metal3 9912 22232 9912 22232 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[109\]
rlabel metal3 18760 36344 18760 36344 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[10\]
rlabel metal2 5600 24584 5600 24584 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[110\]
rlabel metal2 6440 23184 6440 23184 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[111\]
rlabel metal2 6440 21616 6440 21616 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[112\]
rlabel metal2 7000 20048 7000 20048 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[113\]
rlabel metal3 7000 18984 7000 18984 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[114\]
rlabel metal3 7672 17640 7672 17640 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[115\]
rlabel metal2 7112 17248 7112 17248 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[116\]
rlabel metal2 4984 16408 4984 16408 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[117\]
rlabel metal2 4760 11088 4760 11088 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[118\]
rlabel metal3 7840 16072 7840 16072 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[119\]
rlabel metal2 18312 42728 18312 42728 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[11\]
rlabel metal3 8008 20552 8008 20552 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[120\]
rlabel metal2 3080 5432 3080 5432 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[121\]
rlabel metal3 8232 14728 8232 14728 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[122\]
rlabel metal3 8848 13720 8848 13720 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[123\]
rlabel metal3 11648 14616 11648 14616 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[124\]
rlabel metal2 11032 11872 11032 11872 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[125\]
rlabel metal3 10696 17416 10696 17416 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[126\]
rlabel metal3 10472 16632 10472 16632 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[127\]
rlabel metal3 19656 10864 19656 10864 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[128\]
rlabel metal2 37128 5544 37128 5544 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[129\]
rlabel metal2 14728 42448 14728 42448 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[12\]
rlabel metal2 39480 6664 39480 6664 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[130\]
rlabel metal2 40264 5936 40264 5936 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[131\]
rlabel metal3 43064 6664 43064 6664 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[132\]
rlabel metal2 46872 6944 46872 6944 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[133\]
rlabel metal3 47992 7560 47992 7560 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[134\]
rlabel metal3 46760 6552 46760 6552 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[135\]
rlabel metal3 16688 40488 16688 40488 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[13\]
rlabel metal2 15288 40824 15288 40824 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[14\]
rlabel metal2 19264 41272 19264 41272 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[15\]
rlabel metal2 19264 45640 19264 45640 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[16\]
rlabel metal3 18424 47320 18424 47320 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[17\]
rlabel metal3 21672 47992 21672 47992 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[18\]
rlabel metal2 26936 47040 26936 47040 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[19\]
rlabel metal2 9016 39592 9016 39592 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[1\]
rlabel metal3 29232 45304 29232 45304 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[20\]
rlabel metal3 30408 41832 30408 41832 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[21\]
rlabel metal3 33096 43624 33096 43624 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[22\]
rlabel metal3 37800 45304 37800 45304 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[23\]
rlabel metal2 38640 46760 38640 46760 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[24\]
rlabel metal3 42056 47208 42056 47208 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[25\]
rlabel metal2 40264 44016 40264 44016 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[26\]
rlabel metal2 40712 42280 40712 42280 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[27\]
rlabel metal3 40376 40488 40376 40488 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[28\]
rlabel metal2 43176 40712 43176 40712 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[29\]
rlabel metal2 10584 40152 10584 40152 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[2\]
rlabel metal2 43848 42392 43848 42392 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[30\]
rlabel metal2 31640 45472 31640 45472 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[31\]
rlabel metal2 33488 47992 33488 47992 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[32\]
rlabel metal2 34104 48272 34104 48272 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[33\]
rlabel metal2 27720 47544 27720 47544 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[34\]
rlabel metal2 25704 46032 25704 46032 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[35\]
rlabel metal2 25760 44856 25760 44856 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[36\]
rlabel metal2 25704 41048 25704 41048 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[37\]
rlabel metal2 26936 42280 26936 42280 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[38\]
rlabel metal3 23744 38808 23744 38808 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[39\]
rlabel metal2 7672 40600 7672 40600 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[3\]
rlabel metal2 19656 39144 19656 39144 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[40\]
rlabel metal2 18256 31528 18256 31528 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[41\]
rlabel metal2 20664 24696 20664 24696 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[42\]
rlabel metal2 20552 28448 20552 28448 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[43\]
rlabel metal2 22680 32480 22680 32480 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[44\]
rlabel metal2 24248 30968 24248 30968 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[45\]
rlabel metal2 24640 26488 24640 26488 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[46\]
rlabel metal2 25368 28616 25368 28616 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[47\]
rlabel metal2 28504 33488 28504 33488 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[48\]
rlabel metal2 30296 39592 30296 39592 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[49\]
rlabel via2 7672 42728 7672 42728 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[4\]
rlabel metal2 31640 40712 31640 40712 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[50\]
rlabel metal2 33376 41160 33376 41160 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[51\]
rlabel metal3 35728 41384 35728 41384 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[52\]
rlabel metal3 36176 38920 36176 38920 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[53\]
rlabel metal3 38892 38024 38892 38024 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[54\]
rlabel metal3 40712 37912 40712 37912 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[55\]
rlabel metal2 43456 36680 43456 36680 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[56\]
rlabel metal3 44856 15848 44856 15848 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[57\]
rlabel metal2 44296 18872 44296 18872 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[58\]
rlabel metal3 43288 15960 43288 15960 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[59\]
rlabel metal2 10528 44408 10528 44408 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[5\]
rlabel metal2 46088 18256 46088 18256 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[60\]
rlabel metal2 47768 18760 47768 18760 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[61\]
rlabel metal2 47208 23240 47208 23240 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[62\]
rlabel metal2 48328 24360 48328 24360 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[63\]
rlabel metal2 24584 25536 24584 25536 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[64\]
rlabel metal2 26488 24304 26488 24304 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[65\]
rlabel metal3 38808 28616 38808 28616 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[66\]
rlabel metal2 43400 29848 43400 29848 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[67\]
rlabel metal2 42392 30464 42392 30464 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[68\]
rlabel metal2 43960 33712 43960 33712 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[69\]
rlabel metal2 11256 45416 11256 45416 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[6\]
rlabel metal2 46984 31696 46984 31696 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[70\]
rlabel metal2 47936 15120 47936 15120 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[71\]
rlabel metal2 47768 14056 47768 14056 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[72\]
rlabel metal2 46536 11256 46536 11256 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[73\]
rlabel metal2 45192 16408 45192 16408 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[74\]
rlabel metal2 43736 19152 43736 19152 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[75\]
rlabel metal3 46200 23240 46200 23240 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[76\]
rlabel metal3 42112 24696 42112 24696 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[77\]
rlabel metal2 45248 24920 45248 24920 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[78\]
rlabel metal2 44968 29792 44968 29792 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[79\]
rlabel metal2 12824 46480 12824 46480 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[7\]
rlabel metal2 36344 30464 36344 30464 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[80\]
rlabel metal2 35896 34160 35896 34160 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[81\]
rlabel metal2 38920 34664 38920 34664 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[82\]
rlabel metal2 23128 40824 23128 40824 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[83\]
rlabel metal2 22456 40936 22456 40936 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[84\]
rlabel metal3 22344 43400 22344 43400 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[85\]
rlabel metal3 23464 39592 23464 39592 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[86\]
rlabel metal2 23240 39256 23240 39256 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[87\]
rlabel metal3 22680 23352 22680 23352 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[88\]
rlabel metal2 17752 23688 17752 23688 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[89\]
rlabel metal2 15904 38696 15904 38696 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[8\]
rlabel metal2 16856 23576 16856 23576 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[90\]
rlabel metal2 15232 26264 15232 26264 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[91\]
rlabel metal2 14056 24752 14056 24752 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[92\]
rlabel metal2 15288 21168 15288 21168 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[93\]
rlabel metal2 14056 30576 14056 30576 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[94\]
rlabel metal2 12600 30184 12600 30184 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[95\]
rlabel metal2 8120 32592 8120 32592 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[96\]
rlabel metal2 9016 33488 9016 33488 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[97\]
rlabel metal2 6888 36736 6888 36736 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[98\]
rlabel metal3 7896 38136 7896 38136 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[99\]
rlabel metal3 17920 34104 17920 34104 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_buffer\[9\]
rlabel metal2 36008 24360 36008 24360 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.data_index\[3\]
rlabel metal2 34664 27440 34664 27440 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[0\]
rlabel metal2 35672 27552 35672 27552 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[1\]
rlabel metal2 35280 26488 35280 26488 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[2\]
rlabel metal2 40600 17248 40600 17248 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[4\]
rlabel metal2 40824 18032 40824 18032 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[5\]
rlabel metal2 36120 9800 36120 9800 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[6\]
rlabel metal2 39032 10584 39032 10584 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[7\]
rlabel metal2 29288 8512 29288 8512 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[8\]
rlabel metal3 36624 13048 36624 13048 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.hpos\[9\]
rlabel metal2 28000 8344 28000 8344 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.quad
rlabel metal2 25592 14056 25592 14056 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[0\]
rlabel metal2 21112 15848 21112 15848 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[1\]
rlabel metal2 27552 10584 27552 10584 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[2\]
rlabel metal2 24584 16296 24584 16296 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[3\]
rlabel metal3 16800 17640 16800 17640 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[4\]
rlabel metal3 17808 19320 17808 19320 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[5\]
rlabel metal2 22120 18144 22120 18144 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[6\]
rlabel metal2 35448 17752 35448 17752 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[7\]
rlabel metal2 22008 19600 22008 19600 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.o_vpos\[9\]
rlabel metal2 12488 9688 12488 9688 0 tt_um_algofoogle_vga_spi_rom.vga_spi_rom.vga_sync.vsync
rlabel metal2 12152 2058 12152 2058 0 ui_in[0]
rlabel metal2 11032 910 11032 910 0 ui_in[1]
rlabel metal2 9912 2058 9912 2058 0 ui_in[2]
rlabel metal2 6496 5096 6496 5096 0 ui_in[5]
rlabel metal2 3304 5096 3304 5096 0 ui_in[6]
rlabel metal2 3192 3584 3192 3584 0 ui_in[7]
rlabel metal2 19824 2968 19824 2968 0 uio_in[1]
rlabel metal2 18872 2058 18872 2058 0 uio_in[2]
rlabel metal2 16408 5544 16408 5544 0 uio_in[6]
rlabel metal2 15736 3528 15736 3528 0 uio_in[7]
rlabel metal2 46872 3262 46872 3262 0 uio_oe[1]
rlabel metal3 43512 3640 43512 3640 0 uio_oe[5]
rlabel metal2 39032 854 39032 854 0 uio_out[0]
rlabel metal2 37912 2198 37912 2198 0 uio_out[1]
rlabel metal2 35672 2030 35672 2030 0 uio_out[3]
rlabel metal3 35784 3640 35784 3640 0 uio_out[4]
rlabel metal3 31920 3416 31920 3416 0 uo_out[0]
rlabel metal3 29512 4088 29512 4088 0 uo_out[1]
rlabel metal3 28616 3640 28616 3640 0 uo_out[2]
rlabel metal2 26712 2422 26712 2422 0 uo_out[3]
rlabel metal2 25592 854 25592 854 0 uo_out[4]
rlabel metal2 24696 5208 24696 5208 0 uo_out[5]
rlabel metal2 23352 2058 23352 2058 0 uo_out[6]
rlabel metal2 22232 854 22232 854 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 50087 53671
<< end >>
